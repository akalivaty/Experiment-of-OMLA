//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT64), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT66), .B(G183gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT24), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n204), .B1(new_n206), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT23), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT23), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n212), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n218), .ZN(new_n221));
  NOR2_X1   g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(new_n208), .B2(new_n210), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n204), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n220), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT27), .B(G183gat), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT28), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(new_n205), .B2(KEYINPUT27), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(G190gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n229), .B1(new_n232), .B2(KEYINPUT28), .ZN(new_n233));
  NOR3_X1   g032(.A1(KEYINPUT68), .A2(G169gat), .A3(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI22_X1  g035(.A1(new_n234), .A2(new_n235), .B1(new_n213), .B2(new_n214), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n233), .B(new_n207), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n226), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n240));
  INV_X1    g039(.A(G113gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(G120gat), .ZN(new_n242));
  INV_X1    g041(.A(G120gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(G113gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n240), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(G127gat), .B2(new_n245), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G134gat), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n239), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n239), .A2(new_n248), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n203), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT34), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n254), .A2(KEYINPUT72), .B1(new_n255), .B2(new_n251), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n257), .A3(new_n253), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G15gat), .B(G43gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT70), .ZN(new_n261));
  INV_X1    g060(.A(G71gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(G99gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n203), .A3(new_n250), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT33), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(KEYINPUT32), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n268), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n259), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n256), .A2(new_n258), .A3(new_n269), .A4(new_n270), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT36), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n273), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n275), .ZN(new_n278));
  NAND2_X1  g077(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n226), .A2(new_n238), .ZN(new_n282));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n239), .A2(KEYINPUT75), .A3(G226gat), .A4(G233gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n239), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n283), .B(KEYINPUT74), .Z(new_n289));
  OAI211_X1 g088(.A(new_n284), .B(new_n285), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291));
  INV_X1    g090(.A(G211gat), .ZN(new_n292));
  INV_X1    g091(.A(G218gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n291), .B1(KEYINPUT22), .B2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G211gat), .B(G218gat), .Z(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n287), .A2(new_n283), .B1(new_n239), .B2(new_n289), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n297), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n290), .A2(new_n300), .A3(new_n298), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT30), .ZN(new_n306));
  XNOR2_X1  g105(.A(G8gat), .B(G36gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(G64gat), .B(G92gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n305), .A2(new_n309), .ZN(new_n311));
  INV_X1    g110(.A(new_n309), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n303), .A2(new_n312), .A3(new_n304), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(KEYINPUT30), .A3(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G1gat), .B(G29gat), .Z(new_n315));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322));
  INV_X1    g121(.A(G148gat), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n323), .A2(G141gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(G141gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT2), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n323), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n324), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n329), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n327), .B1(new_n337), .B2(KEYINPUT2), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n330), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AOI211_X1 g138(.A(new_n321), .B(new_n322), .C1(new_n248), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n248), .A2(new_n339), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(new_n322), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n342), .B2(new_n321), .ZN(new_n343));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT79), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n248), .B1(new_n346), .B2(new_n339), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n248), .B(new_n339), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n345), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n351), .A2(KEYINPUT5), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n342), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n350), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n320), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n360));
  OR2_X1    g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n351), .A2(KEYINPUT5), .A3(new_n353), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n319), .A3(new_n357), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n362), .A2(KEYINPUT82), .A3(new_n319), .A4(new_n357), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n365), .A2(new_n359), .A3(new_n360), .A4(new_n366), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n310), .A2(new_n314), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(G78gat), .B(G106gat), .Z(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT31), .B(G50gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT3), .B1(new_n297), .B2(new_n286), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(new_n339), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n339), .A2(new_n346), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n286), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n375), .B2(new_n298), .ZN(new_n376));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G22gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n371), .B1(new_n379), .B2(KEYINPUT83), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n378), .B(G22gat), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n381), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n276), .B(new_n280), .C1(new_n368), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT37), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n309), .B1(new_n305), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n290), .A2(new_n297), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n301), .B2(new_n298), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT38), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n319), .B(KEYINPUT84), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(new_n354), .B2(new_n358), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n365), .A2(new_n395), .A3(new_n360), .A4(new_n366), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n392), .A2(new_n396), .A3(new_n361), .A4(new_n311), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n388), .A2(new_n391), .B1(new_n309), .B2(new_n305), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n400), .A2(KEYINPUT86), .A3(new_n361), .A4(new_n396), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n388), .B1(new_n387), .B2(new_n305), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT38), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n348), .A2(new_n349), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n344), .B1(new_n355), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT39), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n394), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT39), .B1(new_n352), .B2(new_n345), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n409), .B(KEYINPUT85), .Z(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n410), .B2(new_n406), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT40), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n413), .A2(new_n395), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n411), .A2(new_n412), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n314), .A2(new_n414), .A3(new_n310), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n385), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n386), .B1(new_n404), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n277), .A2(new_n384), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n314), .A2(new_n310), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT35), .B1(new_n361), .B2(new_n396), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT35), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n368), .B2(new_n420), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT87), .B1(new_n419), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n368), .A2(new_n420), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT35), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n423), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n397), .A2(new_n398), .B1(KEYINPUT38), .B2(new_n402), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n417), .B1(new_n433), .B2(new_n401), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n431), .B(new_n432), .C1(new_n434), .C2(new_n386), .ZN(new_n435));
  XNOR2_X1  g234(.A(G113gat), .B(G141gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(G197gat), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT11), .B(G169gat), .Z(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n439), .B(KEYINPUT12), .Z(new_n440));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n441));
  NAND2_X1  g240(.A1(G229gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G15gat), .B(G22gat), .ZN(new_n444));
  INV_X1    g243(.A(G1gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT16), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G8gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n444), .A2(G1gat), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT92), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n444), .A2(G1gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n448), .A4(new_n447), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT91), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n456), .A3(new_n447), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n444), .A2(KEYINPUT91), .A3(new_n446), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n458), .A2(G8gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n462));
  INV_X1    g261(.A(G50gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(G43gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(G43gat), .ZN(new_n465));
  INV_X1    g264(.A(G43gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT15), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT14), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(G29gat), .B2(G36gat), .ZN(new_n472));
  INV_X1    g271(.A(G29gat), .ZN(new_n473));
  INV_X1    g272(.A(G36gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT14), .ZN(new_n475));
  NAND2_X1  g274(.A1(G29gat), .A2(G36gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT90), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n479));
  AND4_X1   g278(.A1(new_n472), .A2(new_n475), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n466), .A2(G50gat), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n465), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n482), .A3(new_n481), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n470), .B(new_n480), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n483), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n475), .A2(new_n472), .A3(new_n476), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(KEYINPUT15), .A3(new_n488), .A4(new_n484), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  AOI211_X1 g289(.A(new_n441), .B(new_n443), .C1(new_n461), .C2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(KEYINPUT17), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n486), .A2(new_n494), .A3(new_n489), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n451), .A2(new_n454), .B1(new_n457), .B2(new_n459), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n486), .A2(new_n494), .A3(new_n489), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n494), .B1(new_n486), .B2(new_n489), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n492), .B(new_n497), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n491), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n461), .A2(new_n490), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n497), .A2(new_n489), .A3(new_n486), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n442), .B(KEYINPUT13), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT93), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n501), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n443), .B1(new_n461), .B2(new_n490), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT18), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n440), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n498), .B2(new_n502), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n441), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n512), .A2(new_n491), .B1(new_n506), .B2(new_n507), .ZN(new_n518));
  INV_X1    g317(.A(new_n440), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n428), .A2(new_n435), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT94), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n428), .A2(new_n435), .A3(new_n524), .A4(new_n521), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G57gat), .B(G64gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G78gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n262), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G71gat), .A2(G78gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT9), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n531), .B(new_n530), .C1(new_n527), .C2(new_n533), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G127gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n497), .B1(new_n538), .B2(new_n537), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G183gat), .B(G211gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT95), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n549));
  INV_X1    g348(.A(G155gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n548), .B(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n552), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT8), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(G99gat), .B2(G106gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT99), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  NAND2_X1  g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT8), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G99gat), .B(G106gat), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT7), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT98), .ZN(new_n569));
  AND2_X1   g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n568), .A2(KEYINPUT97), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n568), .A2(KEYINPUT97), .A3(KEYINPUT98), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(new_n570), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n565), .A2(new_n567), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n567), .B1(new_n565), .B2(new_n574), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n577), .A2(new_n490), .B1(KEYINPUT41), .B2(new_n579), .ZN(new_n580));
  OAI22_X1  g379(.A1(new_n499), .A2(new_n500), .B1(new_n575), .B2(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G190gat), .B(G218gat), .Z(new_n583));
  AND2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT96), .Z(new_n588));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(KEYINPUT100), .A3(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(KEYINPUT100), .Z(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n584), .B2(new_n585), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n555), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G230gat), .ZN(new_n596));
  INV_X1    g395(.A(G233gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n537), .B1(new_n575), .B2(new_n576), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g399(.A(new_n564), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n563), .B1(new_n560), .B2(new_n562), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n574), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n566), .ZN(new_n604));
  INV_X1    g403(.A(new_n537), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n565), .A2(new_n567), .A3(new_n574), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n600), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT10), .A4(new_n606), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n598), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n599), .A2(new_n607), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n610), .B1(new_n611), .B2(new_n598), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n612), .B(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n595), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n526), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n361), .A2(new_n367), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n445), .ZN(G1324gat));
  INV_X1    g420(.A(KEYINPUT42), .ZN(new_n622));
  INV_X1    g421(.A(new_n421), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n526), .A2(new_n623), .A3(new_n617), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT16), .B(G8gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT101), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n622), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(G8gat), .B1(new_n618), .B2(new_n421), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n626), .B1(new_n630), .B2(new_n622), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n630), .B2(new_n626), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n628), .A2(new_n629), .B1(new_n624), .B2(new_n632), .ZN(G1325gat));
  NAND2_X1  g432(.A1(new_n280), .A2(new_n276), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(G15gat), .B1(new_n618), .B2(new_n635), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n277), .A2(G15gat), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n618), .B2(new_n637), .ZN(G1326gat));
  NOR2_X1   g437(.A1(new_n618), .A2(new_n385), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT43), .B(G22gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1327gat));
  INV_X1    g440(.A(KEYINPUT45), .ZN(new_n642));
  INV_X1    g441(.A(new_n555), .ZN(new_n643));
  INV_X1    g442(.A(new_n616), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n594), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT103), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n523), .B2(new_n525), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n619), .A2(G29gat), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n650), .B1(new_n649), .B2(new_n651), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n642), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n526), .A2(new_n647), .A3(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT104), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(KEYINPUT45), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n594), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT105), .B1(new_n424), .B2(new_n426), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n430), .A2(new_n661), .A3(new_n423), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n659), .B1(new_n663), .B2(new_n419), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n428), .A2(new_n435), .A3(KEYINPUT44), .A4(new_n659), .ZN(new_n667));
  INV_X1    g466(.A(new_n619), .ZN(new_n668));
  INV_X1    g467(.A(new_n521), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n645), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n666), .A2(new_n667), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n473), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n672), .B2(new_n671), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n654), .A2(new_n658), .A3(new_n674), .ZN(G1328gat));
  INV_X1    g474(.A(new_n649), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n623), .A2(new_n474), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n676), .A2(KEYINPUT46), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT46), .B1(new_n676), .B2(new_n677), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n666), .A2(new_n667), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n680), .A2(new_n623), .A3(new_n670), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n678), .B(new_n679), .C1(new_n474), .C2(new_n681), .ZN(G1329gat));
  NAND4_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n634), .A4(new_n670), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G43gat), .ZN(new_n684));
  INV_X1    g483(.A(new_n277), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n466), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n676), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n684), .B(KEYINPUT47), .C1(new_n676), .C2(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1330gat));
  NAND4_X1  g490(.A1(new_n666), .A2(new_n667), .A3(new_n384), .A4(new_n670), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G50gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n384), .A2(new_n463), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n676), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT48), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n693), .B(KEYINPUT48), .C1(new_n676), .C2(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1331gat));
  OR2_X1    g498(.A1(new_n663), .A2(new_n419), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n595), .A2(new_n521), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n616), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT107), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n668), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g506(.A1(new_n704), .A2(new_n421), .ZN(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  AND2_X1   g508(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n708), .B2(new_n709), .ZN(G1333gat));
  OAI21_X1  g511(.A(G71gat), .B1(new_n704), .B2(new_n635), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n685), .A2(new_n262), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n704), .B2(new_n714), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g515(.A1(new_n704), .A2(new_n385), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(new_n529), .ZN(G1335gat));
  NOR2_X1   g517(.A1(new_n555), .A2(new_n521), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n700), .A2(new_n659), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g521(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n700), .A2(new_n659), .A3(new_n719), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n619), .A2(G85gat), .A3(new_n644), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n555), .A2(new_n521), .A3(new_n644), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n680), .A2(new_n668), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G85gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  NOR3_X1   g532(.A1(new_n421), .A2(G92gat), .A3(new_n644), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT52), .B1(new_n725), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n680), .A2(new_n623), .A3(new_n728), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G92gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(KEYINPUT51), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n720), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n741), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n700), .A2(new_n659), .A3(new_n719), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n734), .B(KEYINPUT110), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n736), .A2(G92gat), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n738), .B1(new_n739), .B2(new_n747), .ZN(G1337gat));
  NAND3_X1  g547(.A1(new_n680), .A2(new_n634), .A3(new_n728), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G99gat), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n277), .A2(G99gat), .A3(new_n644), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n725), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1338gat));
  NOR3_X1   g552(.A1(new_n385), .A2(G106gat), .A3(new_n644), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT53), .B1(new_n725), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n680), .A2(new_n384), .A3(new_n728), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G106gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n756), .A2(G106gat), .B1(new_n745), .B2(new_n754), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(G1339gat));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n608), .A2(new_n609), .ZN(new_n765));
  INV_X1    g564(.A(new_n598), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT54), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n609), .A2(new_n598), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n768), .B1(new_n770), .B2(new_n608), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n764), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n615), .B1(new_n610), .B2(new_n768), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(new_n773), .B1(new_n612), .B2(new_n615), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n767), .A2(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n773), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n764), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n509), .A2(new_n514), .A3(new_n440), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n519), .B1(new_n517), .B2(new_n518), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n774), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n442), .B1(new_n512), .B2(new_n504), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n506), .A2(new_n507), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n439), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n616), .A2(new_n520), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n659), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n774), .A2(new_n777), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n520), .A2(new_n783), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n786), .A2(new_n594), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n763), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n611), .A2(new_n598), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n767), .A2(new_n790), .A3(new_n615), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n599), .A2(new_n600), .A3(new_n607), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT54), .B1(new_n792), .B2(new_n769), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT55), .B1(new_n793), .B2(new_n610), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n765), .A2(new_n768), .A3(new_n766), .ZN(new_n795));
  INV_X1    g594(.A(new_n615), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n791), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT55), .B1(new_n775), .B2(new_n773), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n520), .A2(new_n783), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n659), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n616), .A2(new_n801), .B1(new_n800), .B2(new_n521), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT112), .B(new_n802), .C1(new_n803), .C2(new_n659), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n804), .A3(new_n643), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n701), .A2(new_n644), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n762), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n762), .A3(new_n806), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n385), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n668), .A2(new_n421), .ZN(new_n811));
  OR3_X1    g610(.A1(new_n810), .A2(new_n277), .A3(new_n811), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT114), .Z(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(G113gat), .A3(new_n521), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n805), .A2(new_n762), .A3(new_n806), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n815), .A2(new_n807), .A3(new_n619), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n421), .A3(new_n420), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n241), .B1(new_n817), .B2(new_n669), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n814), .A2(new_n818), .ZN(G1340gat));
  NAND3_X1  g618(.A1(new_n813), .A2(G120gat), .A3(new_n616), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n243), .B1(new_n817), .B2(new_n644), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(G1341gat));
  INV_X1    g621(.A(new_n813), .ZN(new_n823));
  OAI21_X1  g622(.A(G127gat), .B1(new_n823), .B2(new_n643), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n643), .A2(G127gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n817), .B2(new_n825), .ZN(G1342gat));
  OAI21_X1  g625(.A(G134gat), .B1(new_n823), .B2(new_n594), .ZN(new_n827));
  XOR2_X1   g626(.A(KEYINPUT69), .B(G134gat), .Z(new_n828));
  NAND2_X1  g627(.A1(new_n659), .A2(new_n828), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n817), .A2(new_n829), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n830));
  NAND2_X1  g629(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n830), .B(new_n831), .Z(new_n832));
  NAND2_X1  g631(.A1(new_n827), .A2(new_n832), .ZN(G1343gat));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n815), .A2(new_n807), .A3(new_n385), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT116), .B1(new_n835), .B2(KEYINPUT57), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n808), .A2(new_n384), .A3(new_n809), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n776), .A2(KEYINPUT117), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n776), .A2(KEYINPUT117), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT55), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n521), .A2(new_n774), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n784), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n594), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n643), .B1(new_n846), .B2(new_n788), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n806), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT57), .A3(new_n384), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n836), .A2(new_n840), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n634), .A2(new_n811), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n834), .B1(new_n852), .B2(new_n669), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n850), .A2(KEYINPUT120), .A3(new_n851), .A4(new_n521), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(G141gat), .A3(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n816), .A2(KEYINPUT119), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n816), .A2(KEYINPUT119), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n635), .A2(new_n384), .A3(new_n421), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n669), .A2(G141gat), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(KEYINPUT58), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n852), .A2(KEYINPUT118), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n865), .A3(new_n851), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n521), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n861), .B1(new_n867), .B2(G141gat), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT121), .B(new_n863), .C1(new_n868), .C2(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n851), .A2(new_n616), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n835), .A2(KEYINPUT57), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n876), .A2(KEYINPUT122), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n806), .B(KEYINPUT123), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n847), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n879), .B2(new_n384), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n876), .B1(new_n880), .B2(KEYINPUT122), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n875), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT59), .B1(new_n882), .B2(new_n323), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n864), .A2(new_n866), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(new_n616), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n323), .A2(KEYINPUT59), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n859), .A2(new_n323), .A3(new_n616), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1345gat));
  NAND2_X1  g688(.A1(new_n859), .A2(new_n555), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n550), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n643), .A2(new_n550), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n884), .B2(new_n894), .ZN(G1346gat));
  AOI21_X1  g694(.A(G162gat), .B1(new_n859), .B2(new_n659), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n659), .A2(G162gat), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n884), .B2(new_n897), .ZN(G1347gat));
  NOR3_X1   g697(.A1(new_n815), .A2(new_n807), .A3(new_n668), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n899), .A2(new_n623), .A3(new_n420), .ZN(new_n900));
  AOI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n521), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n668), .A2(new_n421), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n810), .A2(new_n277), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n669), .A2(new_n213), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n900), .B2(new_n616), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n644), .A2(new_n214), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n904), .B2(new_n908), .ZN(G1349gat));
  INV_X1    g708(.A(new_n904), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n205), .B1(new_n910), .B2(new_n643), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n900), .A2(new_n227), .A3(new_n555), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g713(.A(new_n228), .B1(new_n904), .B2(new_n659), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT61), .Z(new_n916));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n228), .A3(new_n659), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n634), .A2(new_n385), .A3(new_n421), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n899), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(G197gat), .B1(new_n921), .B2(new_n521), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n635), .A2(new_n902), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n877), .B2(new_n881), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n521), .A2(G197gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1352gat));
  XNOR2_X1  g725(.A(KEYINPUT125), .B(G204gat), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(KEYINPUT126), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n920), .A2(new_n644), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n930), .B(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n924), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(new_n644), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n934), .B2(new_n927), .ZN(G1353gat));
  NAND3_X1  g734(.A1(new_n921), .A2(new_n292), .A3(new_n555), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n924), .A2(new_n555), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n937), .B2(G211gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g741(.A(KEYINPUT127), .B(new_n936), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1354gat));
  OAI21_X1  g743(.A(G218gat), .B1(new_n933), .B2(new_n594), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n921), .A2(new_n293), .A3(new_n659), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1355gat));
endmodule


