

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(G2104), .A2(n517), .ZN(n886) );
  NOR2_X1 U551 ( .A1(n728), .A2(G1966), .ZN(n592) );
  NAND2_X1 U552 ( .A1(n664), .A2(G8), .ZN(n728) );
  NOR2_X1 U553 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U554 ( .A(n522), .B(n521), .ZN(n893) );
  XOR2_X1 U555 ( .A(KEYINPUT70), .B(n595), .Z(n514) );
  NOR2_X1 U556 ( .A1(n726), .A2(n728), .ZN(n515) );
  OR2_X1 U557 ( .A1(n618), .A2(n770), .ZN(n619) );
  INV_X1 U558 ( .A(KEYINPUT30), .ZN(n647) );
  XNOR2_X1 U559 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U560 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n654) );
  INV_X1 U561 ( .A(KEYINPUT103), .ZN(n662) );
  XNOR2_X1 U562 ( .A(n599), .B(KEYINPUT15), .ZN(n968) );
  XOR2_X1 U563 ( .A(KEYINPUT1), .B(n529), .Z(n799) );
  XNOR2_X1 U564 ( .A(n525), .B(KEYINPUT64), .ZN(n890) );
  NOR2_X1 U565 ( .A1(G651), .A2(n579), .ZN(n800) );
  NOR2_X1 U566 ( .A1(n528), .A2(n527), .ZN(G164) );
  AND2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U568 ( .A1(G114), .A2(n885), .ZN(n516) );
  XOR2_X1 U569 ( .A(KEYINPUT88), .B(n516), .Z(n520) );
  INV_X1 U570 ( .A(G2105), .ZN(n517) );
  NAND2_X1 U571 ( .A1(G126), .A2(n886), .ZN(n518) );
  XNOR2_X1 U572 ( .A(KEYINPUT87), .B(n518), .ZN(n519) );
  NOR2_X1 U573 ( .A1(n520), .A2(n519), .ZN(n524) );
  XNOR2_X1 U574 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n522) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n893), .A2(G138), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U578 ( .A1(G2104), .A2(n517), .ZN(n525) );
  NAND2_X1 U579 ( .A1(G102), .A2(n890), .ZN(n526) );
  XNOR2_X1 U580 ( .A(n526), .B(KEYINPUT89), .ZN(n527) );
  INV_X1 U581 ( .A(G651), .ZN(n532) );
  NOR2_X1 U582 ( .A1(G543), .A2(n532), .ZN(n529) );
  NAND2_X1 U583 ( .A1(G64), .A2(n799), .ZN(n531) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n579) );
  NAND2_X1 U585 ( .A1(G52), .A2(n800), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n537) );
  NOR2_X1 U587 ( .A1(n579), .A2(n532), .ZN(n803) );
  NAND2_X1 U588 ( .A1(G77), .A2(n803), .ZN(n534) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n804) );
  NAND2_X1 U590 ( .A1(G90), .A2(n804), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U592 ( .A(KEYINPUT9), .B(n535), .Z(n536) );
  NOR2_X1 U593 ( .A1(n537), .A2(n536), .ZN(G171) );
  NAND2_X1 U594 ( .A1(n804), .A2(G89), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n538), .B(KEYINPUT4), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G76), .A2(n803), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n541), .B(KEYINPUT5), .ZN(n547) );
  NAND2_X1 U599 ( .A1(n800), .A2(G51), .ZN(n542) );
  XNOR2_X1 U600 ( .A(n542), .B(KEYINPUT72), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G63), .A2(n799), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(n545), .Z(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U605 ( .A(n548), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U606 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U607 ( .A1(G62), .A2(n799), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G75), .A2(n803), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G88), .A2(n804), .ZN(n552) );
  NAND2_X1 U611 ( .A1(G50), .A2(n800), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT83), .B(n555), .Z(G166) );
  INV_X1 U615 ( .A(G166), .ZN(G303) );
  NAND2_X1 U616 ( .A1(G101), .A2(n890), .ZN(n556) );
  XNOR2_X1 U617 ( .A(KEYINPUT23), .B(n556), .ZN(n558) );
  AND2_X1 U618 ( .A1(n886), .A2(G125), .ZN(n557) );
  NOR2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n588) );
  INV_X1 U620 ( .A(KEYINPUT66), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G137), .A2(n893), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G113), .A2(n885), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n565) );
  AND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U626 ( .A1(KEYINPUT66), .A2(n563), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n589) );
  AND2_X1 U628 ( .A1(n588), .A2(n589), .ZN(G160) );
  XOR2_X1 U629 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n567) );
  NAND2_X1 U630 ( .A1(G73), .A2(n803), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G61), .A2(n799), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G86), .A2(n804), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n800), .A2(G48), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(G305) );
  NAND2_X1 U638 ( .A1(G651), .A2(G74), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT80), .B(n574), .Z(n575) );
  NOR2_X1 U640 ( .A1(n799), .A2(n575), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n800), .A2(G49), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT81), .ZN(n581) );
  NAND2_X1 U644 ( .A1(G87), .A2(n579), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(G288) );
  NAND2_X1 U646 ( .A1(G72), .A2(n803), .ZN(n583) );
  NAND2_X1 U647 ( .A1(G85), .A2(n804), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U649 ( .A1(G60), .A2(n799), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G47), .A2(n800), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  OR2_X1 U652 ( .A1(n587), .A2(n586), .ZN(G290) );
  NOR2_X1 U653 ( .A1(G164), .A2(G1384), .ZN(n677) );
  AND2_X1 U654 ( .A1(G40), .A2(n588), .ZN(n590) );
  AND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X2 U656 ( .A1(n677), .A2(n591), .ZN(n664) );
  NOR2_X1 U657 ( .A1(G2084), .A2(n664), .ZN(n645) );
  NAND2_X1 U658 ( .A1(G8), .A2(n645), .ZN(n660) );
  XNOR2_X1 U659 ( .A(n592), .B(KEYINPUT97), .ZN(n644) );
  NAND2_X1 U660 ( .A1(G54), .A2(n800), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G79), .A2(n803), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G92), .A2(n804), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n799), .A2(G66), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n514), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  INV_X1 U667 ( .A(n968), .ZN(n770) );
  INV_X1 U668 ( .A(n664), .ZN(n638) );
  NOR2_X1 U669 ( .A1(n638), .A2(G1348), .ZN(n601) );
  NOR2_X1 U670 ( .A1(G2067), .A2(n664), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n618) );
  NAND2_X1 U672 ( .A1(n770), .A2(n618), .ZN(n617) );
  NAND2_X1 U673 ( .A1(G56), .A2(n799), .ZN(n602) );
  XOR2_X1 U674 ( .A(KEYINPUT14), .B(n602), .Z(n609) );
  NAND2_X1 U675 ( .A1(n804), .A2(G81), .ZN(n603) );
  XOR2_X1 U676 ( .A(KEYINPUT12), .B(n603), .Z(n606) );
  NAND2_X1 U677 ( .A1(n803), .A2(G68), .ZN(n604) );
  XOR2_X1 U678 ( .A(KEYINPUT68), .B(n604), .Z(n605) );
  NOR2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT13), .ZN(n608) );
  NOR2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n800), .A2(G43), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n983) );
  INV_X1 U684 ( .A(G1996), .ZN(n945) );
  NOR2_X1 U685 ( .A1(n664), .A2(n945), .ZN(n612) );
  XOR2_X1 U686 ( .A(n612), .B(KEYINPUT26), .Z(n614) );
  NAND2_X1 U687 ( .A1(n664), .A2(G1341), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U689 ( .A1(n983), .A2(n615), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U692 ( .A(KEYINPUT99), .B(n621), .ZN(n632) );
  NAND2_X1 U693 ( .A1(n638), .A2(G2072), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n622), .B(KEYINPUT27), .ZN(n624) );
  INV_X1 U695 ( .A(G1956), .ZN(n917) );
  NOR2_X1 U696 ( .A1(n917), .A2(n638), .ZN(n623) );
  NOR2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n633) );
  NAND2_X1 U698 ( .A1(G65), .A2(n799), .ZN(n626) );
  NAND2_X1 U699 ( .A1(G53), .A2(n800), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U701 ( .A1(G78), .A2(n803), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G91), .A2(n804), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n811) );
  NAND2_X1 U705 ( .A1(n633), .A2(n811), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n636) );
  NOR2_X1 U707 ( .A1(n633), .A2(n811), .ZN(n634) );
  XOR2_X1 U708 ( .A(n634), .B(KEYINPUT28), .Z(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U710 ( .A(KEYINPUT29), .B(n637), .Z(n643) );
  XOR2_X1 U711 ( .A(KEYINPUT25), .B(G2078), .Z(n951) );
  NAND2_X1 U712 ( .A1(n638), .A2(n951), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G1961), .A2(n664), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U715 ( .A(KEYINPUT98), .B(n641), .Z(n651) );
  NAND2_X1 U716 ( .A1(n651), .A2(G171), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n657) );
  NAND2_X1 U718 ( .A1(G8), .A2(n644), .ZN(n646) );
  NOR2_X1 U719 ( .A1(G168), .A2(n649), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n650), .B(KEYINPUT100), .ZN(n653) );
  NOR2_X1 U721 ( .A1(n651), .A2(G171), .ZN(n652) );
  NOR2_X2 U722 ( .A1(n653), .A2(n652), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U725 ( .A1(n644), .A2(n661), .ZN(n658) );
  XOR2_X1 U726 ( .A(KEYINPUT102), .B(n658), .Z(n659) );
  NAND2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n673) );
  NAND2_X1 U728 ( .A1(G286), .A2(n661), .ZN(n663) );
  XNOR2_X1 U729 ( .A(n663), .B(n662), .ZN(n669) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n728), .ZN(n666) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U733 ( .A1(G303), .A2(n667), .ZN(n668) );
  NAND2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n670), .A2(G8), .ZN(n671) );
  XNOR2_X1 U736 ( .A(n671), .B(KEYINPUT32), .ZN(n672) );
  NAND2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X2 U738 ( .A(n674), .B(KEYINPUT104), .ZN(n724) );
  NOR2_X1 U739 ( .A1(G2090), .A2(G303), .ZN(n675) );
  NAND2_X1 U740 ( .A1(G8), .A2(n675), .ZN(n713) );
  NAND2_X1 U741 ( .A1(G160), .A2(G40), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n751) );
  XNOR2_X1 U743 ( .A(G2067), .B(KEYINPUT37), .ZN(n749) );
  XNOR2_X1 U744 ( .A(KEYINPUT93), .B(KEYINPUT36), .ZN(n690) );
  NAND2_X1 U745 ( .A1(G104), .A2(n890), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n678), .B(KEYINPUT90), .ZN(n680) );
  NAND2_X1 U747 ( .A1(G140), .A2(n893), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n681), .B(KEYINPUT34), .ZN(n682) );
  XNOR2_X1 U750 ( .A(n682), .B(KEYINPUT91), .ZN(n688) );
  XNOR2_X1 U751 ( .A(KEYINPUT35), .B(KEYINPUT92), .ZN(n686) );
  NAND2_X1 U752 ( .A1(G116), .A2(n885), .ZN(n684) );
  NAND2_X1 U753 ( .A1(G128), .A2(n886), .ZN(n683) );
  NAND2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n690), .B(n689), .ZN(n898) );
  NOR2_X1 U758 ( .A1(n749), .A2(n898), .ZN(n998) );
  NAND2_X1 U759 ( .A1(n751), .A2(n998), .ZN(n746) );
  NAND2_X1 U760 ( .A1(G117), .A2(n885), .ZN(n692) );
  NAND2_X1 U761 ( .A1(G129), .A2(n886), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U763 ( .A1(n890), .A2(G105), .ZN(n693) );
  XOR2_X1 U764 ( .A(KEYINPUT38), .B(n693), .Z(n694) );
  NOR2_X1 U765 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U766 ( .A1(n893), .A2(G141), .ZN(n696) );
  NAND2_X1 U767 ( .A1(n697), .A2(n696), .ZN(n880) );
  NAND2_X1 U768 ( .A1(G1996), .A2(n880), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n698), .B(KEYINPUT95), .ZN(n707) );
  NAND2_X1 U770 ( .A1(n893), .A2(G131), .ZN(n700) );
  NAND2_X1 U771 ( .A1(G95), .A2(n890), .ZN(n699) );
  NAND2_X1 U772 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U773 ( .A(KEYINPUT94), .B(n701), .Z(n705) );
  NAND2_X1 U774 ( .A1(G107), .A2(n885), .ZN(n703) );
  NAND2_X1 U775 ( .A1(G119), .A2(n886), .ZN(n702) );
  AND2_X1 U776 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U777 ( .A1(n705), .A2(n704), .ZN(n901) );
  AND2_X1 U778 ( .A1(G1991), .A2(n901), .ZN(n706) );
  NOR2_X1 U779 ( .A1(n707), .A2(n706), .ZN(n1002) );
  XOR2_X1 U780 ( .A(n751), .B(KEYINPUT96), .Z(n708) );
  NOR2_X1 U781 ( .A1(n1002), .A2(n708), .ZN(n742) );
  INV_X1 U782 ( .A(n742), .ZN(n709) );
  AND2_X1 U783 ( .A1(n746), .A2(n709), .ZN(n725) );
  NOR2_X1 U784 ( .A1(G1981), .A2(G305), .ZN(n710) );
  XOR2_X1 U785 ( .A(n710), .B(KEYINPUT24), .Z(n711) );
  NOR2_X1 U786 ( .A1(n728), .A2(n711), .ZN(n712) );
  NAND2_X1 U787 ( .A1(n725), .A2(n712), .ZN(n715) );
  AND2_X1 U788 ( .A1(n713), .A2(n715), .ZN(n714) );
  NAND2_X1 U789 ( .A1(n724), .A2(n714), .ZN(n719) );
  INV_X1 U790 ( .A(n715), .ZN(n717) );
  AND2_X1 U791 ( .A1(n728), .A2(n725), .ZN(n716) );
  OR2_X1 U792 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U793 ( .A1(n719), .A2(n718), .ZN(n736) );
  NOR2_X1 U794 ( .A1(G1971), .A2(G303), .ZN(n720) );
  NOR2_X1 U795 ( .A1(G1976), .A2(G288), .ZN(n977) );
  NOR2_X1 U796 ( .A1(n720), .A2(n977), .ZN(n722) );
  INV_X1 U797 ( .A(KEYINPUT33), .ZN(n721) );
  AND2_X1 U798 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U799 ( .A1(n724), .A2(n723), .ZN(n734) );
  XOR2_X1 U800 ( .A(G1981), .B(G305), .Z(n963) );
  AND2_X1 U801 ( .A1(n963), .A2(n725), .ZN(n732) );
  NAND2_X1 U802 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U803 ( .A(n974), .ZN(n726) );
  NOR2_X1 U804 ( .A1(KEYINPUT33), .A2(n515), .ZN(n730) );
  NAND2_X1 U805 ( .A1(n977), .A2(KEYINPUT33), .ZN(n727) );
  NOR2_X1 U806 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U807 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U808 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n738) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n970) );
  NAND2_X1 U812 ( .A1(n970), .A2(n751), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n738), .A2(n737), .ZN(n754) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n880), .ZN(n739) );
  XOR2_X1 U815 ( .A(KEYINPUT105), .B(n739), .Z(n994) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n740) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n901), .ZN(n1004) );
  NOR2_X1 U818 ( .A1(n740), .A2(n1004), .ZN(n741) );
  NOR2_X1 U819 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U820 ( .A1(n994), .A2(n743), .ZN(n744) );
  XNOR2_X1 U821 ( .A(KEYINPUT106), .B(n744), .ZN(n745) );
  XNOR2_X1 U822 ( .A(n745), .B(KEYINPUT39), .ZN(n747) );
  NAND2_X1 U823 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U824 ( .A(KEYINPUT107), .B(n748), .Z(n750) );
  NAND2_X1 U825 ( .A1(n749), .A2(n898), .ZN(n1011) );
  NAND2_X1 U826 ( .A1(n750), .A2(n1011), .ZN(n752) );
  NAND2_X1 U827 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U828 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n755), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U830 ( .A(G2427), .B(KEYINPUT108), .ZN(n765) );
  XOR2_X1 U831 ( .A(KEYINPUT109), .B(G2446), .Z(n757) );
  XNOR2_X1 U832 ( .A(G2435), .B(G2438), .ZN(n756) );
  XNOR2_X1 U833 ( .A(n757), .B(n756), .ZN(n761) );
  XOR2_X1 U834 ( .A(G2454), .B(G2430), .Z(n759) );
  XNOR2_X1 U835 ( .A(G1348), .B(G1341), .ZN(n758) );
  XNOR2_X1 U836 ( .A(n759), .B(n758), .ZN(n760) );
  XOR2_X1 U837 ( .A(n761), .B(n760), .Z(n763) );
  XNOR2_X1 U838 ( .A(G2451), .B(G2443), .ZN(n762) );
  XNOR2_X1 U839 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U840 ( .A(n765), .B(n764), .ZN(n766) );
  AND2_X1 U841 ( .A1(n766), .A2(G14), .ZN(G401) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U843 ( .A(G57), .ZN(G237) );
  INV_X1 U844 ( .A(G132), .ZN(G219) );
  INV_X1 U845 ( .A(G82), .ZN(G220) );
  INV_X1 U846 ( .A(n811), .ZN(G299) );
  XOR2_X1 U847 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n768) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U849 ( .A(n768), .B(n767), .ZN(G223) );
  INV_X1 U850 ( .A(G223), .ZN(n837) );
  NAND2_X1 U851 ( .A1(n837), .A2(G567), .ZN(n769) );
  XOR2_X1 U852 ( .A(KEYINPUT11), .B(n769), .Z(G234) );
  INV_X1 U853 ( .A(G860), .ZN(n777) );
  OR2_X1 U854 ( .A1(n983), .A2(n777), .ZN(G153) );
  XNOR2_X1 U855 ( .A(G171), .B(KEYINPUT69), .ZN(G301) );
  INV_X1 U856 ( .A(G868), .ZN(n774) );
  NAND2_X1 U857 ( .A1(n770), .A2(n774), .ZN(n772) );
  NAND2_X1 U858 ( .A1(G868), .A2(G301), .ZN(n771) );
  NAND2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U860 ( .A(KEYINPUT71), .B(n773), .Z(G284) );
  NOR2_X1 U861 ( .A1(G286), .A2(n774), .ZN(n776) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n776), .A2(n775), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n777), .A2(G559), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n778), .A2(n968), .ZN(n779) );
  XNOR2_X1 U866 ( .A(n779), .B(KEYINPUT16), .ZN(n780) );
  XOR2_X1 U867 ( .A(KEYINPUT73), .B(n780), .Z(G148) );
  NOR2_X1 U868 ( .A1(G868), .A2(n983), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n968), .A2(G868), .ZN(n781) );
  NOR2_X1 U870 ( .A1(G559), .A2(n781), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(G282) );
  XNOR2_X1 U872 ( .A(G2100), .B(KEYINPUT79), .ZN(n797) );
  XOR2_X1 U873 ( .A(KEYINPUT74), .B(KEYINPUT18), .Z(n785) );
  NAND2_X1 U874 ( .A1(G123), .A2(n886), .ZN(n784) );
  XNOR2_X1 U875 ( .A(n785), .B(n784), .ZN(n794) );
  NAND2_X1 U876 ( .A1(n885), .A2(G111), .ZN(n786) );
  XNOR2_X1 U877 ( .A(n786), .B(KEYINPUT76), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G99), .A2(n890), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U880 ( .A(n789), .B(KEYINPUT77), .ZN(n792) );
  NAND2_X1 U881 ( .A1(G135), .A2(n893), .ZN(n790) );
  XOR2_X1 U882 ( .A(KEYINPUT75), .B(n790), .Z(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n1000) );
  XNOR2_X1 U885 ( .A(n1000), .B(G2096), .ZN(n795) );
  XNOR2_X1 U886 ( .A(n795), .B(KEYINPUT78), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(G156) );
  NAND2_X1 U888 ( .A1(n968), .A2(G559), .ZN(n821) );
  XNOR2_X1 U889 ( .A(n983), .B(n821), .ZN(n798) );
  NOR2_X1 U890 ( .A1(n798), .A2(G860), .ZN(n809) );
  NAND2_X1 U891 ( .A1(G67), .A2(n799), .ZN(n802) );
  NAND2_X1 U892 ( .A1(G55), .A2(n800), .ZN(n801) );
  NAND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n808) );
  NAND2_X1 U894 ( .A1(G80), .A2(n803), .ZN(n806) );
  NAND2_X1 U895 ( .A1(G93), .A2(n804), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U897 ( .A1(n808), .A2(n807), .ZN(n817) );
  XNOR2_X1 U898 ( .A(n809), .B(n817), .ZN(G145) );
  NOR2_X1 U899 ( .A1(G868), .A2(n817), .ZN(n810) );
  XOR2_X1 U900 ( .A(n810), .B(KEYINPUT86), .Z(n824) );
  XOR2_X1 U901 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n813) );
  XNOR2_X1 U902 ( .A(n811), .B(KEYINPUT85), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n813), .B(n812), .ZN(n816) );
  XNOR2_X1 U904 ( .A(G166), .B(G305), .ZN(n814) );
  XNOR2_X1 U905 ( .A(n814), .B(G288), .ZN(n815) );
  XNOR2_X1 U906 ( .A(n816), .B(n815), .ZN(n819) );
  XNOR2_X1 U907 ( .A(G290), .B(n817), .ZN(n818) );
  XNOR2_X1 U908 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U909 ( .A(n820), .B(n983), .ZN(n905) );
  XNOR2_X1 U910 ( .A(n905), .B(n821), .ZN(n822) );
  NAND2_X1 U911 ( .A1(G868), .A2(n822), .ZN(n823) );
  NAND2_X1 U912 ( .A1(n824), .A2(n823), .ZN(G295) );
  NAND2_X1 U913 ( .A1(G2084), .A2(G2078), .ZN(n825) );
  XOR2_X1 U914 ( .A(KEYINPUT20), .B(n825), .Z(n826) );
  NAND2_X1 U915 ( .A1(G2090), .A2(n826), .ZN(n827) );
  XNOR2_X1 U916 ( .A(KEYINPUT21), .B(n827), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n828), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U918 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U919 ( .A1(G220), .A2(G219), .ZN(n829) );
  XOR2_X1 U920 ( .A(KEYINPUT22), .B(n829), .Z(n830) );
  NOR2_X1 U921 ( .A1(G218), .A2(n830), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G96), .A2(n831), .ZN(n841) );
  NAND2_X1 U923 ( .A1(n841), .A2(G2106), .ZN(n835) );
  NAND2_X1 U924 ( .A1(G120), .A2(G69), .ZN(n832) );
  NOR2_X1 U925 ( .A1(G237), .A2(n832), .ZN(n833) );
  NAND2_X1 U926 ( .A1(G108), .A2(n833), .ZN(n842) );
  NAND2_X1 U927 ( .A1(n842), .A2(G567), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n843) );
  NAND2_X1 U929 ( .A1(G483), .A2(G661), .ZN(n836) );
  NOR2_X1 U930 ( .A1(n843), .A2(n836), .ZN(n840) );
  NAND2_X1 U931 ( .A1(n840), .A2(G36), .ZN(G176) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U934 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(G188) );
  XOR2_X1 U937 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  XNOR2_X1 U938 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  NOR2_X1 U941 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  INV_X1 U943 ( .A(n843), .ZN(G319) );
  XOR2_X1 U944 ( .A(G2096), .B(G2100), .Z(n845) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2072), .Z(n847) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2090), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U950 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U951 ( .A(G2084), .B(G2078), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(G227) );
  XNOR2_X1 U953 ( .A(G1996), .B(KEYINPUT112), .ZN(n861) );
  XOR2_X1 U954 ( .A(G1976), .B(G1956), .Z(n853) );
  XNOR2_X1 U955 ( .A(G1991), .B(G1961), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U957 ( .A(G1981), .B(G1971), .Z(n855) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1966), .ZN(n854) );
  XNOR2_X1 U959 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U960 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U961 ( .A(G2474), .B(KEYINPUT41), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U964 ( .A1(n890), .A2(G100), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n862), .B(KEYINPUT114), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G112), .A2(n885), .ZN(n863) );
  XOR2_X1 U967 ( .A(KEYINPUT113), .B(n863), .Z(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n886), .A2(G124), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G136), .A2(n893), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U973 ( .A1(n870), .A2(n869), .ZN(G162) );
  XNOR2_X1 U974 ( .A(G164), .B(G162), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G118), .A2(n885), .ZN(n872) );
  NAND2_X1 U976 ( .A1(G130), .A2(n886), .ZN(n871) );
  NAND2_X1 U977 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n893), .A2(G142), .ZN(n874) );
  NAND2_X1 U979 ( .A1(G106), .A2(n890), .ZN(n873) );
  NAND2_X1 U980 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U981 ( .A(KEYINPUT45), .B(n875), .Z(n876) );
  NOR2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U983 ( .A(n879), .B(n878), .ZN(n884) );
  XNOR2_X1 U984 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n880), .B(n1000), .ZN(n881) );
  XNOR2_X1 U986 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n900) );
  NAND2_X1 U988 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n889), .B(KEYINPUT47), .ZN(n892) );
  NAND2_X1 U992 ( .A1(G103), .A2(n890), .ZN(n891) );
  NAND2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n896) );
  NAND2_X1 U994 ( .A1(G139), .A2(n893), .ZN(n894) );
  XNOR2_X1 U995 ( .A(KEYINPUT115), .B(n894), .ZN(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U997 ( .A(KEYINPUT116), .B(n897), .Z(n1007) );
  XNOR2_X1 U998 ( .A(n898), .B(n1007), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n901), .B(G160), .Z(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n904), .ZN(G395) );
  XOR2_X1 U1003 ( .A(n905), .B(G286), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G171), .B(n968), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n908), .ZN(n909) );
  XOR2_X1 U1007 ( .A(KEYINPUT117), .B(n909), .Z(G397) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n912), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(KEYINPUT119), .B(n914), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1018 ( .A(G20), .B(n917), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G19), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(G1981), .B(G6), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1023 ( .A(KEYINPUT59), .B(G1348), .Z(n922) );
  XNOR2_X1 U1024 ( .A(G4), .B(n922), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(KEYINPUT60), .B(n925), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G21), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(G5), .B(G1961), .ZN(n926) );
  NOR2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G22), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(G23), .B(G1976), .ZN(n930) );
  NOR2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n933) );
  XOR2_X1 U1034 ( .A(G1986), .B(G24), .Z(n932) );
  NAND2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1036 ( .A(KEYINPUT58), .B(n934), .ZN(n935) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(n937), .B(KEYINPUT61), .ZN(n939) );
  INV_X1 U1039 ( .A(G16), .ZN(n938) );
  NAND2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n962) );
  XNOR2_X1 U1041 ( .A(KEYINPUT54), .B(G34), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(n940), .B(KEYINPUT123), .ZN(n941) );
  XNOR2_X1 U1043 ( .A(G2084), .B(n941), .ZN(n959) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n957) );
  XNOR2_X1 U1045 ( .A(G1991), .B(G25), .ZN(n943) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n942) );
  NOR2_X1 U1047 ( .A1(n943), .A2(n942), .ZN(n950) );
  XOR2_X1 U1048 ( .A(G2067), .B(G26), .Z(n944) );
  NAND2_X1 U1049 ( .A1(n944), .A2(G28), .ZN(n948) );
  XOR2_X1 U1050 ( .A(G32), .B(n945), .Z(n946) );
  XNOR2_X1 U1051 ( .A(KEYINPUT122), .B(n946), .ZN(n947) );
  NOR2_X1 U1052 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1053 ( .A1(n950), .A2(n949), .ZN(n954) );
  XOR2_X1 U1054 ( .A(G27), .B(n951), .Z(n952) );
  XNOR2_X1 U1055 ( .A(KEYINPUT121), .B(n952), .ZN(n953) );
  NOR2_X1 U1056 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1058 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n989) );
  NOR2_X1 U1060 ( .A1(G29), .A2(KEYINPUT55), .ZN(n960) );
  NAND2_X1 U1061 ( .A1(n989), .A2(n960), .ZN(n961) );
  NAND2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n1022) );
  XOR2_X1 U1063 ( .A(KEYINPUT56), .B(G16), .Z(n988) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n964) );
  NAND2_X1 U1065 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1066 ( .A(n965), .B(KEYINPUT57), .ZN(n982) );
  XOR2_X1 U1067 ( .A(G171), .B(G1961), .Z(n967) );
  XNOR2_X1 U1068 ( .A(G299), .B(G1956), .ZN(n966) );
  NOR2_X1 U1069 ( .A1(n967), .A2(n966), .ZN(n972) );
  XOR2_X1 U1070 ( .A(G1348), .B(n968), .Z(n969) );
  NOR2_X1 U1071 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G166), .B(G1971), .ZN(n973) );
  XNOR2_X1 U1074 ( .A(n973), .B(KEYINPUT124), .ZN(n975) );
  NAND2_X1 U1075 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1076 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1077 ( .A(KEYINPUT125), .B(n978), .ZN(n979) );
  NOR2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(G1341), .B(n983), .ZN(n984) );
  NOR2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(KEYINPUT126), .B(n986), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n992) );
  INV_X1 U1084 ( .A(KEYINPUT55), .ZN(n1016) );
  OR2_X1 U1085 ( .A1(n1016), .A2(n989), .ZN(n990) );
  NAND2_X1 U1086 ( .A1(G11), .A2(n990), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n1020) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1090 ( .A(KEYINPUT120), .B(n995), .Z(n996) );
  XOR2_X1 U1091 ( .A(KEYINPUT51), .B(n996), .Z(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(G2084), .B(G160), .Z(n999) );
  NOR2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1014) );
  XOR2_X1 U1098 ( .A(G164), .B(G2078), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(G2072), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(n1010), .B(KEYINPUT50), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT52), .B(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(G29), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1023), .Z(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1024), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

