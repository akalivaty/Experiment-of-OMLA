//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n202), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G68), .Z(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n213), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n207), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n254), .A2(new_n256), .B1(new_n201), .B2(new_n207), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n248), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n247), .B(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n261), .B1(new_n206), .B2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n259), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  AND2_X1   g0069(.A1(G1), .A2(G13), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n274), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n206), .A2(new_n278), .B1(new_n270), .B2(new_n271), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(G226), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G179), .ZN(new_n281));
  AND2_X1   g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n282), .A2(new_n283), .A3(new_n213), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT66), .B1(new_n270), .B2(new_n271), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G222), .A2(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G223), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n286), .B(new_n291), .C1(G77), .C2(new_n287), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n280), .A2(new_n281), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n280), .A2(new_n292), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n268), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(G200), .B2(new_n294), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT9), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n263), .A2(new_n301), .A3(new_n267), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n263), .B2(new_n267), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n294), .A2(G200), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(KEYINPUT69), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n307), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n300), .C1(new_n302), .C2(new_n303), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n297), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n252), .B1(new_n206), .B2(G20), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n265), .A2(new_n259), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n252), .A2(new_n260), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n247), .ZN(new_n316));
  XNOR2_X1  g0116(.A(G58), .B(G68), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(G20), .B1(G159), .B2(new_n255), .ZN(new_n318));
  INV_X1    g0118(.A(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n207), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n321), .A2(G33), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT72), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT72), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n324), .A2(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n318), .B1(new_n333), .B2(new_n218), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n316), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(G20), .B1(new_n320), .B2(new_n322), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  OAI21_X1  g0138(.A(G68), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n323), .A2(new_n327), .A3(new_n207), .ZN(new_n340));
  OAI211_X1 g0140(.A(KEYINPUT16), .B(new_n318), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n315), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n278), .A2(new_n206), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n270), .A2(new_n271), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(G232), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n276), .ZN(new_n346));
  INV_X1    g0146(.A(G226), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G1698), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G223), .B2(G1698), .ZN(new_n349));
  INV_X1    g0149(.A(G87), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n349), .A2(new_n323), .B1(new_n319), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n346), .B1(new_n286), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G179), .ZN(new_n353));
  INV_X1    g0153(.A(new_n346), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n286), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G169), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT18), .B1(new_n342), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n318), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n331), .A2(new_n332), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n327), .B1(new_n287), .B2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n360), .B1(new_n363), .B2(G68), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n247), .B(new_n341), .C1(new_n364), .C2(KEYINPUT16), .ZN(new_n365));
  INV_X1    g0165(.A(new_n315), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT18), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n353), .A2(new_n357), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n354), .A2(new_n298), .A3(new_n355), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n352), .B2(G200), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n365), .A2(new_n372), .A3(new_n366), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n365), .A2(new_n372), .A3(KEYINPUT17), .A4(new_n366), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n359), .A2(new_n370), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n251), .B2(new_n202), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(KEYINPUT11), .A3(new_n248), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT12), .B1(new_n259), .B2(G68), .ZN(new_n382));
  OR3_X1    g0182(.A1(new_n259), .A2(KEYINPUT12), .A3(G68), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n260), .A2(new_n247), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n218), .B1(new_n206), .B2(G20), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n382), .A2(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT11), .B1(new_n380), .B2(new_n248), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n347), .A2(new_n289), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n231), .A2(G1698), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n320), .A2(new_n390), .A3(new_n322), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G97), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n286), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n279), .A2(G238), .B1(new_n272), .B2(new_n275), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n395), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g0199(.A(G200), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n283), .B1(new_n282), .B2(new_n213), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n270), .A2(KEYINPUT66), .A3(new_n271), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n393), .B2(new_n392), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n279), .A2(G238), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n276), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT13), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(G190), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n389), .A2(new_n400), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(G179), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT70), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT70), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n407), .A2(new_n414), .A3(G179), .A4(new_n408), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(G169), .B1(new_n398), .B2(new_n399), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT14), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(G169), .C1(new_n398), .C2(new_n399), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n389), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n411), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n350), .A2(KEYINPUT15), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT15), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G87), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n249), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n252), .A2(new_n256), .B1(new_n207), .B2(new_n202), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n247), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n384), .A2(new_n432), .B1(new_n202), .B2(new_n260), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n277), .B1(G244), .B2(new_n279), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n219), .A2(G1698), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(G232), .B2(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n287), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n286), .B(new_n438), .C1(G107), .C2(new_n287), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n434), .B1(new_n295), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n435), .A2(new_n281), .A3(new_n439), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(G200), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n434), .C1(new_n298), .C2(new_n440), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n311), .A2(new_n378), .A3(new_n423), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT5), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT74), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(G41), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n274), .A2(G1), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n273), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(G270), .A3(new_n344), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n272), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n459));
  OAI21_X1  g0259(.A(G303), .B1(new_n329), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G257), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n289), .ZN(new_n462));
  INV_X1    g0262(.A(G264), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G1698), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n320), .A2(new_n462), .A3(new_n322), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n466), .A2(new_n286), .A3(KEYINPUT79), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT79), .B1(new_n466), .B2(new_n286), .ZN(new_n468));
  OAI211_X1 g0268(.A(G190), .B(new_n458), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT75), .A2(G116), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT75), .A2(G116), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n259), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n319), .A2(G1), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n384), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(G20), .B1(G33), .B2(G283), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n319), .A2(G97), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n477), .A2(new_n478), .B1(new_n246), .B2(new_n213), .ZN(new_n479));
  OR2_X1    g0279(.A1(KEYINPUT75), .A2(G116), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT75), .A2(G116), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(G20), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT20), .B1(new_n479), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n476), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT79), .ZN(new_n487));
  INV_X1    g0287(.A(G303), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n320), .B2(new_n322), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n462), .A2(new_n464), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n287), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n491), .B2(new_n403), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n466), .A2(new_n286), .A3(KEYINPUT79), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n457), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G200), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n469), .B(new_n486), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(G179), .A3(new_n485), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n485), .A2(G169), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n494), .A2(new_n498), .A3(KEYINPUT21), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT21), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n458), .B1(new_n467), .B2(new_n468), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT20), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n477), .A2(new_n478), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n247), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n470), .A2(new_n471), .A3(new_n207), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n295), .B1(new_n508), .B2(new_n476), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n500), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n496), .B(new_n497), .C1(new_n499), .C2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT80), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n485), .A2(G179), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n501), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT21), .B1(new_n494), .B2(new_n498), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n501), .A2(new_n509), .A3(new_n500), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(KEYINPUT80), .A3(new_n496), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n473), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n265), .A2(new_n259), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n427), .B(KEYINPUT78), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR3_X1   g0325(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n526));
  INV_X1    g0326(.A(new_n393), .ZN(new_n527));
  AND2_X1   g0327(.A1(KEYINPUT76), .A2(KEYINPUT19), .ZN(new_n528));
  NOR2_X1   g0328(.A1(KEYINPUT76), .A2(KEYINPUT19), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n526), .B1(new_n530), .B2(new_n207), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n320), .A2(new_n322), .A3(new_n207), .A4(G68), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n533));
  OR2_X1    g0333(.A1(KEYINPUT76), .A2(KEYINPUT19), .ZN(new_n534));
  NAND2_X1  g0334(.A1(KEYINPUT76), .A2(KEYINPUT19), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n247), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n428), .A2(new_n260), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n538), .A2(KEYINPUT77), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT77), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n525), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G250), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n206), .B2(G45), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n272), .A2(new_n452), .B1(new_n344), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G238), .A2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n220), .B2(G1698), .ZN(new_n547));
  XNOR2_X1  g0347(.A(KEYINPUT75), .B(G116), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n547), .A2(new_n287), .B1(new_n548), .B2(G33), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n545), .B1(new_n549), .B2(new_n403), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n295), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n281), .B(new_n545), .C1(new_n549), .C2(new_n403), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n542), .A2(new_n554), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n556));
  INV_X1    g0356(.A(new_n249), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n548), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT81), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT81), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT24), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n320), .A2(new_n322), .A3(new_n207), .A4(G87), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n287), .A2(new_n568), .A3(new_n207), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n564), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n565), .B1(new_n564), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n247), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G107), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n260), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT25), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n523), .B2(G107), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n454), .A2(G264), .A3(new_n344), .ZN(new_n578));
  INV_X1    g0378(.A(G294), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n319), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(G250), .A2(G1698), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n461), .B2(G1698), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n580), .B1(new_n582), .B2(new_n287), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n578), .B(new_n456), .C1(new_n583), .C2(new_n403), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n495), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G190), .B2(new_n584), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n573), .A2(new_n577), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n550), .A2(new_n495), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G190), .B2(new_n550), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n523), .A2(G87), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n541), .C2(new_n540), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n555), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n454), .A2(new_n344), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n456), .B1(new_n593), .B2(new_n461), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT73), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n220), .A2(G1698), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n320), .A3(new_n322), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G250), .A2(G1698), .ZN(new_n601));
  NAND2_X1  g0401(.A1(KEYINPUT4), .A2(G244), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(G1698), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n287), .A2(new_n603), .B1(G33), .B2(G283), .ZN(new_n604));
  AOI211_X1 g0404(.A(new_n596), .B(new_n403), .C1(new_n600), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n600), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT73), .B1(new_n606), .B2(new_n286), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n281), .B(new_n595), .C1(new_n605), .C2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n574), .B1(new_n361), .B2(new_n362), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n255), .A2(G77), .ZN(new_n610));
  NAND2_X1  g0410(.A1(KEYINPUT6), .A2(G97), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(G107), .ZN(new_n612));
  XNOR2_X1  g0412(.A(G97), .B(G107), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT6), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n610), .B1(new_n615), .B2(new_n207), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n247), .B1(new_n609), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n265), .A2(G97), .A3(new_n259), .A4(new_n521), .ZN(new_n618));
  INV_X1    g0418(.A(G97), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n260), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n403), .B1(new_n604), .B2(new_n600), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n295), .B1(new_n594), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n608), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n622), .B(KEYINPUT73), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n495), .B1(new_n625), .B2(new_n595), .ZN(new_n626));
  INV_X1    g0426(.A(new_n622), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n595), .A2(new_n627), .A3(G190), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(new_n618), .A3(new_n617), .A4(new_n620), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n624), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n580), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n461), .A2(G1698), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(G250), .B2(G1698), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n633), .B2(new_n323), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n286), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(G179), .A3(new_n456), .A4(new_n578), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT83), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT82), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n584), .A2(new_n639), .A3(G169), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n584), .B2(G169), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n638), .A2(new_n642), .B1(new_n573), .B2(new_n577), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n592), .A2(new_n630), .A3(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n448), .A2(new_n520), .A3(new_n644), .ZN(G372));
  NAND2_X1  g0445(.A1(new_n375), .A2(new_n376), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n413), .A2(new_n415), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n418), .A2(new_n420), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n422), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n443), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n410), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n646), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n359), .A2(new_n370), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n310), .B2(new_n308), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n297), .ZN(new_n656));
  INV_X1    g0456(.A(new_n555), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n555), .A2(new_n591), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n624), .ZN(new_n660));
  INV_X1    g0460(.A(new_n624), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(new_n555), .A3(KEYINPUT26), .A4(new_n591), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n657), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n573), .A2(new_n577), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n640), .A2(new_n641), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n636), .B(KEYINPUT83), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n518), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n555), .A2(new_n587), .A3(new_n591), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n621), .A2(new_n623), .ZN(new_n670));
  AND4_X1   g0470(.A1(new_n628), .A2(new_n618), .A3(new_n617), .A4(new_n620), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n595), .B1(new_n605), .B2(new_n607), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G200), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n670), .A2(new_n608), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n668), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n663), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n656), .B1(new_n447), .B2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  INV_X1    g0479(.A(G13), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n680), .A2(G1), .A3(G20), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(G213), .B1(new_n682), .B2(KEYINPUT27), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT27), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n681), .A2(KEYINPUT84), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT84), .B1(new_n681), .B2(new_n684), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G343), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n520), .B1(new_n486), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n518), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n486), .A2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n679), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT85), .ZN(new_n695));
  INV_X1    g0495(.A(new_n689), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n664), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n587), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n695), .B1(new_n698), .B2(new_n643), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n667), .A2(KEYINPUT85), .A3(new_n697), .A4(new_n587), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n667), .A2(new_n689), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n694), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n518), .A2(new_n696), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n699), .A2(new_n700), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n643), .A2(new_n689), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n706), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n210), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G1), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n526), .A2(new_n474), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(new_n216), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n676), .A2(new_n689), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n630), .A2(KEYINPUT87), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT87), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n624), .B(new_n723), .C1(new_n626), .C2(new_n629), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n668), .A2(new_n722), .A3(new_n669), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n696), .B1(new_n663), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n511), .A2(new_n512), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT80), .B1(new_n518), .B2(new_n496), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n669), .A2(new_n674), .A3(new_n667), .A4(new_n689), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g0534(.A(G179), .B(new_n545), .C1(new_n549), .C2(new_n403), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n578), .B1(new_n583), .B2(new_n403), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n492), .A2(new_n493), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n594), .A2(new_n622), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n737), .A2(new_n738), .A3(new_n458), .A4(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n550), .A2(new_n281), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n672), .A2(new_n501), .A3(new_n584), .A4(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n494), .A2(KEYINPUT30), .A3(new_n737), .A4(new_n739), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n746), .A2(new_n696), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n746), .A2(new_n696), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(G330), .B1(new_n734), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n729), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n719), .B1(new_n757), .B2(G1), .ZN(G364));
  NOR2_X1   g0558(.A1(new_n680), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n206), .B1(new_n759), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n714), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n713), .A2(new_n323), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n764), .A2(G355), .B1(new_n474), .B2(new_n713), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n713), .A2(new_n287), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G45), .B2(new_n216), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n244), .A2(new_n274), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT89), .Z(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n213), .B1(G20), .B2(new_n295), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n763), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n773), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n207), .A2(G179), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G190), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT32), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(G20), .A2(G179), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n298), .A3(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n298), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n781), .B1(new_n218), .B2(new_n784), .C1(new_n787), .C2(new_n261), .ZN(new_n788));
  OR3_X1    g0588(.A1(new_n779), .A2(KEYINPUT32), .A3(new_n780), .ZN(new_n789));
  INV_X1    g0589(.A(G58), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n495), .A2(G190), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n782), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n783), .A2(new_n778), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n789), .B1(new_n790), .B2(new_n793), .C1(new_n202), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n791), .A2(G20), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT91), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n796), .A2(new_n797), .A3(new_n782), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(new_n796), .B2(new_n782), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n788), .B(new_n795), .C1(G97), .C2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n777), .A2(new_n298), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G107), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n805), .B(new_n287), .C1(new_n350), .C2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT90), .ZN(new_n808));
  INV_X1    g0608(.A(new_n779), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n809), .A2(G329), .B1(new_n792), .B2(G322), .ZN(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n810), .B(new_n323), .C1(new_n811), .C2(new_n794), .ZN(new_n812));
  INV_X1    g0612(.A(G326), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n787), .A2(new_n813), .B1(new_n806), .B2(new_n488), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT33), .B(G317), .Z(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n784), .A2(new_n815), .B1(new_n803), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n812), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n801), .A2(G294), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n802), .A2(new_n808), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n690), .A2(new_n693), .ZN(new_n821));
  INV_X1    g0621(.A(new_n772), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n775), .B1(new_n776), .B2(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n821), .A2(G330), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT88), .ZN(new_n825));
  INV_X1    g0625(.A(new_n694), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n763), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n823), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT92), .ZN(G396));
  OAI21_X1  g0629(.A(new_n445), .B1(new_n434), .B2(new_n689), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n443), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n650), .A2(new_n689), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n720), .B(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n755), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n762), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n838), .B2(KEYINPUT95), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(KEYINPUT95), .B2(new_n838), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n773), .A2(new_n770), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT93), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(G77), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n803), .A2(new_n350), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n787), .A2(new_n488), .B1(new_n806), .B2(new_n574), .ZN(new_n845));
  INV_X1    g0645(.A(new_n784), .ZN(new_n846));
  XNOR2_X1  g0646(.A(KEYINPUT94), .B(G283), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n848), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n793), .A2(new_n579), .B1(new_n779), .B2(new_n811), .ZN(new_n850));
  INV_X1    g0650(.A(new_n794), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n287), .B(new_n850), .C1(new_n548), .C2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n849), .B(new_n852), .C1(new_n619), .C2(new_n800), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n851), .A2(G159), .B1(G143), .B2(new_n792), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n854), .B1(new_n254), .B2(new_n784), .C1(new_n855), .C2(new_n787), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT34), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n287), .B1(new_n779), .B2(new_n859), .C1(new_n261), .C2(new_n806), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G68), .B2(new_n804), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n858), .B(new_n861), .C1(new_n790), .C2(new_n800), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n856), .A2(new_n857), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n853), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n763), .B(new_n843), .C1(new_n864), .C2(new_n773), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n771), .B2(new_n834), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n840), .A2(new_n866), .ZN(G384));
  NOR2_X1   g0667(.A1(new_n759), .A2(new_n206), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n341), .A2(new_n248), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n337), .A2(new_n327), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n870), .B(G68), .C1(new_n338), .C2(new_n337), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT16), .B1(new_n871), .B2(new_n318), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n366), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n688), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n377), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n369), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n874), .A3(new_n373), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n367), .A2(new_n369), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n367), .A2(new_n688), .ZN(new_n881));
  XNOR2_X1  g0681(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n373), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n876), .A2(new_n884), .A3(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n422), .A2(new_n696), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n649), .A2(new_n410), .A3(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n422), .B(new_n696), .C1(new_n421), .C2(new_n411), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n696), .B(new_n833), .C1(new_n663), .C2(new_n675), .ZN(new_n894));
  INV_X1    g0694(.A(new_n832), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n889), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n688), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n653), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n649), .A2(new_n696), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n884), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n876), .B2(new_n884), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n881), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n377), .A2(KEYINPUT98), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n880), .A2(new_n881), .A3(new_n373), .ZN(new_n907));
  INV_X1    g0707(.A(new_n882), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n883), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT98), .B1(new_n377), .B2(new_n905), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n886), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n888), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n904), .B1(new_n914), .B2(new_n903), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n899), .B1(new_n900), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n448), .B1(new_n721), .B2(new_n728), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n656), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n916), .B(new_n918), .Z(new_n919));
  AOI21_X1  g0719(.A(new_n749), .B1(new_n746), .B2(new_n696), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n689), .A2(new_n752), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n746), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT99), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT99), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n746), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n920), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n520), .A2(new_n644), .A3(new_n689), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n833), .B1(new_n891), .B2(new_n892), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(KEYINPUT40), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n914), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n901), .A2(new_n902), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n746), .A2(new_n924), .A3(new_n921), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n924), .B1(new_n746), .B2(new_n921), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n935), .A2(new_n936), .B1(new_n747), .B2(new_n749), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n929), .B1(new_n734), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n933), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n928), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n447), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n679), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n940), .B2(new_n942), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n868), .B1(new_n919), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n919), .B2(new_n944), .ZN(new_n946));
  INV_X1    g0746(.A(new_n615), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n474), .B(new_n215), .C1(new_n947), .C2(KEYINPUT35), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(KEYINPUT35), .B2(new_n947), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n202), .B(new_n216), .C1(G58), .C2(G68), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT96), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n951), .A2(new_n952), .B1(new_n261), .B2(G68), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n952), .B2(new_n951), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n680), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n946), .A2(new_n950), .A3(new_n955), .ZN(G367));
  NAND2_X1  g0756(.A1(new_n621), .A2(new_n696), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n722), .A2(new_n724), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n661), .A2(new_n696), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n711), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT45), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n710), .B2(new_n960), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT44), .B1(new_n710), .B2(new_n960), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n960), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n705), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n701), .B(new_n703), .C1(new_n518), .C2(new_n696), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT102), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n708), .B(new_n970), .C1(new_n694), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n708), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(new_n826), .A3(KEYINPUT102), .ZN(new_n974));
  AND4_X1   g0774(.A1(new_n729), .A2(new_n755), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n965), .B(new_n706), .C1(new_n966), .C2(new_n967), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n969), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT103), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n969), .A2(new_n975), .A3(KEYINPUT103), .A4(new_n976), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n756), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n714), .B(KEYINPUT41), .Z(new_n982));
  OAI21_X1  g0782(.A(new_n760), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n960), .B(KEYINPUT101), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n705), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT100), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n590), .B1(new_n540), .B2(new_n541), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n696), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n555), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n555), .A2(new_n989), .A3(new_n591), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT100), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n705), .A2(new_n985), .A3(new_n994), .ZN(new_n995));
  AND4_X1   g0795(.A1(new_n984), .A2(new_n987), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n987), .A2(new_n995), .B1(new_n984), .B2(new_n993), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n960), .A2(new_n708), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT42), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n661), .B1(new_n985), .B2(new_n643), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n696), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n998), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n983), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n774), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n713), .B2(new_n427), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n766), .A2(new_n237), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n763), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n787), .A2(new_n811), .B1(new_n803), .B2(new_n619), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G294), .B2(new_n846), .ZN(new_n1012));
  INV_X1    g0812(.A(G317), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n794), .A2(new_n847), .B1(new_n779), .B2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n287), .B(new_n1014), .C1(G303), .C2(new_n792), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n801), .A2(G107), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT46), .B1(new_n806), .B2(new_n474), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n548), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT46), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1017), .B1(new_n1019), .B2(new_n806), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .A4(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n779), .A2(new_n855), .B1(new_n794), .B2(new_n261), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n323), .B(new_n1022), .C1(G150), .C2(new_n792), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n801), .A2(G68), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n806), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G58), .A2(new_n1025), .B1(new_n846), .B2(G159), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n803), .A2(new_n202), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G143), .B2(new_n786), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1021), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT104), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT47), .Z(new_n1032));
  OAI221_X1 g0832(.A(new_n1010), .B1(new_n822), .B2(new_n992), .C1(new_n1032), .C2(new_n776), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1006), .A2(new_n1033), .ZN(G387));
  NOR2_X1   g0834(.A1(new_n975), .A2(new_n715), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n974), .A2(new_n972), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n757), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n761), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n764), .A2(new_n717), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(G107), .B2(new_n210), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n234), .A2(new_n274), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n766), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n252), .A2(G50), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT50), .ZN(new_n1044));
  AOI211_X1 g0844(.A(G45), .B(new_n717), .C1(G68), .C2(G77), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1040), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n762), .B1(new_n1047), .B2(new_n1007), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n323), .B1(new_n779), .B2(new_n813), .C1(new_n1018), .C2(new_n803), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n851), .A2(G303), .B1(G317), .B2(new_n792), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT105), .B(G322), .Z(new_n1051));
  OAI221_X1 g0851(.A(new_n1050), .B1(new_n811), .B2(new_n784), .C1(new_n787), .C2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT106), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1054), .A2(KEYINPUT48), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(KEYINPUT48), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n800), .A2(new_n847), .B1(new_n579), .B2(new_n806), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1049), .B1(new_n1058), .B2(KEYINPUT49), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(KEYINPUT49), .B2(new_n1058), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n787), .A2(new_n780), .B1(new_n806), .B2(new_n202), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n803), .A2(new_n619), .B1(new_n784), .B2(new_n252), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n801), .A2(new_n524), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n323), .B1(new_n851), .B2(G68), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n809), .A2(G150), .B1(new_n792), .B2(G50), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1060), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1048), .B1(new_n1068), .B2(new_n773), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n704), .B2(new_n822), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1037), .A2(new_n1038), .A3(new_n1070), .ZN(G393));
  AOI21_X1  g0871(.A(new_n715), .B1(new_n979), .B2(new_n980), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT107), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n969), .A2(new_n1073), .A3(new_n976), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1073), .B2(new_n976), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1072), .B1(new_n975), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n985), .A2(new_n822), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1042), .A2(new_n241), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n774), .B1(new_n619), .B2(new_n210), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n323), .B1(new_n794), .B2(new_n579), .C1(new_n1051), .C2(new_n779), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n805), .B1(new_n488), .B2(new_n784), .C1(new_n806), .C2(new_n847), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(new_n548), .C2(new_n801), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n786), .A2(G317), .B1(G311), .B2(new_n792), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT52), .Z(new_n1084));
  AOI22_X1  g0884(.A1(new_n786), .A2(G150), .B1(G159), .B2(new_n792), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT51), .Z(new_n1086));
  AOI21_X1  g0886(.A(new_n844), .B1(G50), .B2(new_n846), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n218), .B2(new_n806), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n800), .A2(new_n202), .ZN(new_n1089));
  INV_X1    g0889(.A(G143), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n287), .B1(new_n779), .B2(new_n1090), .C1(new_n252), .C2(new_n794), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1082), .A2(new_n1084), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n762), .B1(new_n1078), .B2(new_n1079), .C1(new_n1093), .C2(new_n776), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1077), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1075), .B2(new_n761), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1076), .A2(new_n1096), .ZN(G390));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n784), .A2(new_n855), .B1(new_n794), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n801), .B2(G159), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT110), .Z(new_n1101));
  NOR2_X1   g0901(.A1(new_n806), .A2(new_n254), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n793), .A2(new_n859), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n323), .B(new_n1104), .C1(G125), .C2(new_n809), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G128), .A2(new_n786), .B1(new_n804), .B2(G50), .ZN(new_n1106));
  AND4_X1   g0906(.A1(new_n1101), .A2(new_n1103), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n851), .A2(G97), .B1(G116), .B2(new_n792), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1108), .B(new_n323), .C1(new_n579), .C2(new_n779), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n787), .A2(new_n816), .B1(new_n574), .B2(new_n784), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n218), .A2(new_n803), .B1(new_n806), .B2(new_n350), .ZN(new_n1111));
  NOR4_X1   g0911(.A1(new_n1089), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n773), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n842), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n763), .B1(new_n1114), .B2(new_n252), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT111), .Z(new_n1117));
  INV_X1    g0917(.A(new_n915), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n771), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT112), .Z(new_n1121));
  INV_X1    g0921(.A(new_n900), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n895), .B1(new_n726), .B2(new_n831), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n893), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n914), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n676), .A2(new_n689), .A3(new_n834), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n832), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n900), .B1(new_n1127), .B2(new_n893), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1125), .B1(new_n915), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n928), .A2(G330), .A3(new_n929), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT108), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n928), .A2(KEYINPUT108), .A3(G330), .A4(new_n929), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n927), .A2(new_n753), .A3(new_n750), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1136), .A2(G330), .A3(new_n834), .A4(new_n893), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1135), .B1(new_n1129), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1121), .B1(new_n761), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1124), .B1(new_n755), .B2(new_n833), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1137), .A2(new_n1123), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n928), .A2(G330), .A3(new_n834), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1124), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1143), .A2(new_n1127), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n941), .A2(new_n679), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n448), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n917), .A2(new_n1149), .A3(new_n656), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n715), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT109), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1154), .B(new_n1135), .C1(new_n1129), .C2(new_n1138), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1153), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1141), .B1(new_n1156), .B2(new_n1157), .ZN(G378));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n268), .A2(new_n688), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n311), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n311), .A2(new_n1161), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1160), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n311), .A2(new_n1161), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1162), .A3(new_n1159), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1167), .A3(new_n1119), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n762), .B1(G50), .B2(new_n841), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n287), .A2(G41), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G50), .B(new_n1170), .C1(new_n319), .C2(new_n273), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1170), .B1(new_n816), .B2(new_n779), .C1(new_n793), .C2(new_n574), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n524), .B2(new_n851), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1025), .A2(G77), .B1(new_n804), .B2(G58), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G116), .A2(new_n786), .B1(new_n846), .B2(G97), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1173), .A2(new_n1024), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1171), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n792), .A2(G128), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n855), .B2(new_n794), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G132), .B2(new_n846), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1098), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n786), .A2(G125), .B1(new_n1025), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(new_n1183), .C1(new_n254), .C2(new_n800), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n804), .A2(G159), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1178), .B1(new_n1177), .B2(new_n1176), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1169), .B1(new_n1190), .B2(new_n773), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1168), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT113), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT114), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1165), .A2(new_n1167), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n939), .A2(G330), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n930), .B1(new_n888), .B2(new_n913), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n928), .B(new_n929), .C1(new_n901), .C2(new_n902), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n679), .B1(new_n1200), .B2(new_n933), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n932), .A3(new_n1195), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n916), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT117), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1203), .B(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1201), .A2(new_n932), .A3(new_n1195), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1195), .B1(new_n1201), .B2(new_n932), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT115), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT115), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1199), .A2(new_n1209), .A3(new_n1202), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n916), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT116), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT116), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1214), .B(new_n916), .C1(new_n1208), .C2(new_n1210), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1205), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1193), .B1(new_n1216), .B2(new_n761), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1150), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1155), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT57), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1212), .B1(new_n1207), .B2(new_n1206), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1203), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(KEYINPUT57), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n714), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1220), .B2(new_n1224), .ZN(G375));
  INV_X1    g1025(.A(new_n982), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1151), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n763), .B1(new_n1114), .B2(new_n218), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n770), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n803), .A2(new_n202), .B1(new_n784), .B2(new_n1018), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n323), .B1(new_n574), .B2(new_n794), .C1(new_n793), .C2(new_n816), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(G294), .C2(new_n786), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n806), .A2(new_n619), .B1(new_n779), .B2(new_n488), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT118), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1064), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n287), .B1(new_n803), .B2(new_n790), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT119), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n793), .A2(new_n855), .B1(new_n794), .B2(new_n254), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G128), .B2(new_n809), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n806), .A2(new_n780), .B1(new_n784), .B2(new_n1098), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G132), .B2(new_n786), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(new_n261), .C2(new_n800), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1236), .B1(new_n1238), .B2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(KEYINPUT120), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(KEYINPUT120), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n773), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1229), .B1(new_n893), .B2(new_n1230), .C1(new_n1245), .C2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1147), .B2(new_n760), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1228), .A2(new_n1250), .ZN(G381));
  INV_X1    g1051(.A(G390), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1141), .A2(new_n1253), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  OR3_X1    g1056(.A1(new_n1256), .A2(G375), .A3(G387), .ZN(G407));
  INV_X1    g1057(.A(G375), .ZN(new_n1258));
  INV_X1    g1058(.A(G213), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(G343), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1254), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT121), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1261), .B(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(G213), .A3(G407), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT122), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1264), .B(new_n1265), .ZN(G409));
  NAND3_X1  g1066(.A1(new_n1216), .A2(new_n1226), .A3(new_n1219), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1193), .B1(new_n1222), .B2(new_n761), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1254), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G378), .B(new_n1217), .C1(new_n1220), .C2(new_n1224), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1260), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT60), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n715), .B1(new_n1274), .B2(new_n1227), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1147), .A2(KEYINPUT60), .A3(new_n1150), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(KEYINPUT123), .A3(new_n1276), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1281), .B2(new_n1250), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1283), .B(new_n1249), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1272), .A2(new_n1273), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1260), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1285), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1006), .A2(G390), .A3(new_n1033), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G390), .B1(new_n1006), .B2(new_n1033), .ZN(new_n1294));
  XOR2_X1   g1094(.A(G393), .B(G396), .Z(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1293), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(new_n1252), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1298), .B2(new_n1292), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1288), .A2(new_n1289), .A3(new_n1291), .A4(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1290), .A2(KEYINPUT124), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT124), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1303), .B(new_n1260), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1280), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT123), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1250), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1283), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1281), .A2(G384), .A3(new_n1250), .ZN(new_n1309));
  INV_X1    g1109(.A(G2897), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1273), .A2(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1308), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1311), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1302), .A2(new_n1304), .A3(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1301), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT125), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1296), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1298), .A2(new_n1295), .A3(new_n1292), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(new_n1320), .A3(KEYINPUT125), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1286), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1290), .A2(KEYINPUT62), .A3(new_n1285), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT61), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1322), .B1(new_n1326), .B2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(KEYINPUT126), .B1(new_n1316), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1303), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1290), .A2(KEYINPUT124), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1327), .A3(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1319), .A2(new_n1320), .A3(new_n1289), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1335), .B1(new_n1287), .B2(new_n1286), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1334), .A2(new_n1336), .A3(new_n1291), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT126), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1289), .B1(new_n1314), .B2(new_n1290), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1339), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1337), .B(new_n1338), .C1(new_n1340), .C2(new_n1322), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1331), .A2(new_n1341), .ZN(G405));
  INV_X1    g1142(.A(new_n1285), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(G375), .A2(new_n1254), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1343), .B1(new_n1344), .B2(new_n1271), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1345), .B1(new_n1300), .B2(KEYINPUT127), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1343), .A2(new_n1271), .A3(new_n1344), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1300), .A2(KEYINPUT127), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1348), .B(new_n1349), .ZN(G402));
endmodule


