//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT73), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT26), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n208), .B(new_n209), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT27), .B(G183gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT28), .A3(new_n219), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n214), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n219), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(new_n212), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G190gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT23), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n234), .B(new_n235), .C1(new_n236), .C2(KEYINPUT25), .ZN(new_n237));
  AND2_X1   g036(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n238), .A2(new_n219), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  OR2_X1    g038(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(G190gat), .A3(new_n230), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n239), .A2(new_n241), .A3(new_n236), .A4(new_n227), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n239), .A2(new_n241), .A3(new_n227), .A4(new_n235), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n225), .B1(new_n237), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n205), .B1(new_n246), .B2(KEYINPUT29), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT74), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(KEYINPUT74), .B(new_n205), .C1(new_n246), .C2(KEYINPUT29), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n243), .B1(new_n244), .B2(new_n242), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n222), .A2(new_n224), .ZN(new_n253));
  OAI22_X1  g052(.A1(new_n251), .A2(new_n252), .B1(new_n253), .B2(new_n214), .ZN(new_n254));
  INV_X1    g053(.A(new_n203), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n249), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(G218gat), .ZN(new_n259));
  INV_X1    g058(.A(G211gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT70), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G211gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n259), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT69), .B(KEYINPUT22), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n258), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n267), .B(new_n258), .C1(new_n264), .C2(new_n265), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(new_n272), .A3(new_n268), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT72), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n255), .B1(new_n254), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n246), .A2(new_n205), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n281), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n202), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n283), .B1(new_n278), .B2(new_n257), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT75), .A3(new_n288), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n289), .B1(new_n285), .B2(KEYINPUT37), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT38), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n271), .A2(new_n276), .A3(new_n273), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n276), .B1(new_n271), .B2(new_n273), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n249), .A2(new_n297), .A3(new_n250), .A4(new_n256), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n274), .B1(new_n281), .B2(new_n282), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT37), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n294), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n290), .B(new_n292), .C1(new_n293), .C2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n288), .B1(new_n291), .B2(new_n301), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n285), .A2(KEYINPUT37), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n294), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT76), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(G155gat), .A3(G162gat), .ZN(new_n311));
  INV_X1    g110(.A(G155gat), .ZN(new_n312));
  INV_X1    g111(.A(G162gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n309), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n308), .A2(KEYINPUT2), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G141gat), .ZN(new_n318));
  INV_X1    g117(.A(G141gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(G148gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n316), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n315), .A2(KEYINPUT77), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n317), .A2(G141gat), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n324), .A2(new_n325), .B1(KEYINPUT2), .B2(new_n308), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n311), .A3(new_n314), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  INV_X1    g129(.A(G113gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(G120gat), .ZN(new_n332));
  INV_X1    g131(.A(G120gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(G113gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT65), .ZN(new_n336));
  NAND2_X1  g135(.A1(G127gat), .A2(G134gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(G127gat), .A2(G134gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n333), .A2(G113gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n331), .A2(G120gat), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT1), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n339), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n337), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT65), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n314), .A2(new_n308), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n342), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n333), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n343), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n345), .A2(KEYINPUT67), .A3(new_n337), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n338), .B2(new_n339), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n358));
  NAND4_X1  g157(.A1(new_n354), .A2(new_n355), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n329), .A2(new_n348), .A3(new_n350), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT4), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n354), .A2(new_n362), .B1(new_n341), .B2(new_n347), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n322), .A2(new_n328), .B1(new_n326), .B2(new_n349), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n359), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n370), .B1(new_n364), .B2(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n326), .A2(new_n327), .A3(new_n323), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT77), .B1(new_n315), .B2(new_n321), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n350), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n369), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n368), .A2(new_n377), .A3(KEYINPUT5), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n363), .A2(new_n364), .A3(new_n380), .A4(new_n365), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n361), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n366), .A2(KEYINPUT78), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n377), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n375), .A2(new_n370), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n360), .ZN(new_n387));
  INV_X1    g186(.A(new_n369), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n375), .A2(new_n370), .A3(KEYINPUT79), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT5), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n379), .B1(new_n384), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n383), .A2(new_n381), .A3(new_n361), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n363), .B1(KEYINPUT3), .B2(new_n375), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n364), .A2(new_n371), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n388), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n397), .A2(KEYINPUT80), .A3(KEYINPUT5), .A4(new_n390), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n378), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT0), .ZN(new_n401));
  XNOR2_X1  g200(.A(G57gat), .B(G85gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  NOR2_X1   g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT6), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n392), .A2(new_n398), .ZN(new_n406));
  INV_X1    g205(.A(new_n378), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n403), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT84), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT6), .B1(new_n399), .B2(new_n403), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n399), .B2(new_n403), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n307), .A2(new_n405), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416));
  INV_X1    g215(.A(G228gat), .ZN(new_n417));
  INV_X1    g216(.A(G233gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n395), .A2(new_n280), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n274), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n269), .B2(new_n270), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n375), .B1(new_n422), .B2(KEYINPUT3), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n420), .B1(new_n295), .B2(new_n296), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(KEYINPUT81), .B(new_n420), .C1(new_n295), .C2(new_n296), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n271), .A2(new_n280), .A3(new_n273), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n371), .ZN(new_n431));
  AOI211_X1 g230(.A(new_n417), .B(new_n418), .C1(new_n431), .C2(new_n375), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n424), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G22gat), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n416), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G78gat), .B(G106gat), .Z(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT31), .B(G50gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n431), .A2(new_n375), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n419), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n427), .B2(new_n428), .ZN(new_n441));
  OAI21_X1  g240(.A(G22gat), .B1(new_n441), .B2(new_n424), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT81), .B1(new_n278), .B2(new_n420), .ZN(new_n443));
  INV_X1    g242(.A(new_n428), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n432), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n424), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n434), .A3(new_n446), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n435), .A2(new_n438), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n442), .A2(new_n447), .A3(KEYINPUT82), .A4(new_n438), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n290), .A2(new_n452), .A3(new_n292), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n291), .A2(new_n288), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n285), .A2(new_n289), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(KEYINPUT30), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n394), .A2(new_n395), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n369), .B1(new_n459), .B2(new_n367), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT39), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n388), .B1(new_n387), .B2(new_n389), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n461), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n403), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n403), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT40), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n410), .A2(new_n413), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n451), .B1(new_n458), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT85), .B1(new_n415), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n434), .B1(new_n445), .B2(new_n446), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n438), .B1(new_n474), .B2(KEYINPUT82), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n442), .A2(new_n447), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n449), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n410), .A2(new_n413), .A3(new_n470), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(new_n457), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n307), .A2(new_n405), .A3(new_n414), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n448), .A2(new_n450), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT83), .B1(new_n477), .B2(new_n449), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n411), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n405), .B1(new_n489), .B2(new_n404), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n458), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n254), .A2(new_n363), .ZN(new_n492));
  INV_X1    g291(.A(G227gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(new_n418), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n246), .A2(new_n370), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT32), .ZN(new_n497));
  XOR2_X1   g296(.A(G15gat), .B(G43gat), .Z(new_n498));
  XNOR2_X1  g297(.A(G71gat), .B(G99gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT33), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n492), .A2(new_n495), .ZN(new_n505));
  INV_X1    g304(.A(new_n494), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI211_X1 g306(.A(KEYINPUT34), .B(new_n494), .C1(new_n492), .C2(new_n495), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n497), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n502), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n500), .ZN(new_n514));
  INV_X1    g313(.A(new_n508), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n505), .A2(new_n506), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT34), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n497), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n509), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n512), .A2(KEYINPUT36), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n518), .A2(new_n519), .A3(new_n509), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n519), .B1(new_n518), .B2(new_n509), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n488), .A2(new_n491), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n484), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n523), .A2(new_n524), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n478), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n531));
  AND3_X1   g330(.A1(new_n530), .A2(new_n458), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n414), .A2(new_n405), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n490), .A2(new_n458), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n530), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n527), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT101), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT15), .ZN(new_n541));
  INV_X1    g340(.A(G43gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n543));
  XOR2_X1   g342(.A(G43gat), .B(G50gat), .Z(new_n544));
  OAI211_X1 g343(.A(new_n541), .B(new_n543), .C1(new_n544), .C2(KEYINPUT89), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  OR3_X1    g345(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n548));
  INV_X1    g347(.A(G29gat), .ZN(new_n549));
  INV_X1    g348(.A(G36gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(KEYINPUT88), .A2(G29gat), .A3(G36gat), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n546), .A2(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n544), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(KEYINPUT15), .A3(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT7), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  INV_X1    g364(.A(G92gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G99gat), .B(G106gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT95), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n561), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT41), .ZN(new_n573));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  OAI22_X1  g373(.A1(new_n559), .A2(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  OAI22_X1  g376(.A1(new_n572), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n574), .A2(new_n573), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(G57gat), .B(G64gat), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n593), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n594), .A2(new_n586), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G127gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G15gat), .B(G22gat), .ZN(new_n604));
  INV_X1    g403(.A(G1gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT16), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(G1gat), .B2(new_n604), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G8gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n599), .B2(new_n598), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n603), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n312), .ZN(new_n614));
  XOR2_X1   g413(.A(G183gat), .B(G211gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n585), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT91), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n610), .A2(new_n559), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n609), .B(KEYINPUT90), .Z(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n624), .B2(new_n561), .ZN(new_n625));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT18), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n610), .B(new_n559), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n626), .B(KEYINPUT13), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G113gat), .B(G141gat), .Z(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G169gat), .B(G197gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n629), .A2(new_n630), .A3(new_n633), .A4(new_n640), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT92), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT92), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n634), .A2(new_n645), .A3(new_n641), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n570), .A2(new_n598), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  OR3_X1    g448(.A1(new_n648), .A2(KEYINPUT98), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT98), .B1(new_n648), .B2(new_n649), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n570), .A2(new_n598), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(KEYINPUT97), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n570), .A2(new_n598), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT10), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT99), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT100), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n654), .A2(new_n660), .A3(new_n656), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n658), .B2(new_n660), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n662), .A2(new_n663), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n666), .ZN(new_n670));
  INV_X1    g469(.A(new_n663), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n661), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n621), .A2(new_n647), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n539), .A2(new_n540), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n540), .B1(new_n539), .B2(new_n674), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n490), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n605), .ZN(G1324gat));
  OR2_X1    g479(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  AND3_X1   g481(.A1(new_n681), .A2(new_n457), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(G8gat), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n681), .B2(new_n457), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT42), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(KEYINPUT42), .B2(new_n683), .ZN(G1325gat));
  AOI21_X1  g486(.A(G15gat), .B1(new_n681), .B2(new_n528), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n523), .A2(new_n524), .A3(new_n522), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT36), .B1(new_n512), .B2(new_n520), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n525), .A2(KEYINPUT102), .A3(new_n521), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT103), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G15gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT104), .Z(new_n698));
  AOI21_X1  g497(.A(new_n688), .B1(new_n681), .B2(new_n698), .ZN(G1326gat));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n681), .A2(new_n700), .A3(new_n488), .ZN(new_n701));
  INV_X1    g500(.A(new_n487), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n451), .A2(KEYINPUT83), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT105), .B1(new_n678), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  AOI21_X1  g507(.A(new_n585), .B1(new_n527), .B2(new_n538), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n647), .A2(new_n620), .A3(new_n673), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(G29gat), .A3(new_n490), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT45), .Z(new_n713));
  AOI22_X1  g512(.A1(new_n533), .A2(new_n532), .B1(new_n536), .B2(KEYINPUT35), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n694), .B1(new_n488), .B2(new_n491), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n457), .A2(new_n413), .A3(new_n410), .A4(new_n470), .ZN(new_n716));
  AND4_X1   g515(.A1(new_n481), .A2(new_n482), .A3(new_n451), .A4(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n481), .B1(new_n480), .B2(new_n482), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT106), .B(new_n715), .C1(new_n717), .C2(new_n718), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n714), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n585), .A2(KEYINPUT44), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n723), .A2(new_n725), .B1(new_n726), .B2(new_n709), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n710), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n490), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n729), .ZN(G1328gat));
  NOR3_X1   g529(.A1(new_n711), .A2(G36gat), .A3(new_n458), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT107), .B1(new_n728), .B2(new_n458), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G36gat), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n728), .A2(KEYINPUT107), .A3(new_n458), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n694), .ZN(new_n737));
  OAI21_X1  g536(.A(G43gat), .B1(new_n728), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n711), .A2(G43gat), .A3(new_n529), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n721), .A2(new_n722), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n725), .B1(new_n743), .B2(new_n538), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n709), .A2(new_n726), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n696), .B(new_n710), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n746), .A2(new_n747), .A3(G43gat), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n746), .B2(G43gat), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n748), .A2(new_n749), .A3(new_n739), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n742), .B1(new_n750), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  OAI21_X1  g551(.A(G50gat), .B1(new_n728), .B2(new_n451), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n711), .A2(G50gat), .A3(new_n704), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT109), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n752), .B(G50gat), .C1(new_n728), .C2(new_n704), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(KEYINPUT109), .B2(KEYINPUT48), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(G1331gat));
  NAND4_X1  g558(.A1(new_n647), .A2(new_n620), .A3(new_n585), .A4(new_n673), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n723), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n490), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  OR3_X1    g563(.A1(new_n723), .A2(KEYINPUT110), .A3(new_n760), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT110), .B1(new_n723), .B2(new_n760), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n457), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT49), .B(G64gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(G1333gat));
  NAND3_X1  g569(.A1(new_n765), .A2(new_n696), .A3(new_n766), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n529), .A2(G71gat), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n771), .A2(G71gat), .B1(new_n761), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g573(.A1(new_n765), .A2(new_n488), .A3(new_n766), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777));
  INV_X1    g576(.A(new_n722), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT106), .B1(new_n484), .B2(new_n715), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n538), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n704), .A2(new_n535), .B1(new_n690), .B2(new_n691), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n473), .B2(new_n483), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n584), .B1(new_n782), .B2(new_n714), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n780), .A2(new_n724), .B1(new_n783), .B2(KEYINPUT44), .ZN(new_n784));
  INV_X1    g583(.A(new_n620), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n647), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n673), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n777), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n727), .A2(KEYINPUT111), .A3(new_n788), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n790), .A2(new_n762), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n786), .A2(new_n585), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n723), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n794), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n762), .A2(new_n565), .A3(new_n673), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n792), .A2(new_n565), .B1(new_n799), .B2(new_n800), .ZN(G1336gat));
  NAND3_X1  g600(.A1(new_n790), .A2(new_n457), .A3(new_n791), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n787), .A2(G92gat), .A3(new_n458), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n802), .A2(G92gat), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  XOR2_X1   g604(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n798), .B2(new_n803), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n457), .B(new_n788), .C1(new_n744), .C2(new_n745), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G92gat), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n807), .B2(new_n810), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n804), .A2(new_n805), .B1(new_n811), .B2(new_n812), .ZN(G1337gat));
  NAND3_X1  g612(.A1(new_n790), .A2(new_n696), .A3(new_n791), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT114), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n790), .A2(new_n816), .A3(new_n791), .A4(new_n696), .ZN(new_n817));
  XOR2_X1   g616(.A(KEYINPUT115), .B(G99gat), .Z(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n798), .A2(new_n528), .A3(new_n673), .A4(new_n818), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1338gat));
  NOR3_X1   g621(.A1(new_n787), .A2(new_n451), .A3(G106gat), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT53), .B1(new_n798), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(G106gat), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n784), .A2(new_n451), .A3(new_n789), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n790), .A2(new_n488), .A3(new_n791), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n828), .A2(G106gat), .B1(new_n798), .B2(new_n823), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(G1339gat));
  INV_X1    g630(.A(new_n639), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n625), .A2(new_n626), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n631), .A2(new_n632), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT116), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(KEYINPUT116), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n643), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n658), .B2(new_n660), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n662), .A2(new_n668), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n666), .B1(new_n661), .B2(new_n839), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n841), .B2(new_n843), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n838), .B(new_n669), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n620), .B1(new_n846), .B2(new_n584), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n584), .B1(new_n838), .B2(new_n673), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n669), .B1(new_n844), .B2(new_n845), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n647), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n621), .A2(new_n673), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n647), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n762), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(new_n478), .A3(new_n529), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n856), .A2(new_n458), .ZN(new_n857));
  INV_X1    g656(.A(new_n647), .ZN(new_n858));
  AOI21_X1  g657(.A(G113gat), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n850), .A2(new_n847), .B1(new_n852), .B2(new_n647), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n488), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n490), .A2(new_n457), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n528), .A3(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n331), .A3(new_n647), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n859), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n860), .B1(new_n859), .B2(new_n865), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1340gat));
  NAND3_X1  g667(.A1(new_n857), .A2(new_n333), .A3(new_n673), .ZN(new_n869));
  OAI21_X1  g668(.A(G120gat), .B1(new_n864), .B2(new_n787), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(G1341gat));
  INV_X1    g673(.A(G127gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n864), .A2(new_n875), .A3(new_n785), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT119), .Z(new_n877));
  AOI21_X1  g676(.A(G127gat), .B1(new_n857), .B2(new_n620), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1342gat));
  INV_X1    g678(.A(G134gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n584), .A2(new_n458), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT120), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n856), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  OAI21_X1  g683(.A(G134gat), .B1(new_n864), .B2(new_n585), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G1343gat));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT57), .B1(new_n861), .B2(new_n704), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n854), .A2(new_n891), .A3(new_n478), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n737), .A2(new_n863), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n890), .A2(new_n892), .A3(new_n858), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G141gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n695), .A2(new_n478), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n855), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n898), .A2(new_n319), .A3(new_n458), .A4(new_n858), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n889), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n319), .B1(new_n895), .B2(KEYINPUT121), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n889), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n888), .B(new_n901), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n903), .B2(new_n902), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT122), .B1(new_n907), .B2(new_n900), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1344gat));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n855), .A2(new_n897), .A3(new_n457), .ZN(new_n911));
  AOI211_X1 g710(.A(new_n910), .B(G148gat), .C1(new_n911), .C2(new_n673), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n892), .A3(new_n894), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n913), .B2(new_n787), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT57), .B1(new_n861), .B2(new_n451), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n854), .A2(new_n891), .A3(new_n488), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n894), .A2(KEYINPUT59), .A3(new_n673), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n912), .B1(new_n919), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n913), .B2(new_n785), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n911), .A2(new_n312), .A3(new_n620), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n913), .B2(new_n585), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n898), .A2(new_n313), .A3(new_n882), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n762), .A2(new_n458), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n862), .A2(new_n528), .A3(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(new_n206), .A3(new_n647), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n854), .A2(new_n530), .A3(new_n927), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n858), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n932), .B2(new_n206), .ZN(G1348gat));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n207), .A3(new_n673), .ZN(new_n934));
  OAI21_X1  g733(.A(G176gat), .B1(new_n928), .B2(new_n787), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1349gat));
  OAI21_X1  g735(.A(G183gat), .B1(new_n928), .B2(new_n785), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n620), .A2(new_n223), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n930), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n937), .A2(KEYINPUT125), .A3(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n940), .A2(new_n942), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT124), .B1(new_n937), .B2(new_n939), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n928), .B2(new_n585), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n219), .A3(new_n584), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1351gat));
  INV_X1    g749(.A(new_n927), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n696), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n915), .A2(new_n916), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(G197gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n953), .A2(new_n954), .A3(new_n647), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n861), .A2(new_n897), .A3(new_n951), .ZN(new_n956));
  AOI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n858), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n955), .A2(new_n957), .ZN(G1352gat));
  INV_X1    g757(.A(G204gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n956), .A2(new_n959), .A3(new_n673), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT62), .Z(new_n961));
  OAI21_X1  g760(.A(G204gat), .B1(new_n953), .B2(new_n787), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1353gat));
  NAND4_X1  g762(.A1(new_n956), .A2(new_n261), .A3(new_n263), .A4(new_n620), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n915), .A2(new_n916), .A3(new_n620), .A4(new_n952), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(G211gat), .A3(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n964), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  OAI21_X1  g772(.A(G218gat), .B1(new_n953), .B2(new_n585), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n259), .A3(new_n584), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1355gat));
endmodule


