

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U546 ( .A1(n633), .A2(n849), .ZN(n615) );
  XOR2_X1 U547 ( .A(KEYINPUT77), .B(n534), .Z(n513) );
  XOR2_X2 U548 ( .A(KEYINPUT15), .B(n614), .Z(n849) );
  XNOR2_X2 U549 ( .A(KEYINPUT78), .B(n542), .ZN(G168) );
  INV_X1 U550 ( .A(n520), .ZN(n907) );
  XOR2_X1 U551 ( .A(G543), .B(KEYINPUT0), .Z(n568) );
  BUF_X1 U552 ( .A(n645), .Z(n663) );
  XNOR2_X1 U553 ( .A(n679), .B(KEYINPUT32), .ZN(n680) );
  NAND2_X1 U554 ( .A1(n697), .A2(n590), .ZN(n645) );
  NAND2_X1 U555 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U556 ( .A1(n745), .A2(n744), .ZN(n747) );
  NOR2_X1 U557 ( .A1(n526), .A2(n525), .ZN(G164) );
  NOR2_X1 U558 ( .A1(n738), .A2(n737), .ZN(n514) );
  XOR2_X1 U559 ( .A(KEYINPUT93), .B(n621), .Z(n515) );
  NOR2_X1 U560 ( .A1(n818), .A2(n639), .ZN(n632) );
  INV_X1 U561 ( .A(n645), .ZN(n629) );
  INV_X1 U562 ( .A(KEYINPUT97), .ZN(n682) );
  XNOR2_X1 U563 ( .A(n683), .B(n682), .ZN(n736) );
  XNOR2_X1 U564 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n519) );
  INV_X1 U565 ( .A(KEYINPUT100), .ZN(n746) );
  NOR2_X1 U566 ( .A1(G543), .A2(G651), .ZN(n807) );
  XNOR2_X1 U567 ( .A(KEYINPUT64), .B(n533), .ZN(n804) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n536), .Z(n803) );
  AND2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n902) );
  NAND2_X1 U570 ( .A1(G114), .A2(n902), .ZN(n517) );
  INV_X1 U571 ( .A(G2105), .ZN(n522) );
  AND2_X1 U572 ( .A1(n522), .A2(G2104), .ZN(n906) );
  NAND2_X1 U573 ( .A1(G102), .A2(n906), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n517), .A2(n516), .ZN(n526) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  XNOR2_X1 U576 ( .A(n519), .B(n518), .ZN(n543) );
  INV_X1 U577 ( .A(n543), .ZN(n520) );
  NAND2_X1 U578 ( .A1(G138), .A2(n907), .ZN(n521) );
  XNOR2_X1 U579 ( .A(n521), .B(KEYINPUT88), .ZN(n524) );
  NOR2_X1 U580 ( .A1(G2104), .A2(n522), .ZN(n903) );
  NAND2_X1 U581 ( .A1(n903), .A2(G126), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U583 ( .A(G651), .B(KEYINPUT67), .ZN(n535) );
  NOR2_X1 U584 ( .A1(n568), .A2(n535), .ZN(n808) );
  NAND2_X1 U585 ( .A1(G76), .A2(n808), .ZN(n530) );
  XOR2_X1 U586 ( .A(KEYINPUT4), .B(KEYINPUT75), .Z(n528) );
  NAND2_X1 U587 ( .A1(G89), .A2(n807), .ZN(n527) );
  XNOR2_X1 U588 ( .A(n528), .B(n527), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U590 ( .A(n531), .B(KEYINPUT76), .ZN(n532) );
  XNOR2_X1 U591 ( .A(KEYINPUT5), .B(n532), .ZN(n540) );
  NOR2_X1 U592 ( .A1(G651), .A2(n568), .ZN(n533) );
  NAND2_X1 U593 ( .A1(G51), .A2(n804), .ZN(n534) );
  NOR2_X1 U594 ( .A1(G543), .A2(n535), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n803), .A2(G63), .ZN(n537) );
  NAND2_X1 U596 ( .A1(n513), .A2(n537), .ZN(n538) );
  XOR2_X1 U597 ( .A(KEYINPUT6), .B(n538), .Z(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n541), .B(KEYINPUT7), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G137), .A2(n543), .ZN(n545) );
  NAND2_X1 U601 ( .A1(G113), .A2(n902), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n547) );
  INV_X1 U603 ( .A(KEYINPUT66), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n547), .B(n546), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n903), .A2(G125), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G101), .A2(n906), .ZN(n550) );
  XNOR2_X1 U608 ( .A(KEYINPUT23), .B(n550), .ZN(n551) );
  NOR2_X2 U609 ( .A1(n552), .A2(n551), .ZN(G160) );
  NAND2_X1 U610 ( .A1(n803), .A2(G64), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G52), .A2(n804), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U613 ( .A(KEYINPUT69), .B(n555), .Z(n560) );
  NAND2_X1 U614 ( .A1(G90), .A2(n807), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G77), .A2(n808), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U618 ( .A1(n560), .A2(n559), .ZN(G171) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  NAND2_X1 U620 ( .A1(G88), .A2(n807), .ZN(n562) );
  NAND2_X1 U621 ( .A1(G75), .A2(n808), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n803), .A2(G62), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G50), .A2(n804), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U626 ( .A1(n566), .A2(n565), .ZN(G166) );
  INV_X1 U627 ( .A(G166), .ZN(G303) );
  XOR2_X1 U628 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U629 ( .A1(n804), .A2(G49), .ZN(n567) );
  XNOR2_X1 U630 ( .A(n567), .B(KEYINPUT82), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G87), .A2(n568), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U634 ( .A1(n803), .A2(n571), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n573), .A2(n572), .ZN(G288) );
  XOR2_X1 U636 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n575) );
  NAND2_X1 U637 ( .A1(G73), .A2(n808), .ZN(n574) );
  XNOR2_X1 U638 ( .A(n575), .B(n574), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G86), .A2(n807), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G61), .A2(n803), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT83), .B(n578), .Z(n579) );
  NOR2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G48), .A2(n804), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(G305) );
  NAND2_X1 U646 ( .A1(n808), .A2(G72), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n807), .A2(G85), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT68), .B(n585), .Z(n589) );
  NAND2_X1 U650 ( .A1(n804), .A2(G47), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n803), .A2(G60), .ZN(n586) );
  AND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(G290) );
  NOR2_X1 U654 ( .A1(G164), .A2(G1384), .ZN(n697) );
  NAND2_X1 U655 ( .A1(G160), .A2(G40), .ZN(n696) );
  XOR2_X1 U656 ( .A(KEYINPUT90), .B(n696), .Z(n590) );
  NOR2_X1 U657 ( .A1(G2084), .A2(n645), .ZN(n646) );
  NAND2_X1 U658 ( .A1(G8), .A2(n646), .ZN(n662) );
  NAND2_X1 U659 ( .A1(G1961), .A2(n663), .ZN(n592) );
  XOR2_X1 U660 ( .A(G2078), .B(KEYINPUT25), .Z(n1009) );
  NAND2_X1 U661 ( .A1(n629), .A2(n1009), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n652) );
  OR2_X1 U663 ( .A1(G301), .A2(n652), .ZN(n669) );
  AND2_X1 U664 ( .A1(n629), .A2(G1996), .ZN(n593) );
  XOR2_X1 U665 ( .A(n593), .B(KEYINPUT26), .Z(n634) );
  AND2_X1 U666 ( .A1(n663), .A2(G1341), .ZN(n606) );
  NAND2_X1 U667 ( .A1(G81), .A2(n807), .ZN(n594) );
  XNOR2_X1 U668 ( .A(n594), .B(KEYINPUT12), .ZN(n595) );
  XNOR2_X1 U669 ( .A(n595), .B(KEYINPUT70), .ZN(n597) );
  NAND2_X1 U670 ( .A1(G68), .A2(n808), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U672 ( .A(KEYINPUT13), .B(n598), .ZN(n605) );
  NAND2_X1 U673 ( .A1(n804), .A2(G43), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT71), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n803), .A2(G56), .ZN(n600) );
  XNOR2_X1 U676 ( .A(KEYINPUT14), .B(n600), .ZN(n601) );
  INV_X1 U677 ( .A(n601), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n982) );
  NOR2_X1 U680 ( .A1(n606), .A2(n982), .ZN(n633) );
  NAND2_X1 U681 ( .A1(G92), .A2(n807), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G66), .A2(n803), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n613) );
  NAND2_X1 U684 ( .A1(G79), .A2(n808), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G54), .A2(n804), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U687 ( .A(KEYINPUT73), .B(n611), .Z(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n634), .A2(n615), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n616), .B(KEYINPUT92), .ZN(n620) );
  NOR2_X1 U691 ( .A1(n629), .A2(G1348), .ZN(n618) );
  NOR2_X1 U692 ( .A1(G2067), .A2(n663), .ZN(n617) );
  NOR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n803), .A2(G65), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G53), .A2(n804), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G91), .A2(n807), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G78), .A2(n808), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n818) );
  NAND2_X1 U702 ( .A1(n629), .A2(G2072), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT27), .ZN(n631) );
  INV_X1 U704 ( .A(G1956), .ZN(n951) );
  NOR2_X1 U705 ( .A1(n951), .A2(n629), .ZN(n630) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n639) );
  XOR2_X1 U707 ( .A(n632), .B(KEYINPUT28), .Z(n637) );
  AND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  OR2_X1 U709 ( .A1(n635), .A2(n849), .ZN(n636) );
  AND2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n515), .A2(n638), .ZN(n643) );
  INV_X1 U712 ( .A(KEYINPUT28), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n818), .A2(n639), .ZN(n640) );
  OR2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n644), .B(KEYINPUT29), .ZN(n671) );
  NAND2_X1 U717 ( .A1(n669), .A2(n671), .ZN(n658) );
  INV_X1 U718 ( .A(KEYINPUT31), .ZN(n657) );
  NAND2_X1 U719 ( .A1(G8), .A2(n645), .ZN(n737) );
  NOR2_X1 U720 ( .A1(G1966), .A2(n737), .ZN(n659) );
  INV_X1 U721 ( .A(n646), .ZN(n647) );
  NAND2_X1 U722 ( .A1(G8), .A2(n647), .ZN(n648) );
  OR2_X1 U723 ( .A1(n659), .A2(n648), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n649), .B(KEYINPUT30), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(KEYINPUT94), .ZN(n651) );
  NOR2_X1 U726 ( .A1(n651), .A2(G168), .ZN(n655) );
  NAND2_X1 U727 ( .A1(G301), .A2(n652), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT95), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n657), .B(n656), .ZN(n673) );
  AND2_X1 U731 ( .A1(n658), .A2(n673), .ZN(n660) );
  NOR2_X1 U732 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n681) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n737), .ZN(n665) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n663), .ZN(n664) );
  NOR2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n666), .B(KEYINPUT96), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n667), .A2(G303), .ZN(n672) );
  INV_X1 U739 ( .A(n672), .ZN(n668) );
  OR2_X1 U740 ( .A1(n668), .A2(G286), .ZN(n674) );
  AND2_X1 U741 ( .A1(n669), .A2(n674), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n678), .A2(G8), .ZN(n679) );
  NOR2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n692) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n692), .A2(n684), .ZN(n987) );
  INV_X1 U750 ( .A(KEYINPUT33), .ZN(n685) );
  AND2_X1 U751 ( .A1(n987), .A2(n685), .ZN(n686) );
  NAND2_X1 U752 ( .A1(n736), .A2(n686), .ZN(n690) );
  INV_X1 U753 ( .A(n737), .ZN(n687) );
  NAND2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n986) );
  AND2_X1 U755 ( .A1(n687), .A2(n986), .ZN(n688) );
  OR2_X1 U756 ( .A1(KEYINPUT33), .A2(n688), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(KEYINPUT98), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n692), .A2(KEYINPUT33), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n737), .A2(n693), .ZN(n694) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n727) );
  XOR2_X1 U762 ( .A(G1981), .B(G305), .Z(n977) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n759) );
  NAND2_X1 U764 ( .A1(G119), .A2(n903), .ZN(n699) );
  NAND2_X1 U765 ( .A1(G131), .A2(n907), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U767 ( .A1(G107), .A2(n902), .ZN(n701) );
  NAND2_X1 U768 ( .A1(G95), .A2(n906), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  OR2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n884) );
  NAND2_X1 U771 ( .A1(G1991), .A2(n884), .ZN(n713) );
  NAND2_X1 U772 ( .A1(G105), .A2(n906), .ZN(n704) );
  XNOR2_X1 U773 ( .A(n704), .B(KEYINPUT38), .ZN(n711) );
  NAND2_X1 U774 ( .A1(G117), .A2(n902), .ZN(n706) );
  NAND2_X1 U775 ( .A1(G141), .A2(n907), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U777 ( .A1(G129), .A2(n903), .ZN(n707) );
  XNOR2_X1 U778 ( .A(KEYINPUT89), .B(n707), .ZN(n708) );
  NOR2_X1 U779 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n882) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n882), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n935) );
  NAND2_X1 U783 ( .A1(n759), .A2(n935), .ZN(n749) );
  XNOR2_X1 U784 ( .A(G1986), .B(G290), .ZN(n981) );
  NAND2_X1 U785 ( .A1(n759), .A2(n981), .ZN(n714) );
  NAND2_X1 U786 ( .A1(n749), .A2(n714), .ZN(n739) );
  INV_X1 U787 ( .A(n739), .ZN(n715) );
  AND2_X1 U788 ( .A1(n977), .A2(n715), .ZN(n725) );
  NAND2_X1 U789 ( .A1(G104), .A2(n906), .ZN(n717) );
  NAND2_X1 U790 ( .A1(G140), .A2(n907), .ZN(n716) );
  NAND2_X1 U791 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U792 ( .A(KEYINPUT34), .B(n718), .ZN(n723) );
  NAND2_X1 U793 ( .A1(G116), .A2(n902), .ZN(n720) );
  NAND2_X1 U794 ( .A1(G128), .A2(n903), .ZN(n719) );
  NAND2_X1 U795 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U796 ( .A(KEYINPUT35), .B(n721), .Z(n722) );
  NOR2_X1 U797 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U798 ( .A(KEYINPUT36), .B(n724), .ZN(n899) );
  XNOR2_X1 U799 ( .A(KEYINPUT37), .B(G2067), .ZN(n748) );
  NOR2_X1 U800 ( .A1(n899), .A2(n748), .ZN(n942) );
  NAND2_X1 U801 ( .A1(n759), .A2(n942), .ZN(n755) );
  AND2_X1 U802 ( .A1(n725), .A2(n755), .ZN(n726) );
  NAND2_X1 U803 ( .A1(n727), .A2(n726), .ZN(n745) );
  INV_X1 U804 ( .A(n755), .ZN(n743) );
  NAND2_X1 U805 ( .A1(G8), .A2(G166), .ZN(n728) );
  NOR2_X1 U806 ( .A1(G2090), .A2(n728), .ZN(n729) );
  XNOR2_X1 U807 ( .A(n729), .B(KEYINPUT99), .ZN(n734) );
  NOR2_X1 U808 ( .A1(G1981), .A2(G305), .ZN(n730) );
  XOR2_X1 U809 ( .A(n730), .B(KEYINPUT24), .Z(n731) );
  NOR2_X1 U810 ( .A1(n737), .A2(n731), .ZN(n732) );
  XOR2_X1 U811 ( .A(KEYINPUT91), .B(n732), .Z(n738) );
  INV_X1 U812 ( .A(n738), .ZN(n733) );
  AND2_X1 U813 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U814 ( .A1(n736), .A2(n735), .ZN(n741) );
  NOR2_X1 U815 ( .A1(n739), .A2(n514), .ZN(n740) );
  NAND2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n742) );
  OR2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U818 ( .A(n747), .B(n746), .ZN(n762) );
  NAND2_X1 U819 ( .A1(n899), .A2(n748), .ZN(n928) );
  NOR2_X1 U820 ( .A1(G1996), .A2(n882), .ZN(n926) );
  INV_X1 U821 ( .A(n749), .ZN(n752) );
  NOR2_X1 U822 ( .A1(G1991), .A2(n884), .ZN(n937) );
  NOR2_X1 U823 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U824 ( .A1(n937), .A2(n750), .ZN(n751) );
  NOR2_X1 U825 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U826 ( .A1(n926), .A2(n753), .ZN(n754) );
  XNOR2_X1 U827 ( .A(n754), .B(KEYINPUT39), .ZN(n756) );
  NAND2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U829 ( .A(KEYINPUT101), .B(n757), .Z(n758) );
  NAND2_X1 U830 ( .A1(n928), .A2(n758), .ZN(n760) );
  NAND2_X1 U831 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U832 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U833 ( .A(n763), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U834 ( .A(G2451), .B(G2443), .Z(n765) );
  XNOR2_X1 U835 ( .A(KEYINPUT103), .B(G2446), .ZN(n764) );
  XNOR2_X1 U836 ( .A(n765), .B(n764), .ZN(n769) );
  XOR2_X1 U837 ( .A(KEYINPUT104), .B(G2438), .Z(n767) );
  XNOR2_X1 U838 ( .A(G2435), .B(G2454), .ZN(n766) );
  XNOR2_X1 U839 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U840 ( .A(n769), .B(n768), .Z(n771) );
  XNOR2_X1 U841 ( .A(G2427), .B(KEYINPUT102), .ZN(n770) );
  XNOR2_X1 U842 ( .A(n771), .B(n770), .ZN(n774) );
  XOR2_X1 U843 ( .A(G1341), .B(G1348), .Z(n772) );
  XNOR2_X1 U844 ( .A(G2430), .B(n772), .ZN(n773) );
  XOR2_X1 U845 ( .A(n774), .B(n773), .Z(n775) );
  AND2_X1 U846 ( .A1(G14), .A2(n775), .ZN(G401) );
  AND2_X1 U847 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U848 ( .A(n818), .ZN(G299) );
  INV_X1 U849 ( .A(G132), .ZN(G219) );
  INV_X1 U850 ( .A(G82), .ZN(G220) );
  INV_X1 U851 ( .A(G120), .ZN(G236) );
  INV_X1 U852 ( .A(G69), .ZN(G235) );
  INV_X1 U853 ( .A(G108), .ZN(G238) );
  NAND2_X1 U854 ( .A1(G7), .A2(G661), .ZN(n776) );
  XNOR2_X1 U855 ( .A(n776), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U856 ( .A(G223), .ZN(n842) );
  NAND2_X1 U857 ( .A1(n842), .A2(G567), .ZN(n777) );
  XOR2_X1 U858 ( .A(KEYINPUT11), .B(n777), .Z(G234) );
  XOR2_X1 U859 ( .A(G860), .B(KEYINPUT72), .Z(n783) );
  OR2_X1 U860 ( .A1(n783), .A2(n982), .ZN(G153) );
  INV_X1 U861 ( .A(n849), .ZN(n990) );
  NOR2_X1 U862 ( .A1(G868), .A2(n990), .ZN(n779) );
  INV_X1 U863 ( .A(G868), .ZN(n824) );
  NOR2_X1 U864 ( .A1(n824), .A2(G301), .ZN(n778) );
  NOR2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U866 ( .A(KEYINPUT74), .B(n780), .ZN(G284) );
  NAND2_X1 U867 ( .A1(G868), .A2(G286), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G299), .A2(n824), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U870 ( .A1(n783), .A2(G559), .ZN(n784) );
  INV_X1 U871 ( .A(n990), .ZN(n801) );
  NAND2_X1 U872 ( .A1(n784), .A2(n801), .ZN(n785) );
  XNOR2_X1 U873 ( .A(n785), .B(KEYINPUT80), .ZN(n787) );
  XOR2_X1 U874 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n786) );
  XNOR2_X1 U875 ( .A(n787), .B(n786), .ZN(G148) );
  NOR2_X1 U876 ( .A1(G868), .A2(n982), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G868), .A2(n801), .ZN(n788) );
  NOR2_X1 U878 ( .A1(G559), .A2(n788), .ZN(n789) );
  NOR2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U880 ( .A(KEYINPUT81), .B(n791), .Z(G282) );
  NAND2_X1 U881 ( .A1(G123), .A2(n903), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n792), .B(KEYINPUT18), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n902), .A2(G111), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G99), .A2(n906), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G135), .A2(n907), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n936) );
  XNOR2_X1 U889 ( .A(n936), .B(G2096), .ZN(n800) );
  INV_X1 U890 ( .A(G2100), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n800), .A2(n799), .ZN(G156) );
  NAND2_X1 U892 ( .A1(n801), .A2(G559), .ZN(n821) );
  XNOR2_X1 U893 ( .A(n982), .B(n821), .ZN(n802) );
  NOR2_X1 U894 ( .A1(n802), .A2(G860), .ZN(n813) );
  NAND2_X1 U895 ( .A1(n803), .A2(G67), .ZN(n806) );
  NAND2_X1 U896 ( .A1(G55), .A2(n804), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G93), .A2(n807), .ZN(n810) );
  NAND2_X1 U899 ( .A1(G80), .A2(n808), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n823) );
  XNOR2_X1 U902 ( .A(n813), .B(n823), .ZN(G145) );
  XOR2_X1 U903 ( .A(G290), .B(G305), .Z(n814) );
  XNOR2_X1 U904 ( .A(G288), .B(n814), .ZN(n817) );
  XNOR2_X1 U905 ( .A(KEYINPUT19), .B(G303), .ZN(n815) );
  XNOR2_X1 U906 ( .A(n815), .B(n982), .ZN(n816) );
  XOR2_X1 U907 ( .A(n817), .B(n816), .Z(n820) );
  XNOR2_X1 U908 ( .A(n818), .B(n823), .ZN(n819) );
  XNOR2_X1 U909 ( .A(n820), .B(n819), .ZN(n848) );
  XNOR2_X1 U910 ( .A(n821), .B(n848), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n822), .A2(G868), .ZN(n826) );
  NAND2_X1 U912 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U913 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U914 ( .A(KEYINPUT85), .B(n827), .ZN(G295) );
  NAND2_X1 U915 ( .A1(G2078), .A2(G2084), .ZN(n828) );
  XOR2_X1 U916 ( .A(KEYINPUT20), .B(n828), .Z(n829) );
  NAND2_X1 U917 ( .A1(G2090), .A2(n829), .ZN(n830) );
  XNOR2_X1 U918 ( .A(KEYINPUT21), .B(n830), .ZN(n831) );
  NAND2_X1 U919 ( .A1(n831), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U920 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U921 ( .A1(G235), .A2(G236), .ZN(n832) );
  XNOR2_X1 U922 ( .A(n832), .B(KEYINPUT87), .ZN(n833) );
  NOR2_X1 U923 ( .A1(G238), .A2(n833), .ZN(n834) );
  NAND2_X1 U924 ( .A1(G57), .A2(n834), .ZN(n846) );
  NAND2_X1 U925 ( .A1(n846), .A2(G567), .ZN(n840) );
  NOR2_X1 U926 ( .A1(G220), .A2(G219), .ZN(n835) );
  XOR2_X1 U927 ( .A(KEYINPUT22), .B(n835), .Z(n836) );
  NOR2_X1 U928 ( .A1(G218), .A2(n836), .ZN(n837) );
  XNOR2_X1 U929 ( .A(KEYINPUT86), .B(n837), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n838), .A2(G96), .ZN(n847) );
  NAND2_X1 U931 ( .A1(n847), .A2(G2106), .ZN(n839) );
  NAND2_X1 U932 ( .A1(n840), .A2(n839), .ZN(n923) );
  NAND2_X1 U933 ( .A1(G483), .A2(G661), .ZN(n841) );
  NOR2_X1 U934 ( .A1(n923), .A2(n841), .ZN(n845) );
  NAND2_X1 U935 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U938 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  NOR2_X1 U943 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  XOR2_X1 U945 ( .A(KEYINPUT112), .B(n848), .Z(n851) );
  XNOR2_X1 U946 ( .A(G171), .B(n849), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U948 ( .A(n852), .B(G286), .Z(n853) );
  NOR2_X1 U949 ( .A1(G37), .A2(n853), .ZN(G397) );
  XNOR2_X1 U950 ( .A(G1986), .B(G2474), .ZN(n863) );
  XOR2_X1 U951 ( .A(G1956), .B(G1971), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1981), .B(G1976), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(G1961), .B(G1966), .Z(n857) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(G229) );
  XOR2_X1 U961 ( .A(G2678), .B(G2090), .Z(n865) );
  XNOR2_X1 U962 ( .A(G2078), .B(G2084), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U964 ( .A(n866), .B(G2100), .Z(n868) );
  XNOR2_X1 U965 ( .A(G2067), .B(G2072), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U967 ( .A(G2096), .B(KEYINPUT105), .Z(n870) );
  XNOR2_X1 U968 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U970 ( .A(n872), .B(n871), .Z(G227) );
  NAND2_X1 U971 ( .A1(G124), .A2(n903), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G100), .A2(n906), .ZN(n874) );
  XOR2_X1 U974 ( .A(KEYINPUT107), .B(n874), .Z(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G112), .A2(n902), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G136), .A2(n907), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(G162) );
  XOR2_X1 U980 ( .A(G164), .B(n936), .Z(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(KEYINPUT48), .B(n883), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n884), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U985 ( .A(G162), .B(n887), .ZN(n901) );
  XNOR2_X1 U986 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G115), .A2(n902), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G127), .A2(n903), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n898) );
  NAND2_X1 U991 ( .A1(n907), .A2(G139), .ZN(n892) );
  XNOR2_X1 U992 ( .A(KEYINPUT109), .B(n892), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n906), .A2(G103), .ZN(n893) );
  XOR2_X1 U994 ( .A(KEYINPUT108), .B(n893), .Z(n894) );
  NOR2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT110), .B(n896), .Z(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n930) );
  XNOR2_X1 U998 ( .A(n899), .B(n930), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n915) );
  NAND2_X1 U1000 ( .A1(G118), .A2(n902), .ZN(n905) );
  NAND2_X1 U1001 ( .A1(G130), .A2(n903), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(n905), .A2(n904), .ZN(n912) );
  NAND2_X1 U1003 ( .A1(G106), .A2(n906), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(G142), .A2(n907), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(KEYINPUT45), .B(n910), .Z(n911) );
  NOR2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1008 ( .A(G160), .B(n913), .Z(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n923), .ZN(n920) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G397), .A2(n918), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n921), .A2(G395), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n922), .B(KEYINPUT113), .ZN(G225) );
  XOR2_X1 U1018 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1019 ( .A(n923), .ZN(G319) );
  INV_X1 U1020 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n924) );
  XNOR2_X1 U1022 ( .A(KEYINPUT116), .B(n924), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n927), .Z(n929) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n946) );
  XOR2_X1 U1026 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(KEYINPUT50), .B(n933), .ZN(n944) );
  XOR2_X1 U1030 ( .A(G160), .B(G2084), .Z(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n940) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT115), .B(n938), .Z(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1041 ( .A1(n950), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1042 ( .A(G20), .B(n951), .ZN(n955) );
  XNOR2_X1 U1043 ( .A(G1981), .B(G6), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1047 ( .A(KEYINPUT59), .B(G1348), .Z(n956) );
  XNOR2_X1 U1048 ( .A(G4), .B(n956), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(KEYINPUT60), .B(n959), .ZN(n963) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G21), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G5), .B(G1961), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(n963), .A2(n962), .ZN(n972) );
  XOR2_X1 U1055 ( .A(G1986), .B(G24), .Z(n968) );
  XNOR2_X1 U1056 ( .A(G1976), .B(G23), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G22), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(n966), .B(KEYINPUT124), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1061 ( .A(KEYINPUT58), .B(n969), .Z(n970) );
  XNOR2_X1 U1062 ( .A(KEYINPUT125), .B(n970), .ZN(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(KEYINPUT61), .B(n973), .ZN(n975) );
  INV_X1 U1065 ( .A(G16), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n976), .A2(G11), .ZN(n1028) );
  XNOR2_X1 U1068 ( .A(G16), .B(KEYINPUT56), .ZN(n1002) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G168), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1071 ( .A(KEYINPUT57), .B(n979), .Z(n999) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G299), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(G1341), .B(KEYINPUT121), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n983), .B(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n996) );
  AND2_X1 U1077 ( .A1(G303), .A2(G1971), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(G301), .B(G1961), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n990), .B(G1348), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1085 ( .A(KEYINPUT122), .B(n997), .Z(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(KEYINPUT123), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1026) );
  XOR2_X1 U1089 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n1022) );
  XNOR2_X1 U1090 ( .A(G2090), .B(G35), .ZN(n1017) );
  XNOR2_X1 U1091 ( .A(G1991), .B(G25), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G2067), .B(G26), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G2072), .B(G33), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT117), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(G28), .A2(n1008), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1996), .B(G32), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1009), .B(G27), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(KEYINPUT118), .B(n1012), .Z(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(G2084), .B(G34), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT54), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1022), .B(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(G29), .A2(n1023), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(KEYINPUT120), .B(n1024), .Z(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1114 ( .A(n1031), .B(KEYINPUT126), .ZN(n1032) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

