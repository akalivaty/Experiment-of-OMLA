//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  INV_X1    g0007(.A(G264), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G68), .C2(G238), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G50), .A2(G226), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G77), .A2(G244), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n203), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n206), .B(new_n224), .C1(new_n231), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(KEYINPUT67), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n208), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n230), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n252), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n255), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT25), .B1(new_n255), .B2(new_n207), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n260), .A2(new_n207), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G1), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT5), .B(G41), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n211), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n213), .A2(G1698), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n271), .A2(new_n273), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G294), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g0079(.A1(G264), .A2(new_n269), .B1(new_n279), .B2(new_n265), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n268), .A2(G274), .A3(new_n267), .ZN(new_n281));
  AOI21_X1  g0081(.A(G200), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI211_X1 g0082(.A(new_n208), .B(new_n265), .C1(new_n267), .C2(new_n268), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  OAI211_X1 g0084(.A(G1), .B(G13), .C1(new_n270), .C2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n277), .B2(new_n278), .ZN(new_n286));
  INV_X1    g0086(.A(new_n281), .ZN(new_n287));
  NOR4_X1   g0087(.A1(new_n283), .A2(new_n286), .A3(G190), .A4(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n229), .A2(new_n290), .A3(G87), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT23), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n295), .A2(G20), .B1(new_n296), .B2(new_n207), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n226), .A2(new_n228), .A3(new_n296), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(new_n207), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n229), .A2(new_n290), .A3(new_n292), .A4(G87), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n294), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XOR2_X1   g0101(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n294), .A2(new_n299), .A3(new_n302), .A4(new_n300), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n257), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT88), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT88), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n304), .A2(new_n308), .A3(new_n257), .A4(new_n305), .ZN(new_n309));
  AOI211_X1 g0109(.A(new_n264), .B(new_n289), .C1(new_n307), .C2(new_n309), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n283), .A2(new_n286), .A3(new_n287), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G169), .B2(new_n311), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n307), .A2(new_n309), .ZN(new_n315));
  INV_X1    g0115(.A(new_n264), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT89), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n289), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT89), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n264), .B1(new_n307), .B2(new_n309), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n320), .B(new_n321), .C1(new_n322), .C2(new_n314), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT18), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n271), .A2(new_n275), .A3(G226), .A4(G1698), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT76), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n290), .A2(KEYINPUT76), .A3(G226), .A4(G1698), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G87), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n290), .A2(G223), .A3(new_n272), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n265), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT69), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT68), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G45), .ZN(new_n337));
  AOI21_X1  g0137(.A(G41), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n334), .B1(new_n338), .B2(G1), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT68), .B(G45), .ZN(new_n340));
  OAI211_X1 g0140(.A(KEYINPUT69), .B(new_n252), .C1(new_n340), .C2(G41), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n339), .A2(G274), .A3(new_n285), .A4(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(G1), .B1(new_n284), .B2(new_n266), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n265), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G232), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n333), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G169), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n333), .A2(G179), .A3(new_n342), .A4(new_n345), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n274), .A2(G33), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT73), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT73), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n271), .A2(new_n275), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT7), .B1(new_n354), .B2(new_n229), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT7), .B(new_n225), .C1(new_n349), .C2(new_n350), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT74), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n271), .A2(new_n275), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT7), .A4(new_n225), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G68), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n220), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(G58), .A2(G68), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G20), .A2(G33), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n366), .A2(G20), .B1(G159), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n362), .A2(KEYINPUT16), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT64), .B(G20), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT7), .B1(new_n370), .B2(new_n290), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n358), .A2(new_n372), .A3(new_n225), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n368), .B1(new_n374), .B2(new_n363), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n369), .A2(new_n257), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n257), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n253), .ZN(new_n380));
  XOR2_X1   g0180(.A(KEYINPUT8), .B(G58), .Z(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n381), .ZN(new_n383));
  INV_X1    g0183(.A(new_n255), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n386), .B(KEYINPUT75), .ZN(new_n387));
  AOI221_X4 g0187(.A(new_n325), .B1(new_n347), .B2(new_n348), .C1(new_n378), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n378), .A2(new_n387), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n347), .A2(new_n348), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT18), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n387), .ZN(new_n394));
  INV_X1    g0194(.A(new_n368), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n370), .B1(new_n351), .B2(new_n353), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n357), .B(new_n360), .C1(new_n396), .C2(KEYINPUT7), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n397), .B2(G68), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n379), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n394), .B1(new_n399), .B2(new_n377), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n346), .A2(G200), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n333), .A2(G190), .A3(new_n342), .A4(new_n345), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n400), .A2(KEYINPUT17), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n378), .A2(new_n401), .A3(new_n402), .A4(new_n387), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n393), .A2(new_n408), .A3(KEYINPUT77), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n344), .A2(G244), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G238), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n290), .B(new_n411), .C1(new_n221), .C2(G1698), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n412), .B(new_n265), .C1(G107), .C2(new_n290), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n342), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n414), .A2(G200), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n384), .A2(G77), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n381), .A2(new_n367), .B1(new_n370), .B2(G77), .ZN(new_n417));
  XOR2_X1   g0217(.A(KEYINPUT15), .B(G87), .Z(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n229), .A2(G33), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n416), .B1(new_n421), .B2(new_n257), .ZN(new_n422));
  INV_X1    g0222(.A(G77), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n380), .ZN(new_n424));
  INV_X1    g0224(.A(G190), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n414), .A2(new_n425), .ZN(new_n426));
  OR3_X1    g0226(.A1(new_n415), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G50), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n225), .B1(new_n365), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(G150), .B2(new_n367), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n420), .B2(new_n383), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(new_n257), .B1(new_n428), .B2(new_n255), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n428), .B2(new_n380), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT9), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n344), .A2(G226), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n272), .A2(G222), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G223), .A2(G1698), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n290), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(new_n265), .C1(G77), .C2(new_n290), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n342), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G200), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(G190), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n434), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT10), .ZN(new_n447));
  INV_X1    g0247(.A(G169), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n414), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n424), .B(new_n449), .C1(G179), .C2(new_n414), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n409), .A2(new_n427), .A3(new_n447), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n440), .A2(new_n448), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n433), .C1(G179), .C2(new_n440), .ZN(new_n453));
  XOR2_X1   g0253(.A(new_n453), .B(KEYINPUT70), .Z(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G303), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n285), .B1(new_n358), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G264), .A2(G1698), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n290), .B(new_n459), .C1(new_n213), .C2(G1698), .ZN(new_n460));
  AOI22_X1  g0260(.A1(G270), .A2(new_n269), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n281), .ZN(new_n462));
  INV_X1    g0262(.A(G116), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n255), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n229), .B(new_n465), .C1(G33), .C2(new_n212), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n256), .A2(new_n230), .B1(G20), .B2(new_n463), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n466), .A2(KEYINPUT20), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT20), .B1(new_n466), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT85), .B1(new_n260), .B2(new_n463), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n258), .A2(new_n472), .A3(G116), .A4(new_n259), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G169), .B(new_n462), .C1(new_n470), .C2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT21), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n466), .A2(new_n467), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT20), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n466), .A2(KEYINPUT20), .A3(new_n467), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(new_n464), .A3(new_n471), .A4(new_n473), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(KEYINPUT21), .A3(G169), .A4(new_n462), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(G179), .A3(new_n281), .A4(new_n461), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n477), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n483), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n462), .A2(G200), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n489), .C1(new_n425), .C2(new_n462), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n290), .A2(G244), .A3(new_n272), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(KEYINPUT80), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n465), .B1(new_n493), .B2(KEYINPUT80), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n211), .A2(new_n272), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n290), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(KEYINPUT80), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n290), .A2(G244), .A3(new_n272), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n287), .B1(new_n500), .B2(new_n265), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n269), .A2(KEYINPUT81), .A3(G257), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT81), .B1(new_n269), .B2(G257), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(G190), .A3(new_n504), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n384), .A2(G97), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n260), .B2(new_n212), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n212), .A2(new_n207), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n370), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n367), .A2(G77), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT78), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n516), .B(new_n518), .C1(new_n374), .C2(new_n207), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n510), .B1(new_n519), .B2(new_n257), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT79), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI211_X1 g0322(.A(KEYINPUT79), .B(new_n510), .C1(new_n519), .C2(new_n257), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n506), .B(new_n507), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n520), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n501), .A2(G179), .A3(new_n504), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n448), .B1(new_n501), .B2(new_n504), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n272), .A2(G244), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n290), .B(new_n530), .C1(G238), .C2(G1698), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n285), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n267), .A2(G250), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n266), .A2(G1), .A3(G274), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n534), .A2(new_n265), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(G169), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n312), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n358), .A2(new_n370), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n229), .A2(G33), .A3(G97), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  AOI22_X1  g0342(.A1(G68), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT82), .B1(new_n370), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT82), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n229), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n210), .A2(new_n212), .A3(new_n207), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n379), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT83), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n260), .A2(new_n419), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n384), .A2(new_n418), .ZN(new_n554));
  NOR4_X1   g0354(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n540), .A2(G68), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n541), .A2(new_n542), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n550), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n554), .B1(new_n558), .B2(new_n257), .ZN(new_n559));
  INV_X1    g0359(.A(new_n553), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT83), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n539), .B1(new_n555), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n258), .A2(G87), .A3(new_n259), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n537), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT84), .B1(new_n565), .B2(new_n425), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT84), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n537), .A2(new_n568), .A3(G190), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n564), .A2(new_n566), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n524), .A2(new_n529), .A3(new_n562), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n491), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n221), .A2(G1698), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(G226), .B2(G1698), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n574), .A2(new_n358), .B1(new_n270), .B2(new_n212), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n265), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n344), .A2(G238), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n342), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g0378(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n579), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n342), .A2(new_n581), .A3(new_n577), .A4(new_n576), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n578), .A2(KEYINPUT13), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n585), .A2(G190), .A3(new_n582), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n384), .A2(KEYINPUT12), .A3(G68), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT12), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n255), .B2(new_n363), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n587), .A2(new_n589), .B1(new_n363), .B2(new_n380), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n367), .A2(G50), .ZN(new_n591));
  OAI221_X1 g0391(.A(new_n591), .B1(new_n225), .B2(G68), .C1(new_n420), .C2(new_n423), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n257), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n593), .A2(KEYINPUT11), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(KEYINPUT11), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n590), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n584), .A2(new_n586), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT72), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n584), .A2(new_n596), .A3(KEYINPUT72), .A4(new_n586), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n583), .A2(G169), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT14), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n585), .A2(G179), .A3(new_n582), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT14), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n583), .A2(new_n605), .A3(G169), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n596), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT77), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n406), .B(new_n403), .C1(new_n388), .C2(new_n391), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n324), .A2(new_n456), .A3(new_n572), .A4(new_n613), .ZN(G372));
  INV_X1    g0414(.A(new_n601), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n609), .B1(new_n615), .B2(new_n450), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT90), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(KEYINPUT90), .B(new_n609), .C1(new_n615), .C2(new_n450), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n408), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n393), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n455), .B1(new_n621), .B2(new_n447), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n456), .A2(new_n613), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n505), .A2(G169), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n520), .B1(new_n624), .B2(new_n526), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n562), .A3(new_n570), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n320), .B1(new_n317), .B2(new_n486), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n627), .B(new_n562), .C1(new_n628), .C2(new_n571), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n522), .A2(new_n523), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n528), .B2(new_n527), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n562), .A2(new_n570), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n631), .A2(new_n632), .A3(KEYINPUT26), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n622), .B1(new_n623), .B2(new_n634), .ZN(G369));
  NOR2_X1   g0435(.A1(new_n370), .A2(new_n254), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n252), .ZN(new_n637));
  OR3_X1    g0437(.A1(new_n637), .A2(KEYINPUT91), .A3(KEYINPUT27), .ZN(new_n638));
  INV_X1    g0438(.A(G213), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n637), .B2(KEYINPUT27), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT91), .B1(new_n637), .B2(KEYINPUT27), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n318), .B2(new_n323), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n317), .B2(new_n644), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n324), .A2(new_n322), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n644), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n488), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n486), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n491), .B2(new_n651), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n324), .A2(new_n486), .A3(new_n650), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n317), .A2(new_n650), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0461(.A(new_n204), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n549), .A2(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n233), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n664), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n650), .B1(new_n629), .B2(new_n633), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT94), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT26), .B1(new_n631), .B2(new_n632), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n625), .A2(new_n562), .A3(new_n570), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n562), .B1(new_n628), .B2(new_n571), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n650), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  INV_X1    g0480(.A(new_n670), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n671), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n505), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n537), .A2(new_n461), .A3(G179), .A4(new_n281), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT93), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n684), .A2(new_n686), .A3(new_n280), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n501), .A2(new_n280), .A3(new_n504), .ZN(new_n690));
  OAI211_X1 g0490(.A(KEYINPUT93), .B(new_n687), .C1(new_n690), .C2(new_n685), .ZN(new_n691));
  INV_X1    g0491(.A(new_n311), .ZN(new_n692));
  AOI21_X1  g0492(.A(G179), .B1(new_n461), .B2(new_n281), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n505), .A2(new_n692), .A3(new_n565), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n689), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(new_n644), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(KEYINPUT31), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n645), .B2(new_n572), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n683), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n669), .B1(new_n703), .B2(G1), .ZN(G364));
  NAND2_X1  g0504(.A1(new_n636), .A2(G45), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n664), .A2(new_n705), .A3(G1), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n653), .A2(G330), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n654), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n290), .A2(G355), .A3(new_n204), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n250), .A2(new_n266), .B1(new_n667), .B2(new_n340), .ZN(new_n711));
  INV_X1    g0511(.A(new_n354), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n662), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI221_X1 g0514(.A(new_n710), .B1(G116), .B2(new_n204), .C1(new_n711), .C2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G13), .A2(G33), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n230), .B1(G20), .B2(new_n448), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n718), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n229), .A2(new_n312), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G190), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G200), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n290), .B1(new_n726), .B2(new_n220), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n229), .A2(G190), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(G179), .A3(new_n442), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n442), .A2(G179), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT98), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G20), .A3(G190), .ZN(new_n736));
  OAI22_X1  g0536(.A1(new_n733), .A2(new_n423), .B1(new_n210), .B2(new_n736), .ZN(new_n737));
  OR3_X1    g0537(.A1(new_n229), .A2(KEYINPUT97), .A3(G190), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT97), .B1(new_n229), .B2(G190), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n735), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n727), .B(new_n737), .C1(G107), .C2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n728), .A2(G179), .A3(G200), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G68), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n738), .A2(new_n746), .A3(new_n739), .ZN(new_n747));
  INV_X1    g0547(.A(G159), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT32), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT96), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n724), .B2(new_n442), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n723), .A2(KEYINPUT96), .A3(G190), .A4(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n370), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n754), .A2(G50), .B1(G97), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n742), .A2(new_n745), .A3(new_n750), .A4(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G294), .ZN(new_n759));
  INV_X1    g0559(.A(new_n756), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n358), .B1(new_n759), .B2(new_n760), .C1(new_n736), .C2(new_n457), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n725), .A2(G322), .ZN(new_n762));
  INV_X1    g0562(.A(G329), .ZN(new_n763));
  XNOR2_X1  g0563(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(G317), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n762), .B1(new_n763), .B2(new_n747), .C1(new_n743), .C2(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n761), .B(new_n766), .C1(G283), .C2(new_n741), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  INV_X1    g0569(.A(new_n754), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n767), .B1(new_n768), .B2(new_n729), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n758), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n719), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n721), .B1(new_n653), .B2(new_n722), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n709), .B1(new_n774), .B2(new_n707), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT100), .Z(G396));
  NAND2_X1  g0576(.A1(new_n644), .A2(new_n424), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n427), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n450), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n450), .A2(new_n644), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n681), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n650), .B(new_n782), .C1(new_n629), .C2(new_n633), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OR3_X1    g0585(.A1(new_n701), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n701), .B1(new_n783), .B2(new_n785), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n786), .A2(new_n787), .A3(new_n706), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n754), .A2(G137), .B1(G143), .B2(new_n725), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n744), .A2(G150), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n789), .B(new_n790), .C1(new_n748), .C2(new_n733), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT34), .Z(new_n792));
  INV_X1    g0592(.A(new_n747), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(G132), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n741), .A2(G68), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n756), .A2(G58), .ZN(new_n796));
  INV_X1    g0596(.A(new_n736), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n354), .B1(new_n797), .B2(G50), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n744), .A2(KEYINPUT101), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n744), .A2(KEYINPUT101), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n358), .B1(new_n733), .B2(new_n463), .C1(new_n800), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n747), .A2(new_n768), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n726), .A2(new_n759), .B1(new_n212), .B2(new_n760), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(new_n754), .C2(G303), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n741), .A2(G87), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(new_n207), .C2(new_n736), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n799), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n719), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n719), .A2(new_n716), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n423), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n781), .A2(new_n716), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n811), .A2(new_n707), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n788), .A2(new_n815), .ZN(G384));
  NOR2_X1   g0616(.A1(new_n683), .A2(new_n623), .ZN(new_n817));
  INV_X1    g0617(.A(new_n622), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT39), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n400), .A2(new_n642), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT37), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n389), .A2(new_n390), .ZN(new_n825));
  INV_X1    g0625(.A(new_n642), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n389), .A2(new_n826), .ZN(new_n827));
  AND4_X1   g0627(.A1(new_n824), .A2(new_n825), .A3(new_n827), .A4(new_n404), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT104), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n612), .A2(new_n823), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n390), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n404), .B1(new_n400), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT37), .B1(new_n832), .B2(new_n823), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n825), .A2(new_n827), .A3(new_n824), .A4(new_n404), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(KEYINPUT104), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n822), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n362), .A2(new_n368), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n376), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n399), .A2(new_n838), .B1(new_n382), .B2(new_n385), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n642), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n612), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n369), .A2(new_n257), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n398), .A2(KEYINPUT16), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n386), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n347), .A2(new_n348), .A3(new_n642), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n824), .B1(new_n846), .B2(new_n404), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT102), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n845), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n404), .B1(new_n839), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT37), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(new_n834), .A3(KEYINPUT102), .ZN(new_n853));
  AND4_X1   g0653(.A1(KEYINPUT38), .A2(new_n841), .A3(new_n849), .A4(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n820), .B1(new_n836), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n609), .A2(new_n644), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n841), .A2(new_n849), .A3(new_n853), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n612), .A2(new_n840), .B1(new_n848), .B2(new_n847), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(KEYINPUT38), .A3(new_n853), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(KEYINPUT39), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n855), .A2(new_n856), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n859), .A2(new_n861), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n608), .A2(new_n644), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n601), .A2(new_n609), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n601), .B2(new_n609), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n784), .B2(new_n780), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n864), .A2(new_n869), .B1(new_n392), .B2(new_n642), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n819), .B(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n860), .B2(new_n853), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n854), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n645), .A2(new_n572), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT105), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n699), .B(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n697), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n865), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n610), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n601), .A2(new_n609), .A3(new_n865), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n781), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n873), .B1(new_n875), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n823), .B1(new_n392), .B2(new_n407), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n828), .A2(new_n829), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n835), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n821), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n873), .B1(new_n890), .B2(new_n861), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n782), .B1(new_n866), .B2(new_n867), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n698), .B2(new_n878), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n886), .A2(new_n894), .A3(G330), .ZN(new_n895));
  INV_X1    g0695(.A(G330), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n698), .B2(new_n878), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n456), .A2(new_n897), .A3(new_n613), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n864), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n900), .A2(new_n873), .B1(new_n891), .B2(new_n893), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n880), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n899), .B1(new_n902), .B2(new_n623), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n872), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n252), .B2(new_n636), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n463), .B1(new_n515), .B2(KEYINPUT35), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n906), .B(new_n231), .C1(KEYINPUT35), .C2(new_n515), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT36), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n667), .A2(new_n423), .A3(new_n364), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n363), .A2(G50), .ZN(new_n910));
  OAI211_X1 g0710(.A(G1), .B(new_n254), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n905), .A2(new_n908), .A3(new_n911), .ZN(G367));
  OAI221_X1 g0712(.A(new_n720), .B1(new_n204), .B2(new_n419), .C1(new_n243), .C2(new_n714), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT108), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n725), .A2(G150), .B1(G68), .B2(new_n756), .ZN(new_n915));
  INV_X1    g0715(.A(G137), .ZN(new_n916));
  OAI221_X1 g0716(.A(new_n915), .B1(new_n916), .B2(new_n747), .C1(new_n803), .C2(new_n748), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(G143), .B2(new_n754), .ZN(new_n918));
  INV_X1    g0718(.A(new_n733), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G50), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n358), .B1(new_n797), .B2(G58), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n741), .A2(G77), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n918), .A2(new_n920), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT46), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n736), .B2(new_n463), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n797), .A2(KEYINPUT46), .A3(G116), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n925), .B(new_n926), .C1(new_n803), .C2(new_n759), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT109), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n741), .A2(G97), .ZN(new_n929));
  INV_X1    g0729(.A(G317), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n930), .B2(new_n747), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n354), .B1(new_n770), .B2(new_n768), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n931), .B(new_n932), .C1(G107), .C2(new_n756), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n928), .B(new_n933), .C1(new_n457), .C2(new_n726), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n733), .A2(new_n800), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n923), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT47), .Z(new_n937));
  OAI211_X1 g0737(.A(new_n707), .B(new_n914), .C1(new_n937), .C2(new_n773), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT110), .Z(new_n939));
  OR2_X1    g0739(.A1(new_n650), .A2(new_n564), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(new_n562), .A3(new_n570), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n562), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n939), .B1(new_n722), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n705), .A2(G1), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n630), .A2(new_n644), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n529), .A3(new_n524), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n631), .B2(new_n650), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n659), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT45), .Z(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT44), .B1(new_n659), .B2(new_n947), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n659), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n656), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n649), .B1(new_n487), .B2(new_n644), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n954), .A2(new_n654), .A3(new_n657), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n654), .B1(new_n954), .B2(new_n657), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n702), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n703), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n663), .B(KEYINPUT41), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n944), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n947), .B(KEYINPUT106), .Z(new_n963));
  NOR3_X1   g0763(.A1(new_n963), .A2(new_n322), .A3(new_n314), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n650), .B1(new_n964), .B2(new_n625), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n657), .A2(new_n946), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT42), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT107), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n966), .A2(KEYINPUT42), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n965), .A2(KEYINPUT107), .A3(new_n967), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n975), .B1(new_n973), .B2(new_n976), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n978), .A2(new_n979), .B1(new_n656), .B2(new_n963), .ZN(new_n980));
  INV_X1    g0780(.A(new_n979), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n656), .A2(new_n963), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n982), .A3(new_n977), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n943), .B1(new_n962), .B2(new_n984), .ZN(G387));
  OR3_X1    g0785(.A1(new_n383), .A2(KEYINPUT50), .A3(G50), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT50), .B1(new_n383), .B2(G50), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n986), .A2(new_n987), .A3(new_n266), .A4(new_n665), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G68), .B2(G77), .ZN(new_n989));
  INV_X1    g0789(.A(new_n340), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n713), .B1(new_n239), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n290), .B(new_n204), .C1(G116), .C2(new_n549), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n204), .A2(G107), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n720), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n756), .A2(new_n418), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n730), .A2(G68), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n797), .A2(G77), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n929), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n754), .A2(G159), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT111), .Z(new_n1001));
  AOI21_X1  g0801(.A(new_n354), .B1(new_n793), .B2(G150), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n428), .C2(new_n726), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n999), .B(new_n1003), .C1(new_n381), .C2(new_n744), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n754), .A2(G322), .B1(G317), .B2(new_n725), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n733), .B2(new_n457), .C1(new_n768), .C2(new_n803), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT48), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n800), .B2(new_n760), .C1(new_n759), .C2(new_n736), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT49), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n354), .B1(new_n747), .B2(new_n769), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G116), .B2(new_n741), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1004), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n707), .B(new_n995), .C1(new_n1012), .C2(new_n773), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n649), .B2(new_n718), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n957), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n1015), .B2(new_n944), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n663), .B1(new_n1015), .B2(new_n703), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n1017), .B2(new_n958), .ZN(G393));
  INV_X1    g0818(.A(new_n953), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n958), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1021), .A2(new_n959), .A3(new_n663), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n953), .A2(new_n944), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n793), .A2(G143), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n808), .B(new_n1024), .C1(new_n363), .C2(new_n736), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n754), .A2(G150), .B1(G159), .B2(new_n725), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT51), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(new_n381), .C2(new_n919), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n756), .A2(G77), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n803), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(G50), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n712), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT112), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n290), .B1(new_n793), .B2(G322), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n207), .B2(new_n740), .C1(new_n803), .C2(new_n457), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n754), .A2(G317), .B1(G311), .B2(new_n725), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1035), .B(new_n1037), .C1(G116), .C2(new_n756), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n800), .B2(new_n736), .C1(new_n759), .C2(new_n729), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n773), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n720), .B1(new_n212), .B2(new_n204), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n713), .B2(new_n247), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1040), .A2(new_n706), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n963), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1043), .B1(new_n722), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1022), .A2(new_n1023), .A3(new_n1045), .ZN(G390));
  AND3_X1   g0846(.A1(new_n859), .A2(KEYINPUT39), .A3(new_n861), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT39), .B1(new_n890), .B2(new_n861), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n716), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT54), .B(G143), .Z(new_n1050));
  AOI22_X1  g0850(.A1(new_n919), .A2(new_n1050), .B1(G159), .B2(new_n756), .ZN(new_n1051));
  INV_X1    g0851(.A(G125), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1051), .B1(new_n428), .B2(new_n740), .C1(new_n1052), .C2(new_n747), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G137), .B2(new_n1030), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n754), .A2(G128), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n797), .A2(G150), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT53), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1057), .A2(new_n358), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G132), .B2(new_n725), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n919), .A2(G97), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n725), .A2(G116), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1061), .A2(new_n795), .A3(new_n1029), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n754), .A2(G283), .B1(G87), .B2(new_n797), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n759), .B2(new_n747), .C1(new_n207), .C2(new_n803), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1063), .A2(new_n1065), .A3(new_n290), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT114), .Z(new_n1067));
  OAI21_X1  g0867(.A(new_n719), .B1(new_n1060), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n812), .A2(new_n383), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1049), .A2(new_n707), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n784), .A2(new_n780), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n868), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n856), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n855), .A2(new_n862), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n836), .B2(new_n854), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n650), .B(new_n779), .C1(new_n676), .C2(new_n677), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n868), .B1(new_n1077), .B2(new_n780), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n700), .A2(G330), .A3(new_n1072), .A4(new_n782), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1075), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n880), .A2(new_n884), .A3(G330), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT113), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n897), .A2(KEYINPUT113), .A3(new_n884), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1047), .A2(new_n1048), .B1(new_n856), .B2(new_n869), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1077), .A2(new_n780), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1074), .B1(new_n854), .B2(new_n836), .C1(new_n1088), .C2(new_n868), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1081), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n944), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1070), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n868), .B1(new_n701), .B2(new_n781), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1071), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1080), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1072), .B1(new_n897), .B2(new_n782), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1088), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n622), .B(new_n898), .C1(new_n683), .C2(new_n623), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1087), .A2(new_n1089), .A3(new_n1097), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n1086), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n664), .B1(new_n1104), .B2(new_n1091), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1093), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(G378));
  INV_X1    g0912(.A(KEYINPUT57), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n447), .A2(new_n453), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n826), .A2(new_n433), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n447), .A2(new_n453), .A3(new_n1117), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n895), .A2(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1119), .A2(KEYINPUT116), .A3(new_n1121), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT116), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n886), .A2(new_n894), .A3(new_n1127), .A4(G330), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1124), .A2(new_n871), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n871), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1102), .B1(new_n1108), .B2(new_n1101), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1113), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n871), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1123), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n901), .B2(G330), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1128), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1124), .A2(new_n871), .A3(new_n1128), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1095), .A2(new_n1071), .B1(new_n1099), .B2(new_n1088), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1103), .B1(new_n1091), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(KEYINPUT117), .B(new_n1134), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n1143), .A3(KEYINPUT57), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1133), .A2(new_n1145), .A3(new_n663), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n944), .ZN(new_n1148));
  INV_X1    g0948(.A(G132), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n743), .A2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n797), .A2(new_n1050), .B1(new_n725), .B2(G128), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT115), .Z(new_n1152));
  AOI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(G150), .C2(new_n756), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n1052), .B2(new_n770), .C1(new_n916), .C2(new_n729), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT59), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n748), .B2(new_n740), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n712), .A2(G41), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n428), .B1(G33), .B2(G41), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1155), .A2(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n725), .A2(G107), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n756), .A2(G68), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n998), .A2(new_n1161), .A3(new_n1162), .A4(new_n1158), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n741), .A2(G58), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n800), .B2(new_n747), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G116), .C2(new_n754), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n212), .B2(new_n743), .C1(new_n419), .C2(new_n729), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT58), .Z(new_n1168));
  OAI21_X1  g0968(.A(new_n719), .B1(new_n1160), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n812), .A2(new_n428), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1127), .A2(new_n716), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1169), .A2(new_n707), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1148), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1146), .A2(new_n1174), .ZN(G375));
  AOI22_X1  g0975(.A1(new_n1030), .A2(new_n1050), .B1(G137), .B2(new_n725), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1149), .B2(new_n770), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT120), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n354), .B1(new_n793), .B2(G128), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1179), .B(new_n1164), .C1(new_n428), .C2(new_n760), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G150), .B2(new_n730), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1178), .B(new_n1181), .C1(new_n748), .C2(new_n736), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n793), .A2(G303), .B1(new_n797), .B2(G97), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT119), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n358), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G283), .B2(new_n725), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1030), .A2(G116), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1187));
  AND4_X1   g0987(.A1(new_n922), .A2(new_n1186), .A3(new_n996), .A4(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n207), .B2(new_n733), .C1(new_n759), .C2(new_n770), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n773), .B1(new_n1182), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n706), .B(new_n1190), .C1(new_n363), .C2(new_n812), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n868), .A2(new_n716), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT118), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1101), .A2(new_n944), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1096), .A2(new_n1102), .A3(new_n1100), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n961), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n1105), .B2(new_n1196), .ZN(G381));
  OR2_X1    g0997(.A1(G393), .A2(G396), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(G387), .A2(new_n1198), .A3(G384), .A4(G381), .ZN(new_n1199));
  INV_X1    g0999(.A(G390), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n664), .B1(new_n1201), .B2(new_n1113), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1173), .B1(new_n1202), .B2(new_n1145), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1111), .A4(new_n1203), .ZN(G407));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1111), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G407), .B(G213), .C1(G343), .C2(new_n1205), .ZN(G409));
  NOR2_X1   g1006(.A1(new_n639), .A2(G343), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(G2897), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT60), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1195), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1142), .A2(KEYINPUT60), .A3(new_n1102), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n1104), .A4(new_n663), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1213), .A2(G384), .A3(new_n1194), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G384), .B1(new_n1213), .B2(new_n1194), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1209), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(new_n1194), .ZN(new_n1217));
  INV_X1    g1017(.A(G384), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1213), .A2(G384), .A3(new_n1194), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1220), .A3(new_n1208), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1216), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1207), .B1(G375), .B2(G378), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1143), .A2(new_n1147), .A3(new_n961), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT121), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1141), .A2(new_n944), .A3(new_n1144), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(new_n1172), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1228), .A3(new_n1111), .A4(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1222), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT122), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G387), .A2(new_n1200), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G390), .B(new_n943), .C1(new_n962), .C2(new_n984), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(G393), .B(G396), .Z(new_n1236));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G387), .B2(new_n1200), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1235), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1236), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1233), .A2(new_n1234), .A3(new_n1237), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G375), .A2(G378), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1207), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1230), .A4(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT63), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1232), .A2(new_n1242), .A3(new_n1243), .A4(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT124), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1231), .B2(KEYINPUT61), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1216), .A2(new_n1221), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1203), .B2(new_n1111), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1230), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(KEYINPUT124), .A3(new_n1243), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1251), .A2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1223), .A2(KEYINPUT62), .A3(new_n1230), .A4(new_n1246), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT126), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1247), .A2(KEYINPUT125), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT125), .B1(new_n1247), .B2(new_n1260), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1257), .B1(new_n1259), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1249), .B1(new_n1264), .B2(new_n1242), .ZN(G405));
  NAND2_X1  g1065(.A1(new_n1233), .A2(KEYINPUT123), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1266), .A2(new_n1240), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1241), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT127), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1244), .A2(new_n1205), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(new_n1246), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT127), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1239), .A2(new_n1273), .A3(new_n1241), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1269), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1242), .A2(new_n1271), .A3(KEYINPUT127), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(G402));
endmodule


