//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT72), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT31), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G137), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT66), .B1(new_n193), .B2(G137), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  OAI211_X1 g013(.A(KEYINPUT66), .B(KEYINPUT11), .C1(new_n193), .C2(G137), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G134), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n195), .B1(new_n194), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n192), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n196), .ZN(new_n206));
  INV_X1    g020(.A(new_n200), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT11), .B1(new_n203), .B2(KEYINPUT66), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n204), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(KEYINPUT69), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n214));
  OAI21_X1  g028(.A(G128), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(new_n216), .A3(G143), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n221), .A2(new_n218), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n205), .A2(new_n211), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n194), .B1(new_n207), .B2(new_n208), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(new_n195), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI221_X1 g048(.A(new_n194), .B1(new_n232), .B2(new_n195), .C1(new_n207), .C2(new_n208), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  OR2_X1    g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n216), .A2(G143), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n237), .B(new_n238), .C1(new_n213), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n237), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n221), .A2(new_n243), .A3(new_n218), .A4(new_n223), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n219), .A2(KEYINPUT64), .A3(new_n237), .A4(new_n238), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n236), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n205), .A2(new_n211), .A3(KEYINPUT70), .A4(new_n227), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n230), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT30), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n227), .A2(new_n209), .A3(new_n210), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n247), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g069(.A1(KEYINPUT68), .A2(G116), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT68), .A2(G116), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(G119), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G116), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G119), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT2), .B(G113), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n261), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n263), .B(new_n258), .C1(new_n259), .C2(G119), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n255), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(G237), .A2(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n268), .B(KEYINPUT27), .Z(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n265), .B1(new_n236), .B2(new_n246), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n230), .A2(new_n272), .A3(new_n248), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n230), .A2(new_n272), .A3(KEYINPUT71), .A4(new_n248), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI211_X1 g091(.A(new_n190), .B(new_n191), .C1(new_n266), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n276), .ZN(new_n279));
  INV_X1    g093(.A(new_n271), .ZN(new_n280));
  INV_X1    g094(.A(new_n265), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n253), .B1(new_n249), .B2(KEYINPUT30), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n279), .B(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT72), .B1(new_n283), .B2(KEYINPUT31), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n279), .A2(new_n280), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(new_n250), .B2(new_n254), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n272), .A2(new_n228), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n289), .A2(KEYINPUT28), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n247), .A2(new_n252), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(new_n281), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n275), .B2(new_n276), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT73), .B(KEYINPUT28), .Z(new_n294));
  OAI21_X1  g108(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n191), .A2(new_n288), .B1(new_n295), .B2(new_n271), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n189), .B1(new_n285), .B2(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT74), .B(KEYINPUT32), .Z(new_n298));
  OAI21_X1  g112(.A(new_n187), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT31), .B1(new_n286), .B2(new_n287), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n190), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n288), .A2(new_n191), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n295), .A2(new_n271), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n283), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n301), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n188), .ZN(new_n306));
  INV_X1    g120(.A(new_n298), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(KEYINPUT75), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n249), .A2(new_n265), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n249), .A2(KEYINPUT76), .A3(new_n265), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n279), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT28), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n280), .A2(KEYINPUT29), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n290), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n315), .A2(KEYINPUT77), .A3(new_n290), .A4(new_n316), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n279), .B1(new_n282), .B2(new_n281), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT29), .B1(new_n321), .B2(new_n271), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n280), .B(new_n290), .C1(new_n293), .C2(new_n294), .ZN(new_n323));
  AOI21_X1  g137(.A(G902), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n319), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(KEYINPUT32), .A2(new_n297), .B1(new_n325), .B2(G472), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n309), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G119), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G128), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT78), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n328), .A3(G128), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n330), .B(new_n332), .C1(new_n328), .C2(G128), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT24), .B(G110), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n328), .A2(G128), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n336), .B(new_n329), .C1(new_n337), .C2(KEYINPUT23), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT80), .B(G110), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G125), .B(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT16), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT16), .ZN(new_n343));
  INV_X1    g157(.A(G140), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(G125), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(G146), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n341), .A2(new_n216), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n346), .ZN(new_n349));
  AOI21_X1  g163(.A(G146), .B1(new_n342), .B2(new_n345), .ZN(new_n350));
  OAI22_X1  g164(.A1(new_n349), .A2(new_n350), .B1(new_n334), .B2(new_n333), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n338), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n338), .A2(new_n352), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n353), .A2(G110), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n348), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G137), .ZN(new_n357));
  INV_X1    g171(.A(G953), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(G221), .A3(G234), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n357), .B(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G902), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n348), .B(new_n360), .C1(new_n351), .C2(new_n355), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n362), .A2(KEYINPUT25), .A3(new_n363), .A4(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G217), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(G234), .B2(new_n363), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(G902), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n362), .A2(new_n364), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G122), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT8), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G104), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n379), .A3(G104), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n382), .B2(KEYINPUT3), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n379), .A2(G104), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G101), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n384), .B2(new_n380), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n259), .A2(G119), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(G113), .B(new_n393), .C1(new_n260), .C2(new_n392), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n390), .A2(new_n264), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n390), .B1(new_n264), .B2(new_n394), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n378), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G125), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n227), .A2(G125), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT7), .ZN(new_n402));
  INV_X1    g216(.A(G224), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n397), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n401), .A2(new_n404), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n400), .A3(new_n405), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n408), .A2(new_n409), .B1(new_n402), .B2(new_n405), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n383), .A2(new_n386), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT85), .B(KEYINPUT4), .Z(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(G101), .A3(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n265), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(G101), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(KEYINPUT87), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n265), .A3(new_n414), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n390), .A2(new_n264), .A3(new_n394), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n418), .A2(new_n421), .A3(new_n377), .A4(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n411), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n377), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n422), .B1(new_n419), .B2(new_n420), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT87), .B1(new_n415), .B2(new_n417), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT6), .A3(new_n423), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n408), .A2(new_n409), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n431), .B(new_n425), .C1(new_n426), .C2(new_n427), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G210), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n424), .A2(new_n433), .A3(new_n435), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G214), .B1(G237), .B2(G902), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n256), .A2(G122), .A3(new_n257), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n259), .A2(G122), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT14), .ZN(new_n446));
  OAI21_X1  g260(.A(G107), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n444), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n379), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n224), .A2(G143), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n212), .A2(G128), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n193), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n448), .A2(KEYINPUT92), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n450), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n445), .A2(new_n447), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n224), .A2(G143), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(KEYINPUT13), .B2(new_n451), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n193), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT13), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT91), .B1(new_n452), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n453), .A2(new_n193), .ZN(new_n467));
  INV_X1    g281(.A(new_n450), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n449), .A2(new_n379), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n455), .A2(new_n459), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT9), .B(G234), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT81), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(new_n370), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n455), .A2(new_n459), .A3(new_n470), .A4(new_n474), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n363), .ZN(new_n479));
  INV_X1    g293(.A(G478), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(KEYINPUT15), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n479), .B(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n483));
  NOR2_X1   g297(.A1(G475), .A2(G902), .ZN(new_n484));
  XNOR2_X1  g298(.A(G113), .B(G122), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(G104), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n267), .A2(G143), .A3(G214), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G143), .B1(new_n267), .B2(G214), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT18), .A2(G131), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G237), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n358), .A3(G214), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n212), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n487), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT18), .A3(G131), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n341), .B(new_n216), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n492), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(G131), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n502), .A2(new_n350), .A3(new_n349), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n490), .A2(new_n504), .A3(new_n195), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT88), .B1(new_n496), .B2(G131), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n501), .A4(new_n500), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n486), .B(new_n499), .C1(new_n503), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n486), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n506), .A3(new_n500), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n341), .B(KEYINPUT19), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n216), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n346), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n499), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n483), .B(new_n484), .C1(new_n508), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT89), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n514), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n486), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n503), .A2(new_n507), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n509), .A3(new_n514), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n483), .A4(new_n484), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n484), .B1(new_n508), .B2(new_n515), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT20), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n517), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n509), .B1(new_n520), .B2(new_n514), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n363), .B1(new_n528), .B2(new_n508), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT90), .B(G475), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G952), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G953), .ZN(new_n534));
  NAND2_X1  g348(.A1(G234), .A2(G237), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n535), .A2(G902), .A3(G953), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT21), .B(G898), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n482), .A2(new_n532), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n473), .A2(G902), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G221), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n543), .B(KEYINPUT82), .Z(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n388), .A2(new_n389), .ZN(new_n546));
  AND4_X1   g360(.A1(new_n221), .A2(new_n218), .A3(new_n223), .A4(new_n225), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n221), .A2(new_n218), .A3(new_n223), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n215), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n549), .B2(KEYINPUT86), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT86), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n551), .A3(new_n215), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n546), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n390), .A2(new_n227), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n236), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT12), .B(new_n236), .C1(new_n553), .C2(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n553), .A2(KEYINPUT10), .ZN(new_n560));
  INV_X1    g374(.A(new_n236), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n390), .A2(KEYINPUT10), .A3(new_n227), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n417), .A2(new_n246), .A3(new_n414), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G140), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n358), .A2(G227), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT83), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n553), .A2(KEYINPUT10), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n563), .A2(new_n562), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n568), .B1(new_n572), .B2(new_n561), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n236), .B1(new_n570), .B2(new_n571), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n565), .A2(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G469), .ZN(new_n576));
  NAND2_X1  g390(.A1(G469), .A2(G902), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n564), .A2(new_n574), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n568), .A2(new_n579), .B1(new_n573), .B2(new_n559), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n580), .A2(G469), .A3(G902), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n545), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n441), .A2(new_n541), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n327), .A2(new_n376), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT93), .B(G101), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(G3));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n285), .B2(new_n296), .ZN(new_n588));
  INV_X1    g402(.A(G472), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n305), .A2(new_n363), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(KEYINPUT94), .A3(G472), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n582), .A2(new_n375), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n590), .A2(new_n306), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n440), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n437), .B2(new_n438), .ZN(new_n597));
  INV_X1    g411(.A(new_n539), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n480), .A2(G902), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT95), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT33), .B1(new_n478), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  AOI211_X1 g417(.A(KEYINPUT95), .B(new_n603), .C1(new_n476), .C2(new_n477), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n479), .A2(new_n480), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n532), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n599), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n595), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  INV_X1    g426(.A(new_n482), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n526), .A2(new_n516), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n531), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n599), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n595), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT96), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT35), .B(G107), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  NOR2_X1   g434(.A1(new_n361), .A2(KEYINPUT36), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n356), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n373), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT97), .B1(new_n372), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n371), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n367), .B2(new_n368), .ZN(new_n626));
  INV_X1    g440(.A(new_n623), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G469), .B1(new_n575), .B2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n579), .A2(new_n568), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n573), .A2(new_n559), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(G469), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n635), .A3(new_n363), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n544), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n540), .A2(new_n597), .A3(new_n630), .A4(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n638), .A2(new_n590), .A3(new_n306), .A4(new_n592), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  NAND3_X1  g455(.A1(new_n597), .A2(new_n630), .A3(new_n637), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n536), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n537), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n615), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n649), .A2(new_n482), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT75), .B1(new_n306), .B2(new_n307), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n187), .B(new_n298), .C1(new_n305), .C2(new_n188), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n325), .A2(G472), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n188), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n643), .B(new_n650), .C1(new_n653), .C2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  XOR2_X1   g472(.A(new_n439), .B(KEYINPUT38), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n482), .A2(new_n532), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n659), .A2(new_n596), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n626), .A2(new_n627), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n314), .A2(new_n280), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(G902), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n321), .A2(new_n280), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n589), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n297), .B2(KEYINPUT32), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n651), .B2(new_n652), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n661), .A2(new_n662), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT98), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n647), .B(KEYINPUT39), .Z(new_n672));
  OR2_X1    g486(.A1(new_n582), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT99), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n669), .A2(new_n670), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n671), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  NAND3_X1  g492(.A1(new_n607), .A2(new_n532), .A3(new_n647), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n643), .B(new_n680), .C1(new_n653), .C2(new_n656), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  OAI21_X1  g496(.A(G469), .B1(new_n580), .B2(G902), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n683), .A2(new_n636), .A3(new_n543), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n375), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n327), .A2(new_n609), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT100), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n687), .B(new_n689), .ZN(G15));
  NAND3_X1  g504(.A1(new_n327), .A2(new_n616), .A3(new_n686), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  INV_X1    g506(.A(new_n630), .ZN(new_n693));
  NOR4_X1   g507(.A1(new_n541), .A2(new_n685), .A3(new_n693), .A4(new_n441), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n327), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  NAND2_X1  g510(.A1(new_n660), .A2(KEYINPUT101), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n482), .A2(new_n532), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n598), .A3(new_n597), .A4(new_n684), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n302), .A2(new_n300), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n280), .B1(new_n315), .B2(new_n290), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n188), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n376), .B(new_n704), .C1(new_n588), .C2(new_n589), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(G122), .Z(G24));
  NAND2_X1  g521(.A1(new_n591), .A2(G472), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n704), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n680), .A2(new_n597), .A3(new_n684), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n709), .A2(new_n710), .A3(new_n662), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(G125), .Z(G27));
  AOI21_X1  g526(.A(new_n375), .B1(new_n309), .B2(new_n326), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n543), .B1(new_n578), .B2(new_n581), .ZN(new_n714));
  NOR4_X1   g528(.A1(new_n714), .A2(new_n679), .A3(new_n439), .A4(new_n596), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT32), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n306), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n654), .A3(new_n655), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n376), .A3(new_n715), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n713), .A2(new_n717), .B1(new_n721), .B2(KEYINPUT42), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  INV_X1    g537(.A(new_n714), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n439), .A2(new_n596), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n650), .A3(new_n725), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n375), .B(new_n726), .C1(new_n309), .C2(new_n326), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n193), .ZN(G36));
  AOI21_X1  g542(.A(new_n297), .B1(new_n708), .B2(new_n587), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n592), .ZN(new_n730));
  INV_X1    g544(.A(new_n662), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n532), .B1(new_n606), .B2(new_n605), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT43), .Z(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n725), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n575), .A2(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n575), .A2(KEYINPUT45), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(G469), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n577), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT102), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n581), .B1(new_n746), .B2(new_n747), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n543), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n672), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n741), .A2(new_n742), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G137), .ZN(G39));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n752), .B1(new_n756), .B2(KEYINPUT47), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n757), .B1(new_n752), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n656), .B1(new_n299), .B2(new_n308), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n679), .A2(new_n439), .A3(new_n376), .A4(new_n596), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n760), .A2(KEYINPUT105), .A3(new_n761), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n759), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n344), .ZN(G42));
  AND2_X1   g581(.A1(new_n683), .A2(new_n636), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT49), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(KEYINPUT49), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n375), .A2(new_n596), .A3(new_n544), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n732), .A2(new_n770), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(new_n309), .A3(new_n667), .A4(new_n659), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT106), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n734), .A2(new_n536), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n705), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n597), .A3(new_n684), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n725), .A2(new_n684), .ZN(new_n779));
  OR4_X1    g593(.A1(new_n375), .A2(new_n668), .A3(new_n644), .A4(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n778), .B(new_n534), .C1(new_n608), .C2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT113), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n776), .A2(new_n779), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n720), .A2(new_n376), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT48), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n659), .A2(new_n596), .A3(new_n684), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(KEYINPUT111), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n777), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT50), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n709), .A2(new_n662), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n795), .B1(new_n796), .B2(new_n783), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n780), .A2(new_n532), .A3(new_n607), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT112), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n777), .A2(new_n725), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n769), .A2(new_n545), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT110), .Z(new_n803));
  AOI21_X1  g617(.A(new_n801), .B1(new_n759), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n790), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n759), .B1(new_n545), .B2(new_n769), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n725), .A3(new_n777), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n797), .A3(KEYINPUT51), .A4(new_n799), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n789), .A2(new_n805), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n715), .A2(new_n708), .A3(new_n731), .A4(new_n704), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n693), .A2(new_n482), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n725), .A3(new_n637), .A4(new_n649), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n811), .B1(new_n760), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT108), .B1(new_n814), .B2(new_n727), .ZN(new_n815));
  INV_X1    g629(.A(new_n726), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n713), .A2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n812), .A2(new_n637), .A3(new_n649), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n327), .A2(new_n725), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n817), .A2(new_n819), .A3(new_n820), .A4(new_n811), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n706), .B1(new_n327), .B2(new_n694), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n687), .A3(new_n691), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n713), .A2(new_n717), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n721), .A2(KEYINPUT42), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT107), .ZN(new_n829));
  INV_X1    g643(.A(new_n532), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n482), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n599), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n639), .B(new_n829), .C1(new_n594), .C2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n584), .A3(new_n610), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n729), .A2(new_n832), .A3(new_n592), .A4(new_n593), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n829), .B1(new_n836), .B2(new_n639), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n822), .A2(new_n828), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n711), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n597), .A2(new_n700), .A3(new_n724), .A4(new_n647), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n668), .A2(new_n841), .A3(new_n662), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n657), .A2(new_n681), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n642), .B1(new_n309), .B2(new_n326), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n711), .B1(new_n846), .B2(new_n650), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(KEYINPUT52), .A3(new_n681), .A4(new_n842), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT53), .B1(new_n839), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n722), .A2(new_n687), .A3(new_n691), .A4(new_n823), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n815), .B2(new_n821), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n845), .A2(new_n848), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n838), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n852), .A2(new_n854), .A3(new_n838), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT53), .B1(new_n854), .B2(KEYINPUT109), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n859), .B(new_n860), .Z(new_n861));
  OAI21_X1  g675(.A(new_n858), .B1(new_n861), .B2(new_n857), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n810), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(G952), .A2(G953), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n775), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT115), .ZN(G75));
  NOR2_X1   g680(.A1(new_n358), .A2(G952), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n429), .A2(new_n432), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(new_n430), .ZN(new_n869));
  XNOR2_X1  g683(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n856), .A2(new_n363), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(G210), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n872), .B(KEYINPUT117), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n436), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n871), .A2(new_n874), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n867), .B(new_n875), .C1(new_n877), .C2(new_n878), .ZN(G51));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n850), .A2(new_n855), .A3(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n858), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n856), .A2(KEYINPUT118), .A3(new_n857), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n577), .B(KEYINPUT57), .Z(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n634), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(KEYINPUT119), .ZN(new_n887));
  INV_X1    g701(.A(new_n745), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n888), .B2(new_n876), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(KEYINPUT119), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n867), .B1(new_n889), .B2(new_n890), .ZN(G54));
  NAND3_X1  g705(.A1(new_n876), .A2(KEYINPUT58), .A3(G475), .ZN(new_n892));
  INV_X1    g706(.A(new_n522), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n867), .ZN(G60));
  OR2_X1    g710(.A1(new_n602), .A2(new_n604), .ZN(new_n897));
  NAND2_X1  g711(.A1(G478), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT59), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n882), .A2(new_n897), .A3(new_n883), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n867), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n900), .A2(KEYINPUT120), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT120), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n897), .B1(new_n862), .B2(new_n899), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT60), .Z(new_n907));
  NAND3_X1  g721(.A1(new_n850), .A2(new_n855), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n362), .A2(new_n364), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n867), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n850), .A2(new_n855), .A3(new_n622), .A4(new_n907), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(KEYINPUT61), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n908), .A2(new_n909), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n901), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT122), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n918), .A3(new_n911), .ZN(new_n919));
  XOR2_X1   g733(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n920));
  AOI21_X1  g734(.A(new_n913), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n911), .B1(new_n910), .B2(new_n917), .ZN(new_n922));
  AOI211_X1 g736(.A(KEYINPUT122), .B(new_n867), .C1(new_n908), .C2(new_n909), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n913), .B(new_n920), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n912), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(KEYINPUT124), .B(new_n912), .C1(new_n921), .C2(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(G66));
  OAI21_X1  g744(.A(G953), .B1(new_n538), .B2(new_n403), .ZN(new_n931));
  INV_X1    g745(.A(new_n838), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n824), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n933), .B2(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n868), .B1(G898), .B2(new_n358), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G69));
  NAND4_X1  g750(.A1(new_n753), .A2(new_n597), .A3(new_n700), .A4(new_n785), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n722), .A3(new_n817), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n847), .A2(new_n681), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n766), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n754), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT127), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n943), .A3(new_n754), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n358), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n282), .B(KEYINPUT125), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n511), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n945), .B(new_n947), .C1(new_n645), .C2(new_n358), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n831), .A2(new_n608), .ZN(new_n949));
  NOR4_X1   g763(.A1(new_n673), .A2(new_n949), .A3(new_n596), .A4(new_n439), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n766), .B1(new_n713), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n677), .A2(new_n681), .A3(new_n847), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n951), .A2(new_n754), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n947), .B1(new_n955), .B2(new_n358), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n948), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n358), .B1(G227), .B2(G900), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  INV_X1    g778(.A(new_n933), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n955), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n665), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n867), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n266), .A2(new_n271), .A3(new_n279), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n665), .A2(new_n969), .A3(new_n964), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n861), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n942), .A2(new_n933), .A3(new_n944), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n972), .B2(new_n964), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n971), .A2(new_n973), .ZN(G57));
endmodule


