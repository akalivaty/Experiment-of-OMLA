//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n449));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  INV_X1    g026(.A(new_n450), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n452), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n452), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n456), .A2(G2106), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n466), .A2(G101), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n466), .B1(new_n476), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n467), .B2(new_n468), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(new_n496), .C1(new_n468), .C2(new_n467), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n491), .B1(new_n495), .B2(new_n497), .ZN(G164));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT68), .A2(G651), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT68), .A2(KEYINPUT6), .A3(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n501), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  INV_X1    g086(.A(new_n508), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT6), .B1(KEYINPUT68), .B2(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n510), .A2(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n504), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  INV_X1    g093(.A(new_n510), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n521), .B(new_n523), .C1(new_n514), .C2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n520), .A2(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n527), .A2(new_n503), .B1(new_n510), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n507), .B2(new_n508), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n531), .A2(G52), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n503), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(G43), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n509), .A2(new_n501), .A3(G81), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n536), .A2(KEYINPUT69), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(KEYINPUT69), .B1(new_n536), .B2(new_n537), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n501), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n503), .ZN(new_n550));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(new_n500), .ZN(new_n552));
  NOR2_X1   g127(.A1(KEYINPUT5), .A2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n556), .A2(KEYINPUT71), .A3(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(KEYINPUT70), .A2(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n514), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n531), .A2(KEYINPUT70), .A3(new_n561), .A4(G53), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n560), .A2(new_n562), .B1(new_n519), .B2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  NAND2_X1  g141(.A1(new_n519), .A2(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n531), .A2(G49), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  INV_X1    g146(.A(G73), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n554), .A2(new_n571), .B1(new_n572), .B2(new_n530), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n531), .B2(G48), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n509), .A2(new_n501), .A3(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(new_n519), .A2(G85), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  XOR2_X1   g153(.A(KEYINPUT72), .B(G47), .Z(new_n579));
  OAI221_X1 g154(.A(new_n577), .B1(new_n503), .B2(new_n578), .C1(new_n514), .C2(new_n579), .ZN(G290));
  INV_X1    g155(.A(KEYINPUT10), .ZN(new_n581));
  INV_X1    g156(.A(G92), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n510), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n509), .A2(new_n501), .A3(KEYINPUT10), .A4(G92), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n514), .A2(KEYINPUT73), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n531), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n588), .A3(G54), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n501), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n503), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n585), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n593), .B2(G171), .ZN(G284));
  OAI21_X1  g170(.A(new_n594), .B1(new_n593), .B2(G171), .ZN(G321));
  NAND2_X1  g171(.A1(G299), .A2(new_n593), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n593), .B2(G168), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(new_n593), .B2(G168), .ZN(G280));
  INV_X1    g174(.A(new_n592), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT74), .B(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(G860), .B2(new_n601), .ZN(G148));
  NAND2_X1  g177(.A1(new_n541), .A2(new_n593), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n601), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n605), .B2(new_n593), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g182(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT12), .Z(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT13), .Z(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT75), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n478), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n480), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n466), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2096), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n611), .B2(new_n610), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n613), .A2(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2443), .B(G2446), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT77), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n636), .A2(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT78), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  AOI21_X1  g220(.A(KEYINPUT18), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT79), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(G2072), .A2(G2078), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n444), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT80), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n659), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n660), .A2(KEYINPUT20), .A3(new_n659), .ZN(new_n665));
  OAI221_X1 g240(.A(new_n661), .B1(new_n659), .B2(new_n657), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n672), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(G229));
  MUX2_X1   g250(.A(G6), .B(G305), .S(G16), .Z(new_n676));
  XOR2_X1   g251(.A(KEYINPUT32), .B(G1981), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n679));
  NOR2_X1   g254(.A1(G16), .A2(G23), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT84), .Z(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(G288), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT85), .Z(new_n684));
  XOR2_X1   g259(.A(KEYINPUT33), .B(G1976), .Z(new_n685));
  AOI22_X1  g260(.A1(new_n678), .A2(new_n679), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n678), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(G22), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G166), .B2(new_n682), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G1971), .Z(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n684), .B2(new_n685), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n687), .A2(KEYINPUT34), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(KEYINPUT34), .B1(new_n687), .B2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(G25), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n478), .A2(G131), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n480), .A2(G119), .ZN(new_n700));
  OR2_X1    g275(.A1(G95), .A2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n701), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n698), .B1(new_n704), .B2(new_n697), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT35), .B(G1991), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G24), .B(G290), .S(G16), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT82), .B(G1986), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n692), .A2(new_n693), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT36), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n682), .A2(G20), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT23), .ZN(new_n714));
  INV_X1    g289(.A(G299), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n682), .ZN(new_n716));
  INV_X1    g291(.A(G1956), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n697), .A2(G35), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n697), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT29), .ZN(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G168), .A2(new_n682), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n682), .B2(G21), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G171), .A2(new_n682), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G5), .B2(new_n682), .ZN(new_n728));
  INV_X1    g303(.A(G1961), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n726), .A2(G1966), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n728), .ZN(new_n731));
  INV_X1    g306(.A(G1966), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n731), .A2(G1961), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n723), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT31), .B(G11), .Z(new_n735));
  INV_X1    g310(.A(G28), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(KEYINPUT30), .ZN(new_n737));
  AOI21_X1  g312(.A(G29), .B1(new_n736), .B2(KEYINPUT30), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n697), .ZN(new_n740));
  INV_X1    g315(.A(G34), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(KEYINPUT24), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n697), .B1(KEYINPUT24), .B2(new_n741), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(KEYINPUT91), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(KEYINPUT91), .B2(new_n743), .ZN(new_n745));
  NAND2_X1  g320(.A1(G160), .A2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n739), .B1(new_n618), .B2(new_n740), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n748), .B2(new_n747), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n697), .A2(G27), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n697), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G2078), .Z(new_n753));
  XOR2_X1   g328(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT92), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n478), .A2(G141), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n480), .A2(G129), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n756), .A2(new_n758), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G32), .B(new_n761), .S(G29), .Z(new_n762));
  XOR2_X1   g337(.A(KEYINPUT27), .B(G1996), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT94), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n762), .B(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n750), .A2(new_n753), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n740), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n480), .A2(G128), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT87), .Z(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  INV_X1    g346(.A(G116), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G140), .B2(new_n478), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n768), .B1(new_n775), .B2(G29), .ZN(new_n776));
  INV_X1    g351(.A(G2067), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n734), .A2(new_n766), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G33), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(G29), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT88), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT25), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n478), .A2(G139), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT89), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT3), .B(G2104), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G127), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT90), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n466), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n787), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n781), .B1(new_n795), .B2(G29), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2072), .ZN(new_n797));
  NOR2_X1   g372(.A1(G16), .A2(G19), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n542), .B2(G16), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT86), .B(G1341), .Z(new_n800));
  XOR2_X1   g375(.A(new_n799), .B(new_n800), .Z(new_n801));
  NOR2_X1   g376(.A1(G4), .A2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n600), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1348), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AND4_X1   g380(.A1(new_n718), .A2(new_n779), .A3(new_n797), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n712), .A2(new_n806), .ZN(G150));
  INV_X1    g382(.A(G150), .ZN(G311));
  NAND2_X1  g383(.A1(new_n531), .A2(G55), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n503), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT95), .B(G93), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n510), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G860), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n600), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  INV_X1    g394(.A(new_n814), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n541), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n814), .B(new_n535), .C1(new_n540), .C2(new_n539), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n819), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT96), .Z(new_n827));
  OAI21_X1  g402(.A(new_n815), .B1(new_n824), .B2(new_n825), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n817), .B1(new_n827), .B2(new_n828), .ZN(G145));
  XNOR2_X1  g404(.A(G160), .B(new_n484), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT97), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n618), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n775), .B(new_n761), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(G164), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(G164), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n795), .A2(KEYINPUT98), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n795), .A2(KEYINPUT98), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n480), .A2(G130), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n466), .A2(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G142), .B2(new_n478), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(new_n609), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n703), .ZN(new_n847));
  OAI211_X1 g422(.A(KEYINPUT98), .B(new_n795), .C1(new_n835), .C2(new_n836), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n840), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n847), .B1(new_n840), .B2(new_n848), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n833), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n851), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n853), .A2(new_n832), .A3(new_n849), .ZN(new_n854));
  INV_X1    g429(.A(G37), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g432(.A1(new_n820), .A2(new_n593), .ZN(new_n858));
  XOR2_X1   g433(.A(G290), .B(G305), .Z(new_n859));
  AND3_X1   g434(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G303), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n859), .B(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n600), .A2(G299), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n592), .A2(new_n558), .A3(new_n563), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT101), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n866), .A2(new_n867), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n600), .A2(KEYINPUT99), .A3(G299), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(KEYINPUT101), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n871), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n823), .B(new_n604), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n882));
  INV_X1    g457(.A(new_n875), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT100), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n865), .A2(new_n881), .A3(new_n882), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT103), .B1(new_n887), .B2(new_n864), .ZN(new_n888));
  INV_X1    g463(.A(new_n885), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n879), .A2(new_n880), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n864), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT104), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n893), .A3(new_n864), .ZN(new_n894));
  AND4_X1   g469(.A1(new_n886), .A2(new_n888), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n858), .B1(new_n895), .B2(new_n593), .ZN(G295));
  OAI21_X1  g471(.A(new_n858), .B1(new_n895), .B2(new_n593), .ZN(G331));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n821), .A2(new_n822), .A3(G301), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G301), .B1(new_n821), .B2(new_n822), .ZN(new_n902));
  OAI21_X1  g477(.A(G286), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(G168), .A3(new_n900), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n875), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n903), .A2(new_n905), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n878), .B2(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(KEYINPUT105), .ZN(new_n909));
  INV_X1    g484(.A(new_n862), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(KEYINPUT105), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n908), .B2(new_n862), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n899), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n868), .A2(KEYINPUT41), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n883), .B2(KEYINPUT41), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n903), .A2(new_n905), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n906), .A2(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n906), .A2(new_n915), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n910), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n913), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n898), .B1(new_n914), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n898), .B1(new_n922), .B2(KEYINPUT43), .ZN(new_n925));
  INV_X1    g500(.A(new_n911), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n910), .B1(new_n908), .B2(KEYINPUT105), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n899), .B(new_n913), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n925), .A2(KEYINPUT107), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT107), .B1(new_n925), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(G397));
  INV_X1    g506(.A(KEYINPUT57), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n558), .A2(new_n563), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n558), .B2(new_n563), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT50), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  INV_X1    g513(.A(new_n497), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n496), .B1(new_n788), .B2(new_n493), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n937), .B(new_n938), .C1(new_n941), .C2(new_n491), .ZN(new_n942));
  INV_X1    g517(.A(G125), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n476), .B2(new_n477), .ZN(new_n944));
  INV_X1    g519(.A(new_n470), .ZN(new_n945));
  OAI21_X1  g520(.A(G2105), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(G40), .A3(new_n473), .A4(new_n472), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(G160), .A2(KEYINPUT108), .A3(G40), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n936), .A2(new_n942), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n717), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT108), .B1(G160), .B2(G40), .ZN(new_n953));
  INV_X1    g528(.A(G40), .ZN(new_n954));
  NOR4_X1   g529(.A1(new_n471), .A2(new_n474), .A3(new_n948), .A4(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G164), .B2(G1384), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT45), .B(new_n938), .C1(new_n941), .C2(new_n491), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT56), .B(G2072), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n956), .A2(new_n958), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n935), .B1(new_n952), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(G164), .A2(G1384), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(new_n949), .A3(new_n950), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1348), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n965), .A2(new_n777), .B1(new_n951), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(new_n592), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n952), .A2(new_n961), .A3(new_n935), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n951), .A2(new_n966), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n956), .A2(new_n777), .A3(new_n963), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n585), .A2(KEYINPUT120), .A3(new_n591), .A4(new_n589), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n973), .A2(KEYINPUT60), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n600), .A2(KEYINPUT120), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT117), .B(G1996), .Z(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n956), .A2(new_n958), .A3(new_n959), .A4(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT58), .B(G1341), .Z(new_n980));
  NAND2_X1  g555(.A1(new_n964), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n541), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n983));
  AOI22_X1  g558(.A1(new_n975), .A2(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n933), .A2(new_n934), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n495), .A2(new_n497), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n486), .A2(new_n490), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n937), .B1(new_n988), .B2(new_n938), .ZN(new_n989));
  AOI211_X1 g564(.A(KEYINPUT50), .B(G1384), .C1(new_n986), .C2(new_n987), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G1956), .B1(new_n991), .B2(new_n956), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n958), .A2(new_n959), .A3(new_n949), .A4(new_n950), .ZN(new_n993));
  INV_X1    g568(.A(new_n960), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n985), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT119), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT61), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n999), .A3(new_n969), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n979), .A2(new_n981), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n542), .ZN(new_n1002));
  NOR2_X1   g577(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n1005));
  INV_X1    g580(.A(new_n976), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1005), .B(new_n1006), .C1(new_n967), .C2(KEYINPUT60), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n984), .A2(new_n1000), .A3(new_n1004), .A4(new_n1007), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n952), .A2(new_n961), .A3(new_n935), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(new_n962), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n997), .A2(new_n998), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n999), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n970), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT111), .B(G8), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G168), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n951), .B2(G2084), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n991), .A2(KEYINPUT116), .A3(new_n748), .A4(new_n956), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n993), .A2(new_n732), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n1020), .B2(G8), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1014), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(G286), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1015), .A2(KEYINPUT51), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1023), .A2(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G303), .A2(G8), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT55), .ZN(new_n1030));
  AOI21_X1  g605(.A(G2090), .B1(new_n951), .B2(KEYINPUT115), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n991), .A2(new_n1032), .A3(new_n956), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT109), .B(G1971), .Z(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1031), .A2(new_n1033), .B1(new_n993), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1030), .B1(new_n1036), .B2(new_n1014), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT45), .B1(new_n988), .B2(new_n938), .ZN(new_n1038));
  AOI211_X1 g613(.A(new_n957), .B(G1384), .C1(new_n986), .C2(new_n987), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1034), .B1(new_n1040), .B2(new_n956), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n951), .A2(G2090), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT110), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1029), .B(KEYINPUT55), .Z(new_n1044));
  NAND3_X1  g619(.A1(new_n991), .A2(new_n722), .A3(new_n956), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n993), .A2(new_n1035), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1043), .A2(G8), .A3(new_n1044), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n574), .A2(new_n1050), .A3(new_n1051), .A4(new_n575), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n571), .B1(new_n499), .B2(new_n500), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n572), .A2(new_n530), .ZN(new_n1054));
  OAI21_X1  g629(.A(G651), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n531), .A2(G48), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(new_n1051), .A3(new_n1056), .A4(new_n575), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT112), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1052), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G305), .A2(G1981), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1059), .A2(KEYINPUT49), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT49), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n964), .A2(new_n1024), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n860), .A2(G1976), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n964), .A2(new_n1065), .A3(new_n1024), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n964), .A2(new_n1065), .A3(new_n1069), .A4(new_n1024), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1037), .A2(new_n1049), .A3(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n993), .B2(G2078), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n951), .A2(new_n729), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1075), .A2(G2078), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1040), .A2(new_n956), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G171), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n947), .A2(new_n1075), .A3(G2078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1040), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1076), .A2(G301), .A3(new_n1077), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1074), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1073), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1076), .A2(new_n1077), .A3(new_n1083), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G171), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1076), .A2(G301), .A3(new_n1079), .A4(new_n1077), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(KEYINPUT54), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1088), .A2(KEYINPUT122), .A3(KEYINPUT54), .A4(new_n1089), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1013), .A2(new_n1028), .A3(new_n1086), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT63), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1020), .A2(G168), .A3(new_n1024), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n1073), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1096), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1043), .A2(G8), .A3(new_n1048), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n1030), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1099), .A2(new_n1101), .A3(new_n1049), .A4(new_n1072), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1049), .A2(new_n1064), .A3(new_n1071), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n860), .A2(new_n1068), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1059), .B1(new_n1064), .B2(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1106), .A2(KEYINPUT114), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1063), .B(KEYINPUT113), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1106), .B2(KEYINPUT114), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1104), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1095), .A2(new_n1103), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT123), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1095), .A2(new_n1113), .A3(new_n1103), .A4(new_n1110), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1073), .A2(new_n1081), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1028), .B2(KEYINPUT62), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1115), .B(KEYINPUT124), .C1(new_n1028), .C2(KEYINPUT62), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1112), .A2(new_n1114), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n956), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(new_n958), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n775), .B(new_n777), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n761), .B(G1996), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n704), .A2(new_n706), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n704), .A2(new_n706), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(G290), .B(G1986), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1122), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G290), .A2(G1986), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1137));
  XOR2_X1   g712(.A(new_n1136), .B(new_n1137), .Z(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n1131), .B2(new_n1124), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1123), .A2(G1996), .A3(new_n958), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT46), .Z(new_n1141));
  OAI21_X1  g716(.A(new_n1124), .B1(new_n1126), .B2(new_n761), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT47), .Z(new_n1144));
  XNOR2_X1  g719(.A(new_n1129), .B(KEYINPUT125), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1128), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(G2067), .B2(new_n775), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n1139), .B(new_n1144), .C1(new_n1124), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1134), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g724(.A1(new_n914), .A2(new_n923), .ZN(new_n1151));
  OR2_X1    g725(.A1(G227), .A2(new_n464), .ZN(new_n1152));
  AOI21_X1  g726(.A(new_n1152), .B1(new_n636), .B2(new_n638), .ZN(new_n1153));
  AOI22_X1  g727(.A1(new_n1153), .A2(KEYINPUT127), .B1(new_n673), .B2(new_n674), .ZN(new_n1154));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n1155));
  OAI21_X1  g729(.A(new_n1155), .B1(G401), .B2(new_n1152), .ZN(new_n1156));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1156), .A3(new_n856), .ZN(new_n1157));
  NOR2_X1   g731(.A1(new_n1151), .A2(new_n1157), .ZN(G308));
  OR2_X1    g732(.A1(new_n1151), .A2(new_n1157), .ZN(G225));
endmodule


