

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U323 ( .A(n304), .B(n303), .ZN(n309) );
  XNOR2_X1 U324 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U325 ( .A(n493), .B(KEYINPUT28), .Z(n527) );
  XNOR2_X1 U326 ( .A(n415), .B(n414), .ZN(n535) );
  AND2_X1 U327 ( .A1(G225GAT), .A2(G233GAT), .ZN(n291) );
  AND2_X1 U328 ( .A1(G226GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U329 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n467) );
  XNOR2_X1 U330 ( .A(n446), .B(n291), .ZN(n296) );
  XNOR2_X1 U331 ( .A(n468), .B(n467), .ZN(n475) );
  XNOR2_X1 U332 ( .A(n296), .B(n325), .ZN(n297) );
  NOR2_X1 U333 ( .A1(n450), .A2(n583), .ZN(n451) );
  XNOR2_X1 U334 ( .A(n407), .B(n292), .ZN(n408) );
  XNOR2_X1 U335 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U336 ( .A(n409), .B(n408), .ZN(n413) );
  XNOR2_X1 U337 ( .A(n329), .B(n328), .ZN(n472) );
  XNOR2_X1 U338 ( .A(n452), .B(KEYINPUT38), .ZN(n517) );
  XNOR2_X1 U339 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U340 ( .A(n453), .B(G29GAT), .ZN(n454) );
  XNOR2_X1 U341 ( .A(n486), .B(n485), .ZN(G1341GAT) );
  XNOR2_X1 U342 ( .A(n455), .B(n454), .ZN(G1328GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT6), .B(KEYINPUT85), .Z(n294) );
  XNOR2_X1 U344 ( .A(G85GAT), .B(KEYINPUT86), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U346 ( .A(G29GAT), .B(G134GAT), .Z(n446) );
  XNOR2_X1 U347 ( .A(G120GAT), .B(G148GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n295), .B(G57GAT), .ZN(n325) );
  XOR2_X1 U349 ( .A(n298), .B(n297), .Z(n304) );
  XOR2_X1 U350 ( .A(G113GAT), .B(G1GAT), .Z(n334) );
  XOR2_X1 U351 ( .A(KEYINPUT0), .B(G127GAT), .Z(n376) );
  XNOR2_X1 U352 ( .A(n334), .B(n376), .ZN(n302) );
  XOR2_X1 U353 ( .A(KEYINPUT87), .B(KEYINPUT5), .Z(n300) );
  XNOR2_X1 U354 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U356 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n305), .B(KEYINPUT2), .ZN(n306) );
  XOR2_X1 U358 ( .A(n306), .B(KEYINPUT83), .Z(n308) );
  XNOR2_X1 U359 ( .A(G141GAT), .B(G162GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n398) );
  XNOR2_X1 U361 ( .A(n309), .B(n398), .ZN(n430) );
  XOR2_X1 U362 ( .A(KEYINPUT88), .B(n430), .Z(n417) );
  XOR2_X1 U363 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n311) );
  NAND2_X1 U364 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n313) );
  INV_X1 U366 ( .A(KEYINPUT69), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n322) );
  INV_X1 U368 ( .A(G92GAT), .ZN(n314) );
  NAND2_X1 U369 ( .A1(n314), .A2(G64GAT), .ZN(n317) );
  INV_X1 U370 ( .A(G64GAT), .ZN(n315) );
  NAND2_X1 U371 ( .A1(n315), .A2(G92GAT), .ZN(n316) );
  NAND2_X1 U372 ( .A1(n317), .A2(n316), .ZN(n319) );
  XNOR2_X1 U373 ( .A(G176GAT), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n404) );
  XNOR2_X1 U375 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n320), .B(KEYINPUT68), .ZN(n353) );
  XNOR2_X1 U377 ( .A(n404), .B(n353), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U379 ( .A(n323), .B(KEYINPUT33), .Z(n329) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(G78GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n324), .B(KEYINPUT70), .ZN(n394) );
  XOR2_X1 U382 ( .A(n394), .B(n325), .Z(n327) );
  XOR2_X1 U383 ( .A(G99GAT), .B(G85GAT), .Z(n445) );
  XNOR2_X1 U384 ( .A(n445), .B(KEYINPUT31), .ZN(n326) );
  INV_X1 U385 ( .A(n472), .ZN(n577) );
  XOR2_X1 U386 ( .A(G197GAT), .B(G141GAT), .Z(n331) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(G29GAT), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n344) );
  XOR2_X1 U389 ( .A(G43GAT), .B(G50GAT), .Z(n333) );
  XNOR2_X1 U390 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n438) );
  XOR2_X1 U392 ( .A(n438), .B(n334), .Z(n336) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U395 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n338) );
  XNOR2_X1 U396 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U398 ( .A(n340), .B(n339), .Z(n342) );
  XOR2_X1 U399 ( .A(G22GAT), .B(G15GAT), .Z(n359) );
  XOR2_X1 U400 ( .A(G169GAT), .B(G8GAT), .Z(n403) );
  XNOR2_X1 U401 ( .A(n359), .B(n403), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n540) );
  NAND2_X1 U404 ( .A1(n577), .A2(n540), .ZN(n506) );
  XOR2_X1 U405 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n346) );
  XNOR2_X1 U406 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n367) );
  XOR2_X1 U408 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n348) );
  XNOR2_X1 U409 ( .A(G1GAT), .B(KEYINPUT72), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U411 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n350) );
  XNOR2_X1 U412 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U414 ( .A(n352), .B(n351), .Z(n365) );
  XOR2_X1 U415 ( .A(n353), .B(G64GAT), .Z(n355) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n363) );
  XOR2_X1 U418 ( .A(G57GAT), .B(G78GAT), .Z(n357) );
  XNOR2_X1 U419 ( .A(G127GAT), .B(G155GAT), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U421 ( .A(n358), .B(G211GAT), .Z(n361) );
  XNOR2_X1 U422 ( .A(n359), .B(G183GAT), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U426 ( .A(n367), .B(n366), .Z(n580) );
  XOR2_X1 U427 ( .A(G120GAT), .B(KEYINPUT81), .Z(n369) );
  XNOR2_X1 U428 ( .A(G113GAT), .B(KEYINPUT20), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n383) );
  XOR2_X1 U430 ( .A(G134GAT), .B(G99GAT), .Z(n371) );
  XNOR2_X1 U431 ( .A(G43GAT), .B(G190GAT), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U433 ( .A(G176GAT), .B(KEYINPUT79), .Z(n373) );
  XNOR2_X1 U434 ( .A(G169GAT), .B(KEYINPUT80), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U436 ( .A(n375), .B(n374), .Z(n381) );
  XOR2_X1 U437 ( .A(G71GAT), .B(n376), .Z(n378) );
  NAND2_X1 U438 ( .A1(G227GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U440 ( .A(G15GAT), .B(n379), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U443 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n385) );
  XNOR2_X1 U444 ( .A(KEYINPUT82), .B(G183GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U446 ( .A(KEYINPUT19), .B(n386), .ZN(n414) );
  XOR2_X1 U447 ( .A(n387), .B(n414), .Z(n421) );
  XOR2_X1 U448 ( .A(KEYINPUT24), .B(KEYINPUT84), .Z(n389) );
  XNOR2_X1 U449 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n402) );
  XNOR2_X1 U451 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n390), .B(G211GAT), .ZN(n411) );
  XOR2_X1 U453 ( .A(G218GAT), .B(n411), .Z(n392) );
  XNOR2_X1 U454 ( .A(G50GAT), .B(G148GAT), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U456 ( .A(n393), .B(KEYINPUT22), .Z(n400) );
  XOR2_X1 U457 ( .A(n394), .B(G204GAT), .Z(n396) );
  NAND2_X1 U458 ( .A1(G228GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U462 ( .A(n402), .B(n401), .Z(n493) );
  XOR2_X1 U463 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U464 ( .A(KEYINPUT89), .B(KEYINPUT91), .Z(n406) );
  XNOR2_X1 U465 ( .A(KEYINPUT72), .B(KEYINPUT90), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U467 ( .A(G36GAT), .B(G190GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n410), .B(G218GAT), .ZN(n437) );
  XNOR2_X1 U469 ( .A(n411), .B(n437), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n535), .B(KEYINPUT27), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n416), .B(KEYINPUT92), .ZN(n426) );
  NAND2_X1 U473 ( .A1(n426), .A2(n417), .ZN(n418) );
  XOR2_X1 U474 ( .A(KEYINPUT93), .B(n418), .Z(n478) );
  NOR2_X1 U475 ( .A1(n527), .A2(n478), .ZN(n419) );
  NAND2_X1 U476 ( .A1(n421), .A2(n419), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n420), .B(KEYINPUT94), .ZN(n432) );
  INV_X1 U478 ( .A(n421), .ZN(n537) );
  NAND2_X1 U479 ( .A1(n537), .A2(n535), .ZN(n422) );
  NAND2_X1 U480 ( .A1(n422), .A2(n493), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n423), .B(KEYINPUT95), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n424), .B(KEYINPUT25), .ZN(n428) );
  NOR2_X1 U483 ( .A1(n537), .A2(n493), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n425), .B(KEYINPUT26), .ZN(n570) );
  NAND2_X1 U485 ( .A1(n426), .A2(n570), .ZN(n427) );
  NAND2_X1 U486 ( .A1(n428), .A2(n427), .ZN(n429) );
  NAND2_X1 U487 ( .A1(n430), .A2(n429), .ZN(n431) );
  NAND2_X1 U488 ( .A1(n432), .A2(n431), .ZN(n504) );
  NAND2_X1 U489 ( .A1(n580), .A2(n504), .ZN(n433) );
  XOR2_X1 U490 ( .A(KEYINPUT99), .B(n433), .Z(n450) );
  XOR2_X1 U491 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n435) );
  NAND2_X1 U492 ( .A1(G232GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U494 ( .A(n436), .B(KEYINPUT9), .Z(n440) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U497 ( .A(G92GAT), .B(KEYINPUT64), .Z(n442) );
  XNOR2_X1 U498 ( .A(G162GAT), .B(G106GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U500 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U502 ( .A(n448), .B(n447), .Z(n547) );
  XNOR2_X1 U503 ( .A(KEYINPUT36), .B(KEYINPUT98), .ZN(n449) );
  XOR2_X1 U504 ( .A(n547), .B(n449), .Z(n583) );
  XNOR2_X1 U505 ( .A(n451), .B(KEYINPUT37), .ZN(n456) );
  NOR2_X1 U506 ( .A1(n506), .A2(n456), .ZN(n452) );
  NAND2_X1 U507 ( .A1(n417), .A2(n517), .ZN(n455) );
  XOR2_X1 U508 ( .A(KEYINPUT39), .B(KEYINPUT100), .Z(n453) );
  INV_X1 U509 ( .A(n540), .ZN(n572) );
  XOR2_X1 U510 ( .A(KEYINPUT41), .B(n472), .Z(n555) );
  NAND2_X1 U511 ( .A1(n572), .A2(n555), .ZN(n520) );
  NOR2_X1 U512 ( .A1(n520), .A2(n456), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n457), .B(KEYINPUT104), .ZN(n538) );
  NAND2_X1 U514 ( .A1(n527), .A2(n538), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n459) );
  XNOR2_X1 U516 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n461), .B(n460), .ZN(G1339GAT) );
  INV_X1 U519 ( .A(KEYINPUT48), .ZN(n477) );
  XOR2_X1 U520 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n463) );
  NAND2_X1 U521 ( .A1(n540), .A2(n555), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n463), .B(n462), .ZN(n464) );
  AND2_X1 U523 ( .A1(n464), .A2(n580), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT110), .ZN(n466) );
  INV_X1 U525 ( .A(n547), .ZN(n560) );
  NAND2_X1 U526 ( .A1(n466), .A2(n560), .ZN(n468) );
  XOR2_X1 U527 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n470) );
  NOR2_X1 U528 ( .A1(n580), .A2(n583), .ZN(n469) );
  XOR2_X1 U529 ( .A(n470), .B(n469), .Z(n471) );
  NOR2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n473), .A2(n572), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n477), .B(n476), .ZN(n488) );
  NOR2_X1 U534 ( .A1(n478), .A2(n488), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n479), .B(KEYINPUT112), .ZN(n551) );
  NAND2_X1 U536 ( .A1(n551), .A2(n537), .ZN(n480) );
  XOR2_X1 U537 ( .A(n480), .B(KEYINPUT113), .Z(n481) );
  NOR2_X1 U538 ( .A1(n481), .A2(n527), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n482), .B(KEYINPUT114), .ZN(n548) );
  NAND2_X1 U540 ( .A1(n548), .A2(n555), .ZN(n486) );
  XOR2_X1 U541 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n484) );
  INV_X1 U542 ( .A(G120GAT), .ZN(n483) );
  INV_X1 U543 ( .A(G190GAT), .ZN(n500) );
  XNOR2_X1 U544 ( .A(n535), .B(KEYINPUT119), .ZN(n487) );
  NOR2_X1 U545 ( .A1(n488), .A2(n487), .ZN(n491) );
  XNOR2_X1 U546 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(KEYINPUT121), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(n492) );
  NOR2_X1 U549 ( .A1(n492), .A2(n417), .ZN(n571) );
  NAND2_X1 U550 ( .A1(n493), .A2(n571), .ZN(n494) );
  XNOR2_X1 U551 ( .A(n494), .B(KEYINPUT55), .ZN(n495) );
  NAND2_X1 U552 ( .A1(n495), .A2(n537), .ZN(n496) );
  XNOR2_X1 U553 ( .A(n496), .B(KEYINPUT122), .ZN(n568) );
  NOR2_X1 U554 ( .A1(n560), .A2(n568), .ZN(n498) );
  XNOR2_X1 U555 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n500), .B(n499), .ZN(G1351GAT) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U559 ( .A(n501), .B(KEYINPUT96), .ZN(n502) );
  XOR2_X1 U560 ( .A(KEYINPUT97), .B(n502), .Z(n508) );
  NOR2_X1 U561 ( .A1(n580), .A2(n547), .ZN(n503) );
  XNOR2_X1 U562 ( .A(n503), .B(KEYINPUT16), .ZN(n505) );
  NAND2_X1 U563 ( .A1(n505), .A2(n504), .ZN(n519) );
  NOR2_X1 U564 ( .A1(n506), .A2(n519), .ZN(n512) );
  NAND2_X1 U565 ( .A1(n512), .A2(n417), .ZN(n507) );
  XNOR2_X1 U566 ( .A(n508), .B(n507), .ZN(G1324GAT) );
  NAND2_X1 U567 ( .A1(n512), .A2(n535), .ZN(n509) );
  XNOR2_X1 U568 ( .A(n509), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U569 ( .A(G15GAT), .B(KEYINPUT35), .Z(n511) );
  NAND2_X1 U570 ( .A1(n512), .A2(n537), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(G1326GAT) );
  NAND2_X1 U572 ( .A1(n512), .A2(n527), .ZN(n513) );
  XNOR2_X1 U573 ( .A(n513), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U574 ( .A1(n517), .A2(n535), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n514), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U576 ( .A1(n517), .A2(n537), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n515), .B(KEYINPUT40), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G43GAT), .B(n516), .ZN(G1330GAT) );
  NAND2_X1 U579 ( .A1(n517), .A2(n527), .ZN(n518) );
  XNOR2_X1 U580 ( .A(n518), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n522) );
  NOR2_X1 U582 ( .A1(n520), .A2(n519), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n417), .A2(n528), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n522), .B(n521), .ZN(G1332GAT) );
  XOR2_X1 U585 ( .A(G64GAT), .B(KEYINPUT101), .Z(n524) );
  NAND2_X1 U586 ( .A1(n528), .A2(n535), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(G1333GAT) );
  NAND2_X1 U588 ( .A1(n537), .A2(n528), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(KEYINPUT102), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G71GAT), .B(n526), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT103), .B(KEYINPUT43), .Z(n530) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U594 ( .A(G78GAT), .B(n531), .Z(G1335GAT) );
  NAND2_X1 U595 ( .A1(n538), .A2(n417), .ZN(n534) );
  XOR2_X1 U596 ( .A(G85GAT), .B(KEYINPUT105), .Z(n532) );
  XNOR2_X1 U597 ( .A(KEYINPUT106), .B(n532), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1336GAT) );
  NAND2_X1 U599 ( .A1(n538), .A2(n535), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n539), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U603 ( .A1(n548), .A2(n540), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n541), .B(G113GAT), .ZN(G1340GAT) );
  INV_X1 U605 ( .A(n580), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n548), .A2(n542), .ZN(n544) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(n546) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n551), .A2(n570), .ZN(n559) );
  NOR2_X1 U615 ( .A1(n572), .A2(n559), .ZN(n552) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n557) );
  INV_X1 U620 ( .A(n555), .ZN(n564) );
  NOR2_X1 U621 ( .A1(n564), .A2(n559), .ZN(n556) );
  XOR2_X1 U622 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U623 ( .A1(n580), .A2(n559), .ZN(n558) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NOR2_X1 U627 ( .A1(n572), .A2(n568), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G169GAT), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT123), .ZN(G1348GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n568), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U634 ( .A1(n580), .A2(n568), .ZN(n569) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n582) );
  NOR2_X1 U637 ( .A1(n582), .A2(n572), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n582), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n582), .ZN(n581) );
  XOR2_X1 U646 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G218GAT), .B(n586), .Z(G1355GAT) );
endmodule

