//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT75), .Z(new_n189));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT80), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G137), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G119), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G128), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n198), .B2(new_n201), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n199), .B1(new_n203), .B2(new_n197), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G110), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT24), .B(G110), .ZN(new_n206));
  INV_X1    g020(.A(new_n203), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  OR3_X1    g023(.A1(new_n209), .A2(KEYINPUT16), .A3(G140), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT77), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(KEYINPUT76), .B2(G125), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n209), .A2(KEYINPUT77), .ZN(new_n213));
  OAI21_X1  g027(.A(G140), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT76), .A2(G125), .ZN(new_n215));
  AOI21_X1  g029(.A(G140), .B1(new_n215), .B2(KEYINPUT77), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n219));
  OAI211_X1 g033(.A(KEYINPUT78), .B(new_n210), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(KEYINPUT77), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(KEYINPUT77), .B2(new_n209), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n216), .B1(new_n223), .B2(G140), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT16), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n220), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n210), .A2(KEYINPUT78), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(new_n224), .B2(KEYINPUT16), .ZN(new_n229));
  AND4_X1   g043(.A1(new_n225), .A2(new_n214), .A3(KEYINPUT16), .A4(new_n217), .ZN(new_n230));
  OAI21_X1  g044(.A(G146), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n208), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G125), .B(G140), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n221), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT79), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n207), .A2(new_n206), .ZN(new_n236));
  INV_X1    g050(.A(G110), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n237), .B(new_n199), .C1(new_n203), .C2(new_n197), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n235), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n231), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n196), .B1(new_n232), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n227), .A2(new_n231), .ZN(new_n243));
  INV_X1    g057(.A(new_n208), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n240), .A3(new_n195), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n190), .B1(new_n247), .B2(G902), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n246), .ZN(new_n249));
  INV_X1    g063(.A(G902), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n189), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n188), .A2(new_n250), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G104), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G107), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G101), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n256), .A2(G107), .ZN(new_n263));
  OR2_X1    g077(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g078(.A(G107), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G104), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n261), .A2(new_n262), .A3(new_n263), .A4(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n265), .A2(G104), .ZN(new_n269));
  OAI21_X1  g083(.A(G101), .B1(new_n257), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT83), .B(G101), .C1(new_n257), .C2(new_n269), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n268), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT1), .A3(G146), .ZN(new_n276));
  XNOR2_X1  g090(.A(G143), .B(G146), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(G128), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT84), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n221), .A2(G143), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(G146), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT84), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n284), .B(new_n276), .C1(new_n277), .C2(G128), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n279), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n274), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n268), .A2(new_n272), .A3(new_n273), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n283), .B(new_n276), .C1(G128), .C2(new_n277), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G137), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT11), .A3(G134), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT11), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G137), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G131), .ZN(new_n298));
  INV_X1    g112(.A(G134), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT64), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT64), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G134), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n293), .A2(KEYINPUT11), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n297), .A2(new_n298), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n298), .B1(new_n297), .B2(new_n304), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT12), .B1(new_n292), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n281), .A2(new_n282), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT0), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(new_n201), .ZN(new_n311));
  NOR2_X1   g125(.A1(KEYINPUT0), .A2(G128), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n277), .B1(new_n310), .B2(new_n201), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n266), .B1(new_n264), .B2(new_n258), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n263), .B1(new_n257), .B2(new_n260), .ZN(new_n317));
  OAI21_X1  g131(.A(G101), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n315), .B1(new_n318), .B2(KEYINPUT4), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n268), .A2(KEYINPUT4), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(new_n318), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n318), .A2(new_n321), .A3(new_n268), .A4(KEYINPUT4), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n320), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT10), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n290), .A2(new_n327), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n287), .A2(new_n327), .B1(new_n274), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n307), .B(KEYINPUT85), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G110), .B(G140), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n191), .A2(G227), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n307), .B1(new_n287), .B2(new_n291), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT12), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n308), .A2(new_n331), .A3(new_n335), .A4(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT87), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n336), .B(KEYINPUT12), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n342), .A2(KEYINPUT87), .A3(new_n335), .A4(new_n331), .ZN(new_n343));
  INV_X1    g157(.A(new_n331), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n307), .B1(new_n326), .B2(new_n329), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n334), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n341), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G469), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n250), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT86), .ZN(new_n350));
  AND4_X1   g164(.A1(new_n334), .A2(new_n308), .A3(new_n331), .A4(new_n338), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n287), .A2(new_n327), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n328), .A2(new_n274), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n318), .A2(KEYINPUT4), .A3(new_n268), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT82), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n319), .B1(new_n356), .B2(new_n324), .ZN(new_n357));
  OAI22_X1  g171(.A1(new_n354), .A2(new_n357), .B1(new_n305), .B2(new_n306), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n334), .B1(new_n358), .B2(new_n331), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n350), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n335), .B1(new_n344), .B2(new_n345), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n308), .A2(new_n331), .A3(new_n334), .A4(new_n338), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(KEYINPUT86), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(G469), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n348), .A2(new_n250), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n349), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT9), .B(G234), .ZN(new_n368));
  OAI21_X1  g182(.A(G221), .B1(new_n368), .B2(G902), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G214), .B1(G237), .B2(G902), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G210), .B1(G237), .B2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n375));
  XNOR2_X1  g189(.A(G110), .B(G122), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n200), .A2(KEYINPUT66), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT66), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G119), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n380), .A3(G116), .ZN(new_n381));
  INV_X1    g195(.A(G116), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G119), .ZN(new_n383));
  INV_X1    g197(.A(G113), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT2), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT2), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G113), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n381), .A2(new_n383), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n381), .B2(new_n383), .ZN(new_n391));
  OAI22_X1  g205(.A1(new_n318), .A2(KEYINPUT4), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n356), .B2(new_n324), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n381), .A2(KEYINPUT5), .A3(new_n383), .ZN(new_n394));
  OAI21_X1  g208(.A(G113), .B1(new_n381), .B2(KEYINPUT5), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT88), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n381), .A2(KEYINPUT5), .A3(new_n383), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT88), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n198), .A2(new_n399), .A3(G116), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n397), .A2(new_n398), .A3(G113), .A4(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n274), .A2(new_n396), .A3(new_n389), .A4(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n375), .B(new_n377), .C1(new_n393), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT89), .ZN(new_n405));
  INV_X1    g219(.A(new_n392), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n323), .B2(new_n325), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n402), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT89), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n375), .A4(new_n377), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n315), .A2(G125), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n289), .A2(new_n209), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G224), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G953), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n414), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n377), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n407), .A2(new_n376), .A3(new_n402), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(KEYINPUT6), .A3(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n411), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n393), .A2(new_n403), .A3(new_n377), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT7), .B1(new_n415), .B2(G953), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n414), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n376), .B(KEYINPUT8), .Z(new_n429));
  OAI21_X1  g243(.A(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n429), .B1(new_n274), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n396), .A2(new_n389), .A3(new_n288), .A4(new_n401), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n414), .A2(KEYINPUT90), .A3(new_n425), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n412), .A2(new_n413), .A3(new_n424), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n428), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n250), .B1(new_n423), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT91), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(new_n250), .C1(new_n423), .C2(new_n436), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n374), .B1(new_n422), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n411), .A2(new_n418), .A3(new_n421), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n443), .A2(new_n373), .A3(new_n440), .A4(new_n438), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n372), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n370), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(G237), .A2(G953), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(G143), .A3(G214), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(G143), .B1(new_n447), .B2(G214), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT17), .A3(G131), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(G131), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT17), .ZN(new_n454));
  INV_X1    g268(.A(new_n450), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n298), .A3(new_n448), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n227), .A2(new_n231), .A3(new_n452), .A4(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G113), .B(G122), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT92), .B(G104), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n459), .B(new_n460), .Z(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(KEYINPUT18), .A2(G131), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n451), .B(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n224), .A2(new_n221), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n464), .B1(new_n235), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n458), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n462), .B1(new_n458), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n250), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G475), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT20), .ZN(new_n472));
  INV_X1    g286(.A(new_n231), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n453), .A2(new_n456), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT19), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n233), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n224), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n474), .B1(G146), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n466), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n461), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n467), .ZN(new_n481));
  NOR2_X1   g295(.A1(G475), .A2(G902), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n472), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n482), .ZN(new_n484));
  AOI211_X1 g298(.A(KEYINPUT20), .B(new_n484), .C1(new_n480), .C2(new_n467), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n471), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n382), .A2(KEYINPUT14), .A3(G122), .ZN(new_n488));
  XNOR2_X1  g302(.A(G116), .B(G122), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(G107), .B(new_n488), .C1(new_n490), .C2(KEYINPUT14), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n265), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n300), .A2(new_n302), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n275), .A2(G128), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n201), .A2(G143), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n491), .B(new_n492), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n489), .B(new_n265), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n495), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n494), .A2(new_n501), .ZN(new_n504));
  OAI21_X1  g318(.A(G134), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(new_n505), .A3(new_n496), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n368), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(G217), .A3(new_n191), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n507), .B(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n250), .ZN(new_n511));
  INV_X1    g325(.A(G478), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n511), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n487), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n191), .A2(G952), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(G234), .B2(G237), .ZN(new_n518));
  AOI211_X1 g332(.A(new_n250), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT21), .B(G898), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n446), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n447), .A2(G210), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT27), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(G101), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n315), .B1(new_n305), .B2(new_n306), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n297), .A2(new_n298), .A3(new_n304), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n298), .B1(G134), .B2(G137), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n300), .A2(new_n302), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(G137), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n289), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n381), .A2(new_n383), .ZN(new_n535));
  INV_X1    g349(.A(new_n388), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n537), .A2(KEYINPUT67), .A3(new_n389), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT67), .B1(new_n537), .B2(new_n389), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n529), .B(new_n534), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n390), .A2(new_n391), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n294), .A2(new_n296), .ZN(new_n544));
  OAI21_X1  g358(.A(G131), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n545), .A2(new_n530), .B1(new_n313), .B2(new_n314), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n289), .A2(new_n530), .A3(new_n533), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n548), .A3(KEYINPUT68), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT28), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n541), .B1(new_n529), .B2(new_n534), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT68), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT69), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n540), .A2(new_n550), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n554), .B1(new_n549), .B2(new_n553), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n528), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT30), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT65), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(KEYINPUT65), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n562), .B(new_n563), .C1(new_n546), .C2(new_n547), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n529), .A2(KEYINPUT65), .A3(new_n561), .A4(new_n534), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n542), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n528), .A3(new_n540), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT31), .ZN(new_n569));
  INV_X1    g383(.A(new_n540), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n566), .B2(new_n542), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT31), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n528), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT70), .B1(new_n560), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n572), .B1(new_n571), .B2(new_n528), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n541), .B1(new_n564), .B2(new_n565), .ZN(new_n578));
  INV_X1    g392(.A(new_n528), .ZN(new_n579));
  NOR4_X1   g393(.A1(new_n578), .A2(new_n570), .A3(KEYINPUT31), .A4(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n555), .A2(new_n556), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n579), .B1(new_n582), .B2(new_n558), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n576), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT71), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n575), .A2(KEYINPUT71), .A3(new_n576), .A4(new_n585), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT74), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n584), .B1(new_n581), .B2(new_n583), .ZN(new_n594));
  INV_X1    g408(.A(new_n576), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n559), .A2(new_n528), .A3(new_n556), .A4(new_n555), .ZN(new_n597));
  INV_X1    g411(.A(new_n571), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT29), .B1(new_n598), .B2(new_n579), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT72), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n538), .A2(new_n539), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n546), .B2(new_n547), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n550), .B1(new_n603), .B2(new_n540), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n556), .A2(KEYINPUT73), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n556), .A2(KEYINPUT73), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n528), .A2(KEYINPUT29), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT72), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n597), .A2(new_n612), .A3(new_n599), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n601), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n596), .A2(KEYINPUT32), .B1(new_n614), .B2(G472), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n591), .A2(new_n592), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n592), .B1(new_n591), .B2(new_n615), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n255), .B(new_n524), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  INV_X1    g433(.A(new_n370), .ZN(new_n620));
  INV_X1    g434(.A(new_n255), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n521), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n445), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(G478), .A2(G902), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n511), .B2(G478), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n510), .B(KEYINPUT33), .Z(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n627), .B2(G478), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n487), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n575), .A2(new_n250), .A3(new_n585), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n588), .A2(new_n634), .A3(new_n590), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n622), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  NAND2_X1  g452(.A1(new_n487), .A2(new_n514), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n624), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n622), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT93), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  INV_X1    g458(.A(new_n446), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT95), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n195), .A2(KEYINPUT36), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT94), .B1(new_n232), .B2(new_n241), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT94), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n245), .A2(new_n649), .A3(new_n240), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n647), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n648), .A2(new_n647), .A3(new_n650), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n253), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n646), .B1(new_n252), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n189), .ZN(new_n656));
  INV_X1    g470(.A(new_n251), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT25), .B1(new_n249), .B2(new_n250), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n654), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT95), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n645), .A2(new_n522), .A3(new_n635), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT37), .B(G110), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  XNOR2_X1  g481(.A(new_n518), .B(KEYINPUT99), .ZN(new_n668));
  OR2_X1    g482(.A1(KEYINPUT98), .A2(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(KEYINPUT98), .A2(G900), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n519), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n487), .A2(new_n514), .A3(new_n672), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n445), .A2(new_n370), .A3(new_n662), .A4(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n616), .B2(new_n617), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(KEYINPUT100), .B(new_n674), .C1(new_n616), .C2(new_n617), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XOR2_X1   g494(.A(new_n672), .B(KEYINPUT39), .Z(new_n681));
  NOR2_X1   g495(.A1(new_n620), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n596), .A2(KEYINPUT32), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n571), .A2(new_n579), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n603), .A2(new_n579), .A3(new_n540), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n250), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n591), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n442), .A2(new_n444), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n486), .A2(new_n514), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n694), .A2(new_n372), .A3(new_n662), .A4(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n684), .A2(new_n690), .A3(new_n691), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT102), .B(G143), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G45));
  AND3_X1   g513(.A1(new_n486), .A2(new_n628), .A3(new_n672), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n692), .A3(new_n701), .A4(new_n371), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n370), .A3(new_n662), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n701), .B1(new_n445), .B2(new_n700), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n616), .B2(new_n617), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  INV_X1    g522(.A(new_n349), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n348), .B1(new_n347), .B2(new_n250), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n369), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n255), .B(new_n713), .C1(new_n616), .C2(new_n617), .ZN(new_n714));
  INV_X1    g528(.A(new_n632), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n708), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n591), .A2(new_n615), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT74), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n591), .A2(new_n592), .A3(new_n615), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n621), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(KEYINPUT104), .A3(new_n632), .A4(new_n713), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n719), .ZN(new_n725));
  AND4_X1   g539(.A1(new_n725), .A2(new_n255), .A3(new_n640), .A4(new_n713), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n382), .ZN(G18));
  AND4_X1   g541(.A1(new_n445), .A2(new_n713), .A3(new_n522), .A4(new_n662), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  XNOR2_X1  g544(.A(new_n695), .B(KEYINPUT108), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n731), .A2(new_n624), .A3(new_n711), .A4(new_n712), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n574), .B1(new_n608), .B2(new_n579), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT105), .B1(new_n733), .B2(new_n595), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n581), .B1(new_n609), .B2(new_n528), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n576), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n738), .A2(new_n634), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n255), .A2(KEYINPUT106), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n252), .B2(new_n254), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n739), .A2(KEYINPUT107), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT107), .B1(new_n739), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n732), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NAND3_X1  g561(.A1(new_n662), .A2(new_n634), .A3(new_n738), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n445), .A3(new_n700), .A4(new_n713), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  NOR2_X1   g565(.A1(new_n692), .A2(new_n372), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n361), .A2(new_n362), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n365), .B1(new_n753), .B2(G469), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n712), .B1(new_n349), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n752), .A2(new_n700), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n743), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n685), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n589), .B1(new_n614), .B2(G472), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n685), .B(new_n760), .C1(new_n764), .C2(new_n596), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n763), .B1(new_n762), .B2(new_n765), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n758), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n752), .A2(new_n700), .A3(new_n755), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n255), .B(new_n769), .C1(new_n616), .C2(new_n617), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n757), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT109), .B1(new_n720), .B2(new_n769), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n768), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G131), .ZN(G33));
  AND3_X1   g589(.A1(new_n752), .A2(new_n673), .A3(new_n755), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n255), .B(new_n776), .C1(new_n616), .C2(new_n617), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NAND2_X1  g592(.A1(new_n487), .A2(new_n628), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT43), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n662), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(new_n635), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT45), .B1(new_n360), .B2(new_n363), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n753), .A2(KEYINPUT45), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n787), .A2(new_n788), .A3(new_n348), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(new_n365), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n709), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n791), .B2(new_n790), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n369), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n681), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n785), .A2(new_n752), .A3(new_n786), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  XNOR2_X1  g611(.A(new_n794), .B(KEYINPUT47), .ZN(new_n798));
  INV_X1    g612(.A(new_n725), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n621), .A3(new_n700), .A4(new_n752), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n798), .A2(KEYINPUT112), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT112), .B1(new_n798), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  OR2_X1    g618(.A1(new_n766), .A2(new_n767), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n780), .A2(new_n668), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n713), .A2(new_n752), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT48), .Z(new_n810));
  NAND2_X1  g624(.A1(new_n255), .A2(new_n518), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n807), .A2(new_n690), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n630), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n517), .B(KEYINPUT118), .Z(new_n814));
  NOR2_X1   g628(.A1(new_n744), .A2(new_n745), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n806), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n713), .ZN(new_n817));
  INV_X1    g631(.A(new_n445), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n813), .B(new_n814), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n694), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n372), .B1(KEYINPUT116), .B2(KEYINPUT50), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n824));
  OR3_X1    g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n798), .B1(new_n369), .B2(new_n711), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n752), .A3(new_n816), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n808), .A2(new_n749), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT117), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n487), .A2(new_n629), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n830), .B1(new_n812), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n825), .A2(new_n826), .A3(new_n828), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n810), .B(new_n819), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT100), .B1(new_n725), .B2(new_n674), .ZN(new_n838));
  INV_X1    g652(.A(new_n678), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n731), .A2(new_n818), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n659), .A2(new_n660), .A3(new_n672), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n690), .A2(new_n841), .A3(new_n755), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n706), .A2(new_n750), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT52), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n706), .A2(new_n750), .A3(new_n843), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n679), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n729), .A2(new_n746), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n726), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n618), .A2(new_n636), .A3(new_n641), .A4(new_n663), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n769), .A2(new_n853), .A3(new_n662), .A4(new_n739), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT113), .B1(new_n748), .B2(new_n756), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n516), .B1(new_n668), .B2(new_n671), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n370), .A2(new_n857), .A3(new_n662), .A4(new_n752), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n616), .B2(new_n617), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n777), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n774), .A2(new_n722), .A3(new_n851), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n849), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n862), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n679), .A2(new_n846), .A3(new_n847), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n847), .B1(new_n679), .B2(new_n846), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT114), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n845), .B2(new_n848), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n865), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n864), .B1(new_n871), .B2(new_n863), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n866), .A2(new_n867), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n865), .A2(new_n876), .A3(KEYINPUT53), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT114), .B1(new_n866), .B2(new_n867), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n845), .A2(new_n869), .A3(new_n848), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n862), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n877), .B(new_n874), .C1(new_n880), .C2(KEYINPUT53), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT115), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n863), .B1(new_n849), .B2(new_n862), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n871), .B2(new_n863), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n875), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n837), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n711), .B(KEYINPUT49), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n369), .A2(new_n371), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n888), .A2(new_n759), .A3(new_n779), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n694), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n690), .B2(new_n891), .ZN(G75));
  NAND2_X1  g706(.A1(new_n411), .A2(new_n421), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT119), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n417), .ZN(new_n896));
  INV_X1    g710(.A(G210), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n872), .A2(new_n897), .A3(new_n250), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n898), .B2(KEYINPUT56), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n191), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n872), .B2(new_n250), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n877), .B1(new_n880), .B2(KEYINPUT53), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(KEYINPUT120), .A3(G902), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n374), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n902), .B1(new_n907), .B2(new_n908), .ZN(G51));
  XNOR2_X1  g723(.A(new_n365), .B(KEYINPUT57), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n872), .A2(new_n874), .ZN(new_n911));
  INV_X1    g725(.A(new_n881), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n347), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n904), .A2(new_n789), .A3(new_n906), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n900), .B1(new_n914), .B2(new_n915), .ZN(G54));
  AND2_X1   g730(.A1(KEYINPUT58), .A2(G475), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n904), .A2(new_n906), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n919));
  INV_X1    g733(.A(new_n481), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n904), .A2(new_n481), .A3(new_n906), .A4(new_n917), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n901), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(G60));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n627), .B(KEYINPUT122), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n625), .B(KEYINPUT59), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n881), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n926), .B1(new_n932), .B2(new_n901), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n927), .B1(new_n886), .B2(new_n928), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n931), .A2(KEYINPUT123), .A3(new_n900), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G63));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n871), .A2(new_n863), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(new_n877), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n937), .B(new_n901), .C1(new_n941), .C2(new_n249), .ZN(new_n942));
  INV_X1    g756(.A(new_n939), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n249), .B1(new_n905), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT124), .B1(new_n944), .B2(new_n900), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n652), .A2(new_n653), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n905), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n942), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n901), .B1(new_n941), .B2(new_n249), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n944), .A2(new_n900), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(KEYINPUT125), .A3(KEYINPUT61), .A4(new_n947), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n950), .A2(new_n957), .ZN(G66));
  OAI21_X1  g772(.A(G953), .B1(new_n520), .B2(new_n415), .ZN(new_n959));
  INV_X1    g773(.A(new_n852), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n851), .A2(new_n722), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n959), .B1(new_n962), .B2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n894), .B1(G898), .B2(new_n191), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT127), .Z(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(G69));
  XNOR2_X1  g780(.A(new_n566), .B(new_n477), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(G900), .B2(G953), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n805), .A2(new_n795), .A3(new_n841), .ZN(new_n969));
  AND4_X1   g783(.A1(new_n777), .A2(new_n803), .A3(new_n796), .A4(new_n969), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n679), .A2(new_n706), .A3(new_n750), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n774), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n972), .B2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n631), .A2(new_n639), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n720), .A2(new_n682), .A3(new_n752), .A4(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n803), .A2(new_n796), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n971), .A2(new_n697), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n976), .B1(KEYINPUT62), .B2(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n967), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n973), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n973), .B(new_n985), .C1(new_n980), .C2(new_n981), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(G72));
  INV_X1    g801(.A(new_n686), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n978), .A2(new_n962), .A3(new_n979), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n571), .A2(new_n579), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n970), .A2(new_n774), .A3(new_n962), .A4(new_n971), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(new_n991), .ZN(new_n995));
  AND4_X1   g809(.A1(new_n988), .A2(new_n884), .A3(new_n991), .A4(new_n993), .ZN(new_n996));
  NOR4_X1   g810(.A1(new_n992), .A2(new_n995), .A3(new_n996), .A4(new_n900), .ZN(G57));
endmodule


