//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n907, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202));
  AND2_X1   g001(.A1(G15gat), .A2(G22gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G15gat), .A2(G22gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT96), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G15gat), .ZN(new_n206));
  INV_X1    g005(.A(G22gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT96), .ZN(new_n209));
  NAND2_X1  g008(.A1(G15gat), .A2(G22gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G1gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT16), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n205), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(G1gat), .B1(new_n205), .B2(new_n211), .ZN(new_n215));
  OAI21_X1  g014(.A(G8gat), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT96), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n209), .B1(new_n208), .B2(new_n210), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n212), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n205), .A2(new_n211), .A3(new_n213), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT91), .ZN(new_n224));
  INV_X1    g023(.A(G29gat), .ZN(new_n225));
  INV_X1    g024(.A(G36gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT91), .A2(G29gat), .A3(G36gat), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT14), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT14), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(G29gat), .B2(G36gat), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT95), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT95), .B1(new_n230), .B2(new_n232), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n229), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G43gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(G50gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT94), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(G50gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(KEYINPUT94), .A3(G50gat), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT15), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G50gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G43gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n239), .A2(new_n244), .A3(KEYINPUT15), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT93), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n239), .A2(new_n244), .A3(KEYINPUT93), .A4(KEYINPUT15), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n235), .A2(new_n242), .A3(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n227), .A2(new_n230), .A3(new_n232), .A4(new_n228), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT92), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n239), .A2(new_n244), .A3(KEYINPUT15), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT17), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n247), .A2(new_n248), .ZN(new_n258));
  INV_X1    g057(.A(new_n234), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT95), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n239), .A2(new_n238), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(new_n244), .A3(new_n241), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT15), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n258), .A2(new_n261), .A3(new_n229), .A4(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT17), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n253), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT92), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n253), .A3(new_n252), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n223), .B1(new_n257), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT97), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n223), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n216), .A2(new_n222), .A3(KEYINPUT97), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n275), .A2(new_n276), .B1(new_n271), .B2(new_n266), .ZN(new_n277));
  NAND2_X1  g076(.A1(G229gat), .A2(G233gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n273), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n202), .B1(new_n280), .B2(KEYINPUT18), .ZN(new_n281));
  INV_X1    g080(.A(new_n223), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n250), .A2(new_n256), .A3(KEYINPUT17), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n267), .B1(new_n266), .B2(new_n271), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n271), .ZN(new_n286));
  INV_X1    g085(.A(new_n276), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT97), .B1(new_n216), .B2(new_n222), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n285), .A2(new_n289), .A3(KEYINPUT18), .A4(new_n278), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(new_n278), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n287), .A2(new_n286), .A3(new_n288), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(new_n277), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G113gat), .B(G141gat), .ZN(new_n297));
  INV_X1    g096(.A(G197gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT11), .B(G169gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n289), .A3(new_n278), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT18), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(KEYINPUT99), .A3(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n281), .A2(new_n296), .A3(new_n302), .A4(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n302), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n280), .A2(KEYINPUT18), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n295), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n306), .A2(KEYINPUT100), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT100), .B1(new_n306), .B2(new_n310), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT25), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT24), .ZN(new_n319));
  NOR2_X1   g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  OAI211_X1 g119(.A(KEYINPUT65), .B(new_n317), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(G169gat), .B2(G176gat), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n323), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n322), .B(new_n325), .C1(G169gat), .C2(G176gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n320), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(KEYINPUT24), .A3(new_n318), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT65), .B1(new_n329), .B2(new_n317), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n315), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n323), .A2(KEYINPUT23), .ZN(new_n332));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT67), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT67), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n338), .B(new_n317), .C1(new_n319), .C2(new_n320), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT25), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n331), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n344), .A2(KEYINPUT68), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(KEYINPUT68), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n344), .A2(KEYINPUT68), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OR3_X1    g151(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n333), .A3(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n347), .A2(new_n352), .A3(new_n318), .A4(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n341), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358));
  OR3_X1    g157(.A1(new_n357), .A2(KEYINPUT29), .A3(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(KEYINPUT75), .B(KEYINPUT22), .Z(new_n360));
  INV_X1    g159(.A(G211gat), .ZN(new_n361));
  INV_X1    g160(.A(G218gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(new_n366), .A3(new_n364), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n356), .B(KEYINPUT69), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n341), .A3(new_n358), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n359), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n341), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n358), .A2(KEYINPUT29), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n374), .A2(new_n375), .B1(new_n357), .B2(new_n358), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT30), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT30), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n373), .B(new_n379), .C1(new_n370), .C2(new_n376), .ZN(new_n380));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n378), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n377), .A2(KEYINPUT30), .A3(new_n383), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT78), .Z(new_n389));
  XOR2_X1   g188(.A(G127gat), .B(G134gat), .Z(new_n390));
  XNOR2_X1  g189(.A(G113gat), .B(G120gat), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n390), .B(KEYINPUT70), .C1(KEYINPUT1), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT70), .ZN(new_n393));
  INV_X1    g192(.A(G120gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G113gat), .ZN(new_n395));
  INV_X1    g194(.A(G113gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G120gat), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT1), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G127gat), .B(G134gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n392), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n399), .A2(KEYINPUT72), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT71), .B(G113gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n395), .B1(new_n403), .B2(new_n394), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT1), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(KEYINPUT72), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n402), .A2(new_n404), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT77), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n401), .A2(new_n407), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT77), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413));
  INV_X1    g212(.A(G155gat), .ZN(new_n414));
  INV_X1    g213(.A(G162gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT2), .ZN(new_n419));
  INV_X1    g218(.A(G148gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G141gat), .ZN(new_n421));
  INV_X1    g220(.A(G141gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G148gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n418), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n421), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n421), .B2(new_n423), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n417), .B1(new_n416), .B2(KEYINPUT2), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n410), .A2(new_n412), .B1(new_n413), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT3), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n389), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT4), .B1(new_n411), .B2(new_n433), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n431), .A2(new_n438), .A3(new_n401), .A4(new_n407), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n435), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n389), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n433), .A2(new_n411), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n410), .A2(new_n412), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(new_n433), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n441), .B(KEYINPUT5), .C1(new_n442), .C2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G1gat), .B(G29gat), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n449), .B(new_n450), .Z(new_n451));
  INV_X1    g250(.A(KEYINPUT81), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT80), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n439), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n453), .A3(new_n452), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n436), .A3(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n439), .A2(new_n453), .A3(new_n452), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n437), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT5), .ZN(new_n461));
  AND4_X1   g260(.A1(KEYINPUT82), .A2(new_n460), .A3(new_n461), .A4(new_n435), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT5), .B1(new_n457), .B2(new_n459), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT82), .B1(new_n463), .B2(new_n435), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n446), .B(new_n451), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n435), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n463), .A2(KEYINPUT82), .A3(new_n435), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n451), .B1(new_n473), .B2(new_n446), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  AOI221_X4 g274(.A(new_n451), .B1(new_n466), .B2(new_n467), .C1(new_n473), .C2(new_n446), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n387), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT84), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n479), .B(new_n387), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT69), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n356), .B(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n336), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n335), .A2(new_n484), .A3(new_n321), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n334), .B1(KEYINPUT67), .B2(new_n336), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n339), .A2(KEYINPUT25), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n485), .A2(new_n315), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n411), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n356), .A2(KEYINPUT69), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n356), .A2(KEYINPUT69), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n341), .B(new_n408), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G227gat), .A2(G233gat), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n494), .B(KEYINPUT64), .Z(new_n495));
  NOR2_X1   g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n492), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n408), .B1(new_n371), .B2(new_n341), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT33), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(KEYINPUT32), .B2(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(G15gat), .B(G43gat), .Z(new_n503));
  XNOR2_X1  g302(.A(G71gat), .B(G99gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT32), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(new_n493), .B2(new_n495), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(KEYINPUT33), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n495), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(new_n489), .B2(new_n492), .ZN(new_n513));
  INV_X1    g312(.A(new_n510), .ZN(new_n514));
  NOR4_X1   g313(.A1(new_n513), .A2(KEYINPUT73), .A3(new_n508), .A4(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n506), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT34), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n512), .B2(KEYINPUT74), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n500), .A2(KEYINPUT32), .A3(new_n510), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT73), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n509), .A2(new_n507), .A3(new_n510), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n520), .B1(new_n524), .B2(new_n506), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n497), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n370), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n431), .A2(new_n413), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n528), .A2(KEYINPUT86), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT86), .B1(new_n528), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT29), .B1(new_n368), .B2(new_n369), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n433), .B1(new_n533), .B2(KEYINPUT3), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT85), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G228gat), .A2(G233gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(KEYINPUT85), .B(new_n433), .C1(new_n533), .C2(KEYINPUT3), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n532), .A2(new_n536), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n534), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n370), .B1(new_n529), .B2(new_n528), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n207), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n207), .A3(new_n543), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G78gat), .B(G106gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT31), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(new_n243), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n545), .A2(new_n551), .A3(new_n546), .A4(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n516), .A2(new_n518), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n524), .A2(new_n520), .A3(new_n506), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n496), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n526), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n387), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n446), .B1(new_n462), .B2(new_n464), .ZN(new_n561));
  INV_X1    g360(.A(new_n451), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n467), .A3(new_n465), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(KEYINPUT6), .A3(new_n562), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT35), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n559), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n556), .A2(new_n496), .A3(new_n557), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n496), .B1(new_n556), .B2(new_n557), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n526), .A2(KEYINPUT36), .A3(new_n558), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n555), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n478), .B(new_n480), .C1(new_n568), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n445), .A2(new_n442), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT39), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n577), .B1(new_n576), .B2(KEYINPUT39), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n457), .A2(new_n459), .B1(new_n434), .B2(new_n432), .ZN(new_n580));
  OAI22_X1  g379(.A1(new_n578), .A2(new_n579), .B1(new_n442), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n442), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT88), .B(KEYINPUT39), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n451), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT40), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n474), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(new_n560), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT38), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT37), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n377), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n373), .B(KEYINPUT37), .C1(new_n370), .C2(new_n376), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI22_X1  g393(.A1(new_n594), .A2(new_n384), .B1(KEYINPUT38), .B2(new_n377), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n376), .A2(new_n527), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT90), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n359), .A2(new_n527), .A3(new_n372), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT37), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n599), .A2(new_n590), .A3(new_n383), .A4(new_n592), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n564), .A2(new_n595), .A3(new_n600), .A4(new_n565), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n589), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n555), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n572), .B2(new_n573), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n526), .A2(new_n555), .A3(new_n558), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n566), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n602), .A2(new_n604), .B1(new_n606), .B2(new_n567), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n314), .B1(new_n575), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT105), .Z(new_n610));
  NOR2_X1   g409(.A1(KEYINPUT102), .A2(G64gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(KEYINPUT102), .A2(G64gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(G57gat), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(G57gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n613), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(G71gat), .A2(G78gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT9), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n614), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n618), .B(KEYINPUT101), .ZN(new_n622));
  OR2_X1    g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n618), .B1(new_n623), .B2(new_n619), .ZN(new_n625));
  INV_X1    g424(.A(G64gat), .ZN(new_n626));
  OR3_X1    g425(.A1(new_n615), .A2(new_n626), .A3(KEYINPUT103), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n615), .B2(KEYINPUT103), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT21), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n632), .A2(new_n275), .A3(new_n276), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n633), .A2(G183gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(G183gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n634), .B2(new_n635), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n610), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  INV_X1    g440(.A(new_n610), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT104), .B(KEYINPUT21), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n630), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G127gat), .B(G155gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G211gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n645), .B(new_n647), .Z(new_n648));
  AND3_X1   g447(.A1(new_n640), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n640), .B2(new_n643), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(KEYINPUT106), .A2(G85gat), .A3(G92gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT7), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT7), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n654), .A2(KEYINPUT106), .A3(G85gat), .A4(G92gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(G99gat), .A2(G106gat), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n653), .A2(new_n655), .B1(KEYINPUT8), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G85gat), .ZN(new_n658));
  INV_X1    g457(.A(G92gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G99gat), .B(G106gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT108), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n653), .A2(new_n655), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n656), .A2(KEYINPUT8), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n666), .A2(new_n662), .A3(new_n660), .A4(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n657), .A2(KEYINPUT107), .A3(new_n662), .A4(new_n660), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n661), .A2(new_n673), .A3(new_n663), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n665), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n283), .B2(new_n284), .ZN(new_n676));
  NAND3_X1  g475(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n665), .A2(new_n674), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n286), .A3(new_n672), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G190gat), .B(G218gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(G134gat), .B(G162gat), .Z(new_n683));
  AOI21_X1  g482(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n681), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n676), .A2(new_n686), .A3(new_n677), .A4(new_n679), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n682), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n685), .B1(new_n682), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691));
  XNOR2_X1  g490(.A(G120gat), .B(G148gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(G176gat), .B(G204gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n630), .B1(new_n670), .B2(new_n671), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n696), .A2(new_n664), .B1(new_n675), .B2(new_n630), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT10), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n631), .A2(KEYINPUT10), .A3(new_n672), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n697), .A2(new_n698), .B1(new_n699), .B2(new_n678), .ZN(new_n700));
  NAND2_X1  g499(.A1(G230gat), .A2(G233gat), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT109), .Z(new_n702));
  OAI21_X1  g501(.A(new_n695), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704));
  INV_X1    g503(.A(new_n702), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n697), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n675), .A2(new_n630), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n631), .A2(new_n672), .A3(new_n664), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(KEYINPUT110), .A3(new_n702), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n691), .B1(new_n703), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n698), .A3(new_n708), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n678), .A3(KEYINPUT10), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n702), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n694), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n716), .A2(KEYINPUT111), .A3(new_n710), .A4(new_n706), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n697), .A2(new_n705), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n694), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n651), .A2(new_n690), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n608), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n475), .ZN(new_n724));
  INV_X1    g523(.A(new_n476), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n212), .ZN(G1324gat));
  NOR2_X1   g527(.A1(new_n723), .A2(new_n387), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n220), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT113), .Z(new_n731));
  INV_X1    g530(.A(KEYINPUT16), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n729), .B1(new_n732), .B2(new_n220), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n733), .A2(new_n734), .B1(KEYINPUT112), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(KEYINPUT42), .ZN(new_n738));
  OAI211_X1 g537(.A(KEYINPUT112), .B(new_n735), .C1(new_n733), .C2(new_n734), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n731), .A2(new_n738), .A3(new_n739), .ZN(G1325gat));
  INV_X1    g539(.A(new_n572), .ZN(new_n741));
  INV_X1    g540(.A(new_n573), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n723), .A2(new_n206), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n570), .A2(new_n571), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n608), .A2(new_n746), .A3(new_n722), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n206), .B2(new_n747), .ZN(G1326gat));
  NOR2_X1   g547(.A1(new_n723), .A2(new_n555), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT43), .B(G22gat), .Z(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1327gat));
  INV_X1    g550(.A(new_n651), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n721), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n306), .A2(new_n310), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n690), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(KEYINPUT44), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n575), .A2(new_n607), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n758), .B1(new_n575), .B2(new_n607), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n756), .B1(new_n575), .B2(new_n607), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n755), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G29gat), .B1(new_n767), .B2(new_n726), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n608), .A2(new_n690), .A3(new_n753), .ZN(new_n769));
  INV_X1    g568(.A(new_n726), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n225), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT45), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n772), .ZN(G1328gat));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n226), .A3(new_n560), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT46), .Z(new_n775));
  OAI21_X1  g574(.A(G36gat), .B1(new_n767), .B2(new_n387), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1329gat));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n769), .A2(KEYINPUT116), .A3(new_n236), .A4(new_n746), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n608), .A2(new_n746), .A3(new_n690), .A4(new_n753), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(G43gat), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n755), .ZN(new_n786));
  INV_X1    g585(.A(new_n757), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n575), .A2(new_n607), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n789), .B2(new_n759), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n763), .A2(new_n764), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n743), .B(new_n786), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G43gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n780), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n783), .A2(G43gat), .ZN(new_n796));
  AOI211_X1 g595(.A(new_n795), .B(new_n796), .C1(new_n792), .C2(G43gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n778), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n236), .B1(new_n766), .B2(new_n743), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n779), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n796), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n793), .A2(KEYINPUT47), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(KEYINPUT117), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n804), .ZN(G1330gat));
  INV_X1    g604(.A(new_n769), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n243), .B1(new_n806), .B2(new_n555), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n603), .A2(G50gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n767), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g609(.A1(new_n789), .A2(new_n759), .ZN(new_n811));
  INV_X1    g610(.A(new_n754), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n718), .A2(new_n720), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n651), .A2(new_n690), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n726), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(new_n615), .ZN(G1332gat));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n387), .ZN(new_n818));
  NOR2_X1   g617(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n819));
  AND2_X1   g618(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n818), .B2(new_n819), .ZN(G1333gat));
  INV_X1    g621(.A(new_n815), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(G71gat), .A3(new_n743), .ZN(new_n824));
  INV_X1    g623(.A(new_n746), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n815), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(G71gat), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g627(.A1(new_n823), .A2(new_n603), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g629(.A1(new_n651), .A2(new_n812), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT118), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n721), .B(new_n833), .C1(new_n790), .C2(new_n791), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n834), .A2(new_n658), .A3(new_n726), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n763), .A2(new_n833), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT51), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n763), .A2(new_n838), .A3(new_n833), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n721), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n770), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n835), .B1(new_n842), .B2(new_n658), .ZN(G1336gat));
  AND4_X1   g642(.A1(new_n659), .A2(new_n840), .A3(new_n560), .A4(new_n721), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846));
  OAI21_X1  g645(.A(G92gat), .B1(new_n834), .B2(new_n387), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n847), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT52), .B1(new_n849), .B2(new_n844), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1337gat));
  INV_X1    g650(.A(G99gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n841), .A2(new_n852), .A3(new_n746), .ZN(new_n853));
  OAI21_X1  g652(.A(G99gat), .B1(new_n834), .B2(new_n744), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1338gat));
  NAND4_X1  g654(.A1(new_n837), .A2(new_n603), .A3(new_n721), .A4(new_n839), .ZN(new_n856));
  INV_X1    g655(.A(G106gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n603), .A2(G106gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n834), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(G1339gat));
  NAND2_X1  g661(.A1(new_n713), .A2(new_n714), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n705), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n713), .A2(new_n702), .A3(new_n714), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n695), .B1(new_n715), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(KEYINPUT55), .A3(new_n868), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n718), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n279), .B1(new_n273), .B2(new_n277), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n275), .A2(new_n276), .A3(new_n271), .A4(new_n266), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n289), .A2(new_n876), .A3(new_n292), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n878), .B2(new_n301), .ZN(new_n879));
  INV_X1    g678(.A(new_n301), .ZN(new_n880));
  AOI211_X1 g679(.A(KEYINPUT119), .B(new_n880), .C1(new_n875), .C2(new_n877), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n690), .A2(new_n882), .A3(new_n306), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n873), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n718), .A2(new_n871), .A3(new_n872), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n690), .A2(new_n882), .A3(new_n306), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT120), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n721), .A2(new_n306), .A3(new_n882), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n754), .A2(new_n718), .A3(new_n871), .A4(new_n872), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n690), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n651), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n722), .A2(new_n812), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n896), .A2(new_n605), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n726), .A2(new_n560), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G113gat), .B1(new_n901), .B2(new_n314), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n812), .A2(new_n403), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(G1340gat));
  NOR2_X1   g703(.A1(new_n901), .A2(new_n813), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(new_n394), .ZN(G1341gat));
  NOR2_X1   g705(.A1(new_n901), .A2(new_n651), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n907), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g707(.A1(new_n901), .A2(new_n756), .ZN(new_n909));
  NOR2_X1   g708(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n910));
  AND2_X1   g709(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n912), .B1(new_n909), .B2(new_n910), .ZN(G1343gat));
  NAND2_X1  g712(.A1(new_n744), .A2(new_n900), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n915), .A2(new_n603), .A3(new_n898), .A4(new_n896), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(G141gat), .A3(new_n314), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(KEYINPUT58), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n885), .A2(new_n888), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n886), .A2(new_n311), .A3(new_n312), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n721), .A2(new_n306), .A3(new_n882), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n756), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n752), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n894), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n603), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n914), .B1(new_n925), .B2(KEYINPUT57), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n896), .A2(new_n927), .A3(new_n603), .A4(new_n898), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G141gat), .B1(new_n929), .B2(new_n314), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n918), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n926), .A2(new_n928), .A3(new_n754), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT122), .A3(G141gat), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT122), .B1(new_n932), .B2(G141gat), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n933), .A2(new_n934), .A3(new_n917), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(KEYINPUT123), .B(new_n931), .C1(new_n935), .C2(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1344gat));
  NOR3_X1   g740(.A1(new_n916), .A2(G148gat), .A3(new_n813), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT124), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n896), .A2(new_n603), .A3(new_n898), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT57), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n873), .A2(new_n883), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n752), .B1(new_n922), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n722), .A2(new_n314), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n927), .B(new_n603), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n946), .A2(new_n721), .A3(new_n915), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n944), .B1(new_n951), .B2(G148gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n944), .B1(new_n929), .B2(new_n813), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(new_n420), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n943), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT125), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n943), .B(new_n957), .C1(new_n952), .C2(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1345gat));
  NOR3_X1   g758(.A1(new_n929), .A2(new_n414), .A3(new_n651), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n916), .A2(new_n651), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n414), .B2(new_n961), .ZN(G1346gat));
  OAI21_X1  g761(.A(new_n415), .B1(new_n916), .B2(new_n756), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n690), .A2(G162gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n929), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT126), .ZN(G1347gat));
  NOR2_X1   g765(.A1(new_n770), .A2(new_n387), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n899), .A2(new_n967), .ZN(new_n968));
  OR3_X1    g767(.A1(new_n968), .A2(G169gat), .A3(new_n812), .ZN(new_n969));
  OAI21_X1  g768(.A(G169gat), .B1(new_n968), .B2(new_n314), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1348gat));
  NOR2_X1   g770(.A1(new_n968), .A2(new_n813), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(G176gat), .Z(G1349gat));
  NOR2_X1   g772(.A1(new_n968), .A2(new_n651), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n342), .ZN(new_n975));
  INV_X1    g774(.A(G183gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n974), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT60), .ZN(G1350gat));
  XNOR2_X1  g777(.A(KEYINPUT61), .B(G190gat), .ZN(new_n979));
  NAND2_X1  g778(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n968), .A2(new_n756), .ZN(new_n981));
  MUX2_X1   g780(.A(new_n979), .B(new_n980), .S(new_n981), .Z(G1351gat));
  INV_X1    g781(.A(new_n967), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n945), .A2(new_n743), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n984), .A2(new_n298), .A3(new_n754), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT127), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n946), .A2(new_n950), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n987), .A2(new_n743), .A3(new_n983), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n298), .B1(new_n988), .B2(new_n313), .ZN(new_n989));
  OR2_X1    g788(.A1(new_n986), .A2(new_n989), .ZN(G1352gat));
  INV_X1    g789(.A(G204gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n984), .A2(new_n991), .A3(new_n721), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n994));
  NOR4_X1   g793(.A1(new_n987), .A2(new_n743), .A3(new_n813), .A4(new_n983), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n993), .B(new_n994), .C1(new_n991), .C2(new_n995), .ZN(G1353gat));
  NAND3_X1  g795(.A1(new_n984), .A2(new_n361), .A3(new_n752), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n988), .A2(new_n752), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n998), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n999));
  AOI21_X1  g798(.A(KEYINPUT63), .B1(new_n998), .B2(G211gat), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(G1354gat));
  NAND3_X1  g800(.A1(new_n984), .A2(new_n362), .A3(new_n690), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n988), .A2(new_n690), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1002), .B1(new_n1003), .B2(new_n362), .ZN(G1355gat));
endmodule


