//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1176, new_n1177, new_n1178, new_n1179;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n449), .B1(new_n457), .B2(new_n454), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n463), .B(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(G137), .A2(new_n462), .B1(new_n465), .B2(G101), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n460), .A2(KEYINPUT68), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n475), .A2(new_n478), .A3(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n467), .B1(new_n477), .B2(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n460), .A2(new_n461), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n460), .A2(G2105), .ZN(new_n486));
  OAI221_X1 g061(.A(new_n482), .B1(new_n483), .B2(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(KEYINPUT4), .B(G138), .C1(new_n468), .C2(new_n469), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n460), .B2(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n494), .B2(new_n461), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n460), .A2(G138), .A3(new_n461), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(G164));
  NAND2_X1  g072(.A1(G75), .A2(G651), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT71), .B(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n499), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(new_n499), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n504), .A2(G543), .B1(G62), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n502), .B2(new_n507), .ZN(new_n511));
  XOR2_X1   g086(.A(KEYINPUT71), .B(KEYINPUT6), .Z(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(new_n507), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n513), .A2(new_n514), .A3(new_n500), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n509), .B1(new_n510), .B2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  AND3_X1   g094(.A1(new_n511), .A2(new_n516), .A3(G89), .ZN(new_n520));
  INV_X1    g095(.A(new_n500), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n521), .B1(new_n512), .B2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(G51), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n508), .A2(G63), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT73), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n523), .B(new_n524), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n520), .A2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n507), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(G651), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n511), .A2(new_n516), .A3(G90), .ZN(new_n539));
  OAI211_X1 g114(.A(G543), .B(new_n500), .C1(new_n501), .C2(new_n499), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n539), .A2(KEYINPUT75), .A3(new_n542), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(G171));
  NAND3_X1  g122(.A1(new_n511), .A2(new_n516), .A3(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n507), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n541), .A2(G43), .B1(new_n551), .B2(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT77), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n522), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n540), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n511), .A2(new_n516), .A3(G91), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n499), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n499), .B1(new_n507), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n541), .B2(G49), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n517), .B2(new_n575), .ZN(G288));
  INV_X1    g151(.A(G48), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n540), .A2(KEYINPUT79), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT79), .B1(new_n540), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n507), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n578), .A2(new_n579), .B1(G651), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n511), .A2(new_n516), .A3(G86), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n511), .A2(new_n516), .A3(KEYINPUT78), .A4(G86), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(G305));
  NAND3_X1  g163(.A1(new_n511), .A2(new_n516), .A3(G85), .ZN(new_n589));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n507), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n541), .A2(G47), .B1(new_n592), .B2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n517), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n511), .A2(new_n516), .A3(KEYINPUT10), .A4(G92), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT81), .B(G66), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n515), .A2(new_n602), .B1(G79), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n499), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(G54), .B2(new_n541), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n595), .A2(KEYINPUT80), .B1(new_n596), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(KEYINPUT80), .B2(new_n595), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT82), .ZN(G284));
  XNOR2_X1  g184(.A(new_n608), .B(KEYINPUT83), .ZN(G321));
  NAND2_X1  g185(.A1(G299), .A2(new_n596), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G168), .B2(new_n596), .ZN(G280));
  XOR2_X1   g187(.A(G280), .B(KEYINPUT84), .Z(G297));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT85), .B(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(G860), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT86), .Z(G148));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n465), .A2(new_n460), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT13), .Z(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  INV_X1    g202(.A(new_n486), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G123), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n462), .A2(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G2096), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n626), .A2(new_n627), .A3(new_n635), .ZN(G156));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT14), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n642), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n651), .A3(G14), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT87), .Z(G401));
  XNOR2_X1  g228(.A(G2072), .B(G2078), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT17), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  OR3_X1    g234(.A1(new_n656), .A2(new_n654), .A3(new_n657), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n656), .A2(new_n654), .A3(new_n657), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n634), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT89), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(new_n673), .ZN(new_n678));
  MUX2_X1   g253(.A(new_n678), .B(new_n677), .S(new_n670), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1986), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n686), .B1(new_n683), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(G229));
  XNOR2_X1  g265(.A(KEYINPUT27), .B(G1996), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT102), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI22_X1  g268(.A1(G129), .A2(new_n628), .B1(new_n465), .B2(G105), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT26), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n462), .A2(G141), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT100), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G29), .B2(G32), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT101), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n704), .A2(new_n705), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n693), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n708), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n710), .A2(new_n706), .A3(new_n692), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G34), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(G29), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G160), .B2(G29), .ZN(new_n715));
  INV_X1    g290(.A(G2084), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n709), .A2(new_n711), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G5), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G171), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(G1961), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n701), .A2(G26), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n628), .A2(G128), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n462), .A2(G140), .ZN(new_n726));
  NOR2_X1   g301(.A1(G104), .A2(G2105), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n725), .B(new_n726), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n724), .B1(new_n729), .B2(G29), .ZN(new_n730));
  INV_X1    g305(.A(G2067), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n701), .A2(G35), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G162), .B2(new_n701), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT29), .B(G2090), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2078), .ZN(new_n737));
  NAND2_X1  g312(.A1(G164), .A2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G27), .B2(G29), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n732), .B(new_n736), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n701), .A2(G33), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  INV_X1    g318(.A(G139), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n483), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n745), .A2(KEYINPUT98), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(KEYINPUT98), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  OAI22_X1  g323(.A1(new_n746), .A2(new_n747), .B1(new_n461), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n741), .B1(new_n749), .B2(G29), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2072), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n740), .B(new_n751), .C1(new_n737), .C2(new_n739), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n719), .A2(G20), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT23), .Z(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G299), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1956), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n718), .A2(new_n722), .A3(new_n752), .A4(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n719), .A2(G21), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G286), .B2(G16), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT103), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n760), .A2(new_n761), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT31), .B(G11), .Z(new_n765));
  INV_X1    g340(.A(G28), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(KEYINPUT30), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT104), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n766), .B2(KEYINPUT30), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n764), .B(new_n770), .C1(new_n701), .C2(new_n633), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n763), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  INV_X1    g348(.A(new_n721), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT105), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n719), .A2(G19), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n554), .B2(new_n719), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT97), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT96), .B(G1341), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n719), .A2(G4), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n614), .B2(new_n719), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT95), .B(G1348), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n775), .A2(new_n776), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n758), .A2(new_n777), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n719), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n719), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  INV_X1    g367(.A(G1971), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G6), .B(G305), .S(G16), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT32), .B(G1981), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n719), .A2(G23), .ZN(new_n798));
  INV_X1    g373(.A(G288), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n719), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT92), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT33), .B(G1976), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n794), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n462), .A2(G131), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT90), .ZN(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n809));
  INV_X1    g384(.A(G95), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n461), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT91), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n628), .A2(G119), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n808), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G25), .B(new_n814), .S(G29), .Z(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G290), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G16), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G16), .B2(G24), .ZN(new_n821));
  INV_X1    g396(.A(G1986), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n818), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n805), .A2(new_n806), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n805), .A2(new_n827), .A3(new_n806), .A4(new_n825), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n789), .B1(new_n829), .B2(new_n830), .ZN(G311));
  INV_X1    g406(.A(KEYINPUT106), .ZN(new_n832));
  NOR2_X1   g407(.A1(G311), .A2(new_n832), .ZN(new_n833));
  AOI211_X1 g408(.A(KEYINPUT106), .B(new_n789), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(G150));
  NAND3_X1  g410(.A1(new_n511), .A2(new_n516), .A3(G93), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  INV_X1    g412(.A(G67), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n507), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n541), .A2(G55), .B1(new_n839), .B2(G651), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n553), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n548), .A2(new_n836), .A3(new_n552), .A4(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT38), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n614), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT107), .B(G860), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n836), .B2(new_n840), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(G145));
  NAND2_X1  g429(.A1(new_n749), .A2(KEYINPUT108), .ZN(new_n855));
  OAI21_X1  g430(.A(G126), .B1(new_n468), .B2(new_n469), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n461), .B1(new_n856), .B2(new_n492), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT4), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n496), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n491), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n729), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n855), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n814), .B(new_n623), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(G106), .A2(G2105), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n486), .A2(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G142), .B2(new_n462), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n700), .B(new_n870), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n865), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(G160), .B(G162), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n633), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n872), .B2(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g453(.A(new_n618), .B(new_n844), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n601), .A2(G299), .A3(new_n605), .ZN(new_n881));
  AOI21_X1  g456(.A(G299), .B1(new_n601), .B2(new_n605), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G299), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n606), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n601), .A2(G299), .A3(new_n605), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n886), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n879), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(G305), .B(new_n819), .ZN(new_n896));
  XNOR2_X1  g471(.A(G303), .B(G288), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(G305), .B(G290), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(KEYINPUT109), .B2(new_n893), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n892), .A2(new_n894), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n895), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n904), .B1(new_n895), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g482(.A(G868), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n841), .A2(new_n596), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(G295));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n909), .ZN(G331));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n912));
  INV_X1    g487(.A(new_n843), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n548), .A2(new_n552), .B1(new_n836), .B2(new_n840), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n912), .B(G286), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  OR3_X1    g490(.A1(new_n520), .A2(new_n529), .A3(new_n912), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n912), .B1(new_n520), .B2(new_n529), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n842), .A3(new_n843), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n915), .A2(G171), .A3(new_n916), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(G171), .A2(new_n916), .ZN(new_n920));
  INV_X1    g495(.A(new_n918), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n917), .B1(new_n842), .B2(new_n843), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n919), .A2(new_n923), .B1(new_n883), .B2(new_n887), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n923), .A2(new_n919), .A3(new_n891), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n903), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n919), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n888), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(new_n919), .A3(new_n891), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n902), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n931), .A2(new_n932), .A3(G37), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n903), .B1(new_n924), .B2(new_n925), .ZN(new_n934));
  INV_X1    g509(.A(G37), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT111), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n927), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n932), .B1(new_n931), .B2(G37), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n934), .A2(KEYINPUT111), .A3(new_n935), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n926), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n931), .A2(G37), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n927), .A2(new_n945), .A3(new_n943), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n938), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI211_X1 g522(.A(KEYINPUT43), .B(new_n926), .C1(new_n940), .C2(new_n941), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n943), .B1(new_n927), .B2(new_n945), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  MUX2_X1   g525(.A(new_n947), .B(new_n950), .S(KEYINPUT44), .Z(G397));
  XNOR2_X1  g526(.A(new_n729), .B(G2067), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n952), .A2(new_n700), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n470), .A2(new_n471), .B1(G113), .B2(G2104), .ZN(new_n954));
  AOI211_X1 g529(.A(KEYINPUT69), .B(new_n461), .C1(new_n954), .C2(new_n473), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n478), .B1(new_n475), .B2(G2105), .ZN(new_n956));
  OAI211_X1 g531(.A(G40), .B(new_n466), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(G164), .B2(G1384), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n953), .A2(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n963), .B2(new_n962), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(new_n822), .A3(new_n819), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT48), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n960), .A2(new_n952), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT113), .Z(new_n971));
  XNOR2_X1  g546(.A(new_n700), .B(G1996), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n960), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n960), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n814), .B(new_n816), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n969), .B1(new_n976), .B2(KEYINPUT126), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(KEYINPUT126), .B2(new_n976), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n814), .A2(new_n817), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n973), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G2067), .B2(new_n729), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n967), .B(new_n978), .C1(new_n960), .C2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1384), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT45), .B1(new_n861), .B2(new_n983), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n958), .B(G1384), .C1(new_n859), .C2(new_n860), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n957), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(G164), .A2(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(G160), .A2(G40), .A3(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT58), .B(G1341), .Z(new_n989));
  AOI22_X1  g564(.A1(new_n986), .A2(new_n961), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT59), .B1(new_n990), .B2(new_n553), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT59), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n993));
  NAND4_X1  g568(.A1(G160), .A2(new_n959), .A3(G40), .A4(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(G1996), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n861), .A2(new_n983), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n957), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n989), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n992), .B(new_n554), .C1(new_n995), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n991), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT61), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT50), .B1(new_n861), .B2(new_n983), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n1004), .B(G1384), .C1(new_n859), .C2(new_n860), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n756), .B1(new_n1006), .B2(new_n957), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n1008));
  XNOR2_X1  g583(.A(G299), .B(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n984), .A2(new_n985), .ZN(new_n1010));
  INV_X1    g585(.A(new_n957), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT56), .B(G2072), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1007), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1009), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1002), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1001), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1007), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT61), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n959), .A2(new_n993), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1012), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1021), .A2(new_n957), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1004), .B1(G164), .B2(G1384), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n861), .A2(KEYINPUT50), .A3(new_n983), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1956), .B1(new_n1026), .B2(new_n1011), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1020), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1007), .A2(KEYINPUT117), .A3(new_n1013), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1009), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1019), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT118), .B1(new_n1017), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1018), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1035), .A2(new_n1002), .B1(new_n991), .B2(new_n1000), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1007), .A2(KEYINPUT117), .A3(new_n1013), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT117), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1031), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1019), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1036), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1026), .A2(new_n1011), .ZN(new_n1044));
  INV_X1    g619(.A(G1348), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1044), .A2(new_n1045), .B1(new_n731), .B2(new_n997), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1046), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n606), .B1(new_n1046), .B2(KEYINPUT60), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1047), .A2(new_n1048), .B1(KEYINPUT60), .B2(new_n1046), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1033), .A2(new_n1043), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1039), .B1(new_n606), .B2(new_n1046), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1018), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n994), .B2(G2078), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT120), .B(new_n1054), .C1(new_n994), .C2(G2078), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1044), .A2(new_n773), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n986), .A2(KEYINPUT53), .A3(new_n737), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G171), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1055), .A2(new_n1056), .B1(new_n773), .B2(new_n1044), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n466), .B(KEYINPUT121), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n737), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1010), .A2(new_n476), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1063), .A2(G301), .A3(new_n1058), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(KEYINPUT122), .A3(new_n1069), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1976), .ZN(new_n1075));
  OAI221_X1 g650(.A(G8), .B1(G288), .B2(new_n1075), .C1(new_n957), .C2(new_n996), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT52), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G303), .A2(G8), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n1082), .B(KEYINPUT55), .Z(new_n1083));
  INV_X1    g658(.A(G8), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n793), .B1(new_n1021), .B2(new_n957), .ZN(new_n1085));
  INV_X1    g660(.A(G2090), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1026), .A2(new_n1011), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1084), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n799), .A2(G1976), .ZN(new_n1090));
  OR3_X1    g665(.A1(new_n1076), .A2(KEYINPUT52), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n583), .A2(new_n584), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G1981), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n583), .A2(new_n586), .A3(new_n685), .A4(new_n587), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT49), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n997), .A2(new_n1084), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n1094), .A3(KEYINPUT49), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1081), .A2(new_n1089), .A3(new_n1091), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1006), .A2(G2084), .A3(new_n957), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1966), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT119), .B(G8), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G168), .A2(new_n1084), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n994), .A2(new_n761), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1026), .A2(new_n1011), .A3(new_n716), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1084), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AND2_X1   g685(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1105), .B(new_n1107), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1110), .B2(new_n1106), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1106), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1085), .A2(new_n1087), .A3(KEYINPUT115), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(G8), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1083), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1117), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1084), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1125));
  AOI211_X1 g700(.A(KEYINPUT116), .B(new_n1083), .C1(new_n1125), .C2(new_n1121), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1102), .B(new_n1116), .C1(new_n1124), .C2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT54), .B1(new_n1061), .B2(G171), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1063), .A2(new_n1058), .A3(new_n1066), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(G171), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1053), .A2(new_n1074), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1102), .B1(new_n1126), .B2(new_n1124), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1112), .A2(new_n1134), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1062), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT123), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1085), .A2(new_n1087), .A3(KEYINPUT115), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT115), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n1084), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT116), .B1(new_n1141), .B2(new_n1083), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1122), .A2(new_n1117), .A3(new_n1123), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1101), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n1136), .A4(new_n1135), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1116), .A2(KEYINPUT62), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1138), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1110), .A2(G168), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1081), .A2(new_n1091), .A3(new_n1100), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT63), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1100), .A2(new_n1075), .A3(new_n799), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1094), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1098), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1157), .B(new_n1149), .C1(new_n1126), .C2(new_n1124), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1089), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1151), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1132), .A2(new_n1148), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n1163));
  XNOR2_X1  g738(.A(G290), .B(G1986), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n976), .B1(new_n960), .B2(new_n1164), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1163), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n982), .B1(new_n1166), .B2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g743(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1170));
  OAI21_X1  g744(.A(new_n1170), .B1(new_n688), .B2(new_n689), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1171), .B1(new_n875), .B2(new_n876), .ZN(new_n1172));
  AND3_X1   g746(.A1(new_n947), .A2(KEYINPUT127), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g747(.A(KEYINPUT127), .B1(new_n947), .B2(new_n1172), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n1173), .A2(new_n1174), .ZN(G308));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n1172), .ZN(new_n1176));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n947), .A2(new_n1172), .A3(KEYINPUT127), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1179), .ZN(G225));
endmodule


