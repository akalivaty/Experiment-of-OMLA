

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582;

  BUF_X2 U322 ( .A(n569), .Z(n290) );
  XOR2_X1 U323 ( .A(n325), .B(n324), .Z(n569) );
  XNOR2_X1 U324 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U325 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U326 ( .A(n307), .B(n341), .ZN(n572) );
  XNOR2_X1 U327 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U328 ( .A(n451), .B(n450), .ZN(G1349GAT) );
  XOR2_X1 U329 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n292) );
  XOR2_X1 U330 ( .A(G176GAT), .B(G92GAT), .Z(n373) );
  XOR2_X1 U331 ( .A(G99GAT), .B(G85GAT), .Z(n352) );
  XNOR2_X1 U332 ( .A(n373), .B(n352), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n298) );
  XOR2_X1 U334 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n294) );
  XNOR2_X1 U335 ( .A(G120GAT), .B(KEYINPUT74), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n296) );
  AND2_X1 U337 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U338 ( .A(KEYINPUT31), .B(n299), .Z(n302) );
  XNOR2_X1 U339 ( .A(G204GAT), .B(G106GAT), .ZN(n300) );
  XNOR2_X1 U340 ( .A(n300), .B(G148GAT), .ZN(n410) );
  XNOR2_X1 U341 ( .A(n410), .B(KEYINPUT33), .ZN(n301) );
  XNOR2_X1 U342 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U343 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n304) );
  XNOR2_X1 U344 ( .A(G71GAT), .B(G57GAT), .ZN(n303) );
  XNOR2_X1 U345 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U346 ( .A(G64GAT), .B(G78GAT), .Z(n305) );
  XNOR2_X1 U347 ( .A(n306), .B(n305), .ZN(n341) );
  XOR2_X1 U348 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n308) );
  XNOR2_X1 U349 ( .A(n572), .B(n308), .ZN(n550) );
  XOR2_X1 U350 ( .A(KEYINPUT108), .B(n550), .Z(n533) );
  XOR2_X1 U351 ( .A(G15GAT), .B(G197GAT), .Z(n310) );
  XNOR2_X1 U352 ( .A(G169GAT), .B(G8GAT), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n325) );
  XOR2_X1 U354 ( .A(G113GAT), .B(G1GAT), .Z(n399) );
  XOR2_X1 U355 ( .A(G29GAT), .B(G43GAT), .Z(n312) );
  XNOR2_X1 U356 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n312), .B(n311), .ZN(n349) );
  XOR2_X1 U358 ( .A(n399), .B(n349), .Z(n314) );
  XNOR2_X1 U359 ( .A(G36GAT), .B(G50GAT), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U361 ( .A(KEYINPUT69), .B(G141GAT), .Z(n316) );
  NAND2_X1 U362 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U364 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U365 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n320) );
  XNOR2_X1 U366 ( .A(KEYINPUT29), .B(G22GAT), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n321), .B(KEYINPUT70), .ZN(n322) );
  XNOR2_X1 U369 ( .A(n323), .B(n322), .ZN(n324) );
  INV_X1 U370 ( .A(n290), .ZN(n499) );
  NOR2_X1 U371 ( .A1(n499), .A2(n550), .ZN(n327) );
  INV_X1 U372 ( .A(KEYINPUT46), .ZN(n326) );
  XNOR2_X1 U373 ( .A(n327), .B(n326), .ZN(n362) );
  XOR2_X1 U374 ( .A(KEYINPUT81), .B(KEYINPUT15), .Z(n329) );
  XNOR2_X1 U375 ( .A(KEYINPUT12), .B(KEYINPUT83), .ZN(n328) );
  XNOR2_X1 U376 ( .A(n329), .B(n328), .ZN(n340) );
  XOR2_X1 U377 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n331) );
  XOR2_X1 U378 ( .A(G15GAT), .B(G127GAT), .Z(n429) );
  XOR2_X1 U379 ( .A(G22GAT), .B(G155GAT), .Z(n411) );
  XNOR2_X1 U380 ( .A(n429), .B(n411), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U382 ( .A(n332), .B(KEYINPUT82), .Z(n338) );
  XNOR2_X1 U383 ( .A(G8GAT), .B(G183GAT), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n333), .B(G211GAT), .ZN(n377) );
  XOR2_X1 U385 ( .A(n377), .B(KEYINPUT84), .Z(n335) );
  NAND2_X1 U386 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U388 ( .A(G1GAT), .B(n336), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n342) );
  XNOR2_X1 U391 ( .A(n342), .B(n341), .ZN(n575) );
  XNOR2_X1 U392 ( .A(KEYINPUT116), .B(n575), .ZN(n557) );
  XOR2_X1 U393 ( .A(KEYINPUT78), .B(G106GAT), .Z(n344) );
  XNOR2_X1 U394 ( .A(G134GAT), .B(G92GAT), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n360) );
  XOR2_X1 U396 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n346) );
  NAND2_X1 U397 ( .A1(G232GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U399 ( .A(n347), .B(KEYINPUT66), .Z(n351) );
  XNOR2_X1 U400 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n348), .B(G162GAT), .ZN(n420) );
  XNOR2_X1 U402 ( .A(n349), .B(n420), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n356) );
  XOR2_X1 U404 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n354) );
  XOR2_X1 U405 ( .A(G36GAT), .B(G190GAT), .Z(n374) );
  XNOR2_X1 U406 ( .A(n352), .B(n374), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U408 ( .A(n356), .B(n355), .Z(n358) );
  XNOR2_X1 U409 ( .A(G218GAT), .B(KEYINPUT79), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U411 ( .A(n360), .B(n359), .Z(n452) );
  INV_X1 U412 ( .A(n452), .ZN(n562) );
  NOR2_X1 U413 ( .A1(n557), .A2(n562), .ZN(n361) );
  NAND2_X1 U414 ( .A1(n362), .A2(n361), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n363), .B(KEYINPUT47), .ZN(n368) );
  INV_X1 U416 ( .A(n575), .ZN(n483) );
  XNOR2_X1 U417 ( .A(KEYINPUT36), .B(n452), .ZN(n580) );
  NOR2_X1 U418 ( .A1(n483), .A2(n580), .ZN(n364) );
  XNOR2_X1 U419 ( .A(KEYINPUT45), .B(n364), .ZN(n365) );
  NAND2_X1 U420 ( .A1(n365), .A2(n572), .ZN(n366) );
  NOR2_X1 U421 ( .A1(n366), .A2(n290), .ZN(n367) );
  NOR2_X1 U422 ( .A1(n368), .A2(n367), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n369), .B(KEYINPUT48), .ZN(n527) );
  XOR2_X1 U424 ( .A(KEYINPUT96), .B(G204GAT), .Z(n371) );
  NAND2_X1 U425 ( .A1(G226GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U427 ( .A(n372), .B(G64GAT), .Z(n376) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n378) );
  XOR2_X1 U430 ( .A(n378), .B(n377), .Z(n384) );
  XOR2_X1 U431 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n380) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n433) );
  XOR2_X1 U434 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n382) );
  XNOR2_X1 U435 ( .A(G197GAT), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n421) );
  XNOR2_X1 U437 ( .A(n433), .B(n421), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n475) );
  NOR2_X1 U439 ( .A1(n527), .A2(n475), .ZN(n386) );
  XNOR2_X1 U440 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n408) );
  XOR2_X1 U442 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n388) );
  XNOR2_X1 U443 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n407) );
  XOR2_X1 U445 ( .A(G162GAT), .B(G85GAT), .Z(n390) );
  XNOR2_X1 U446 ( .A(G29GAT), .B(G148GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U448 ( .A(KEYINPUT95), .B(G155GAT), .Z(n392) );
  XNOR2_X1 U449 ( .A(G127GAT), .B(G57GAT), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U451 ( .A(n394), .B(n393), .Z(n405) );
  XOR2_X1 U452 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n396) );
  XNOR2_X1 U453 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(KEYINPUT92), .B(n397), .ZN(n426) );
  INV_X1 U456 ( .A(n426), .ZN(n403) );
  XNOR2_X1 U457 ( .A(G134GAT), .B(G120GAT), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n398), .B(KEYINPUT0), .ZN(n430) );
  XOR2_X1 U459 ( .A(n430), .B(n399), .Z(n401) );
  NAND2_X1 U460 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n543) );
  NOR2_X1 U465 ( .A1(n408), .A2(n543), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n409), .B(KEYINPUT65), .ZN(n568) );
  XOR2_X1 U467 ( .A(n411), .B(n410), .Z(n413) );
  NAND2_X1 U468 ( .A1(G228GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n425) );
  XOR2_X1 U470 ( .A(KEYINPUT94), .B(KEYINPUT89), .Z(n415) );
  XNOR2_X1 U471 ( .A(G211GAT), .B(G78GAT), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U473 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n417) );
  XNOR2_X1 U474 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U476 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n464) );
  NOR2_X1 U481 ( .A1(n568), .A2(n464), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n428), .B(KEYINPUT55), .ZN(n446) );
  XOR2_X1 U483 ( .A(n430), .B(n429), .Z(n432) );
  XNOR2_X1 U484 ( .A(G99GAT), .B(G190GAT), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n437) );
  XOR2_X1 U486 ( .A(n433), .B(KEYINPUT20), .Z(n435) );
  NAND2_X1 U487 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U489 ( .A(n437), .B(n436), .Z(n445) );
  XOR2_X1 U490 ( .A(G71GAT), .B(G176GAT), .Z(n439) );
  XNOR2_X1 U491 ( .A(G43GAT), .B(G183GAT), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U493 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n441) );
  XNOR2_X1 U494 ( .A(G113GAT), .B(KEYINPUT88), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n528) );
  NOR2_X1 U498 ( .A1(n446), .A2(n528), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n447), .B(KEYINPUT122), .ZN(n563) );
  NAND2_X1 U500 ( .A1(n533), .A2(n563), .ZN(n451) );
  XOR2_X1 U501 ( .A(G176GAT), .B(KEYINPUT57), .Z(n449) );
  XOR2_X1 U502 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n448) );
  XOR2_X1 U503 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n473) );
  NAND2_X1 U504 ( .A1(n290), .A2(n572), .ZN(n487) );
  NAND2_X1 U505 ( .A1(n575), .A2(n452), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n453), .B(KEYINPUT85), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(KEYINPUT16), .ZN(n471) );
  XOR2_X1 U508 ( .A(n475), .B(KEYINPUT97), .Z(n455) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(n455), .ZN(n462) );
  XNOR2_X1 U510 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n456), .B(n464), .ZN(n479) );
  NAND2_X1 U512 ( .A1(n543), .A2(n479), .ZN(n457) );
  NOR2_X1 U513 ( .A1(n462), .A2(n457), .ZN(n530) );
  XNOR2_X1 U514 ( .A(n530), .B(KEYINPUT98), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n458), .A2(n528), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(KEYINPUT99), .ZN(n469) );
  NAND2_X1 U517 ( .A1(n464), .A2(n528), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(KEYINPUT26), .ZN(n461) );
  XNOR2_X1 U519 ( .A(KEYINPUT100), .B(n461), .ZN(n567) );
  NOR2_X1 U520 ( .A1(n567), .A2(n462), .ZN(n544) );
  NOR2_X1 U521 ( .A1(n528), .A2(n475), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  NOR2_X1 U524 ( .A1(n544), .A2(n466), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n543), .A2(n467), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U527 ( .A(KEYINPUT101), .B(n470), .ZN(n482) );
  NAND2_X1 U528 ( .A1(n471), .A2(n482), .ZN(n500) );
  NOR2_X1 U529 ( .A1(n487), .A2(n500), .ZN(n480) );
  NAND2_X1 U530 ( .A1(n480), .A2(n543), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U532 ( .A(G1GAT), .B(n474), .Z(G1324GAT) );
  INV_X1 U533 ( .A(n475), .ZN(n517) );
  NAND2_X1 U534 ( .A1(n517), .A2(n480), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  INV_X1 U537 ( .A(n528), .ZN(n520) );
  NAND2_X1 U538 ( .A1(n480), .A2(n520), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  INV_X1 U540 ( .A(n479), .ZN(n522) );
  NAND2_X1 U541 ( .A1(n480), .A2(n522), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U543 ( .A1(n483), .A2(n482), .ZN(n484) );
  NOR2_X1 U544 ( .A1(n580), .A2(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n485) );
  XOR2_X1 U546 ( .A(n486), .B(n485), .Z(n515) );
  OR2_X1 U547 ( .A1(n487), .A2(n515), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(n488), .Z(n497) );
  NAND2_X1 U549 ( .A1(n543), .A2(n497), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n491), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n517), .A2(n497), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  XNOR2_X1 U555 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n496) );
  XOR2_X1 U556 ( .A(G43GAT), .B(KEYINPUT105), .Z(n494) );
  NAND2_X1 U557 ( .A1(n497), .A2(n520), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n497), .A2(n522), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT107), .Z(n502) );
  NAND2_X1 U563 ( .A1(n499), .A2(n533), .ZN(n514) );
  NOR2_X1 U564 ( .A1(n514), .A2(n500), .ZN(n510) );
  NAND2_X1 U565 ( .A1(n510), .A2(n543), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n517), .A2(n510), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n520), .A2(n510), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT111), .B(KEYINPUT113), .Z(n509) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT112), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n513) );
  NAND2_X1 U577 ( .A1(n510), .A2(n522), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n523), .A2(n543), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n523), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT114), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n519), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n520), .A2(n523), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n525) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U592 ( .A1(n527), .A2(n528), .ZN(n529) );
  NAND2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U594 ( .A(KEYINPUT117), .B(n531), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n540), .A2(n290), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n532), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U598 ( .A1(n540), .A2(n533), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n538) );
  NAND2_X1 U602 ( .A1(n540), .A2(n557), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n562), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U609 ( .A1(n527), .A2(n545), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n554), .A2(n290), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n552) );
  INV_X1 U615 ( .A(n554), .ZN(n549) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(n552), .B(n551), .Z(G1345GAT) );
  NAND2_X1 U618 ( .A1(n575), .A2(n554), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n562), .A2(n554), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n563), .A2(n290), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT124), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(n559), .ZN(G1350GAT) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(KEYINPUT125), .ZN(n561) );
  XOR2_X1 U629 ( .A(KEYINPUT126), .B(n561), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT59), .ZN(n571) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n576), .A2(n290), .ZN(n570) );
  XOR2_X1 U636 ( .A(n571), .B(n570), .Z(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U638 ( .A(n576), .ZN(n579) );
  OR2_X1 U639 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT127), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

