

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789;

  BUF_X1 U380 ( .A(n674), .Z(n357) );
  INV_X1 U381 ( .A(n602), .ZN(n684) );
  NAND2_X2 U382 ( .A1(n453), .A2(n450), .ZN(n383) );
  XNOR2_X1 U383 ( .A(n439), .B(n534), .ZN(n757) );
  NOR2_X1 U384 ( .A1(n626), .A2(n697), .ZN(n627) );
  AND2_X1 U385 ( .A1(n646), .A2(n356), .ZN(n421) );
  NAND2_X1 U386 ( .A1(n424), .A2(n643), .ZN(n356) );
  NOR2_X1 U387 ( .A1(n783), .A2(n789), .ZN(n579) );
  INV_X2 U388 ( .A(G953), .ZN(n775) );
  AND2_X1 U389 ( .A1(n644), .A2(n642), .ZN(n424) );
  BUF_X2 U390 ( .A(n754), .Z(n358) );
  NOR2_X2 U391 ( .A1(n749), .A2(n756), .ZN(n443) );
  NAND2_X2 U392 ( .A1(n374), .A2(n376), .ZN(n380) );
  XNOR2_X2 U393 ( .A(n561), .B(n550), .ZN(n770) );
  XNOR2_X2 U394 ( .A(n536), .B(G134), .ZN(n561) );
  NAND2_X1 U395 ( .A1(n697), .A2(n696), .ZN(n701) );
  XNOR2_X2 U396 ( .A(n516), .B(n758), .ZN(n533) );
  INV_X1 U397 ( .A(KEYINPUT35), .ZN(n623) );
  INV_X1 U398 ( .A(G475), .ZN(n417) );
  NOR2_X1 U399 ( .A1(n737), .A2(n417), .ZN(n414) );
  AND2_X1 U400 ( .A1(n391), .A2(n390), .ZN(n668) );
  NOR2_X1 U401 ( .A1(n655), .A2(n664), .ZN(n420) );
  NOR2_X1 U402 ( .A1(n624), .A2(KEYINPUT71), .ZN(n639) );
  XNOR2_X1 U403 ( .A(n631), .B(n630), .ZN(n636) );
  AND2_X1 U404 ( .A1(n525), .A2(n423), .ZN(n438) );
  XNOR2_X1 U405 ( .A(n499), .B(n498), .ZN(n562) );
  XOR2_X1 U406 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n499) );
  NAND2_X1 U407 ( .A1(n588), .A2(n712), .ZN(n359) );
  NAND2_X1 U408 ( .A1(n588), .A2(n712), .ZN(n382) );
  XOR2_X2 U409 ( .A(KEYINPUT4), .B(KEYINPUT65), .Z(n771) );
  XNOR2_X1 U410 ( .A(n359), .B(KEYINPUT19), .ZN(n360) );
  XNOR2_X1 U411 ( .A(n382), .B(KEYINPUT19), .ZN(n618) );
  XNOR2_X1 U412 ( .A(n669), .B(n446), .ZN(n445) );
  NAND2_X1 U413 ( .A1(n421), .A2(n420), .ZN(n419) );
  NOR2_X1 U414 ( .A1(n658), .A2(n592), .ZN(n610) );
  NOR2_X1 U415 ( .A1(n447), .A2(n737), .ZN(n754) );
  NOR2_X1 U416 ( .A1(n394), .A2(n393), .ZN(n392) );
  INV_X1 U417 ( .A(n589), .ZN(n423) );
  XNOR2_X1 U418 ( .A(n574), .B(n425), .ZN(n714) );
  INV_X1 U419 ( .A(KEYINPUT112), .ZN(n425) );
  NAND2_X2 U420 ( .A1(n402), .A2(n399), .ZN(n587) );
  NAND2_X1 U421 ( .A1(n401), .A2(n400), .ZN(n399) );
  AND2_X1 U422 ( .A1(n404), .A2(n403), .ZN(n402) );
  NOR2_X1 U423 ( .A1(n362), .A2(G902), .ZN(n400) );
  XNOR2_X1 U424 ( .A(KEYINPUT70), .B(G101), .ZN(n485) );
  XNOR2_X1 U425 ( .A(n770), .B(G146), .ZN(n384) );
  XNOR2_X1 U426 ( .A(n409), .B(n408), .ZN(n439) );
  INV_X1 U427 ( .A(KEYINPUT16), .ZN(n408) );
  AND2_X1 U428 ( .A1(n455), .A2(n454), .ZN(n453) );
  NAND2_X1 U429 ( .A1(G472), .A2(n452), .ZN(n451) );
  XNOR2_X1 U430 ( .A(n579), .B(n371), .ZN(n395) );
  XNOR2_X1 U431 ( .A(n587), .B(n586), .ZN(n625) );
  XNOR2_X1 U432 ( .A(n541), .B(n542), .ZN(n483) );
  BUF_X1 U433 ( .A(n625), .Z(n441) );
  XNOR2_X1 U434 ( .A(n526), .B(n428), .ZN(n422) );
  INV_X1 U435 ( .A(KEYINPUT30), .ZN(n428) );
  NOR2_X1 U436 ( .A1(G953), .A2(G237), .ZN(n545) );
  XOR2_X1 U437 ( .A(KEYINPUT5), .B(KEYINPUT80), .Z(n520) );
  XNOR2_X1 U438 ( .A(G137), .B(G116), .ZN(n519) );
  INV_X1 U439 ( .A(G122), .ZN(n410) );
  NOR2_X1 U440 ( .A1(n774), .A2(n367), .ZN(n481) );
  XNOR2_X1 U441 ( .A(n364), .B(n533), .ZN(n474) );
  XNOR2_X1 U442 ( .A(n514), .B(n427), .ZN(n406) );
  INV_X1 U443 ( .A(KEYINPUT28), .ZN(n437) );
  XNOR2_X1 U444 ( .A(KEYINPUT117), .B(KEYINPUT41), .ZN(n575) );
  NOR2_X1 U445 ( .A1(n715), .A2(n714), .ZN(n576) );
  AND2_X1 U446 ( .A1(n528), .A2(n365), .ZN(n464) );
  NAND2_X1 U447 ( .A1(n465), .A2(n462), .ZN(n461) );
  NOR2_X1 U448 ( .A1(n467), .A2(n365), .ZN(n465) );
  BUF_X1 U449 ( .A(n588), .Z(n593) );
  INV_X1 U450 ( .A(n441), .ZN(n702) );
  NOR2_X1 U451 ( .A1(n714), .A2(n628), .ZN(n629) );
  INV_X1 U452 ( .A(KEYINPUT6), .ZN(n426) );
  NOR2_X1 U453 ( .A1(n716), .A2(n603), .ZN(n605) );
  NAND2_X1 U454 ( .A1(n609), .A2(n388), .ZN(n393) );
  AND2_X1 U455 ( .A1(n608), .A2(n385), .ZN(n386) );
  AND2_X1 U456 ( .A1(n609), .A2(n694), .ZN(n385) );
  NAND2_X1 U457 ( .A1(n694), .A2(n388), .ZN(n387) );
  OR2_X1 U458 ( .A1(G237), .A2(G902), .ZN(n540) );
  NAND2_X1 U459 ( .A1(n362), .A2(G902), .ZN(n403) );
  XOR2_X1 U460 ( .A(KEYINPUT103), .B(KEYINPUT20), .Z(n506) );
  XOR2_X1 U461 ( .A(G140), .B(KEYINPUT11), .Z(n544) );
  XNOR2_X1 U462 ( .A(KEYINPUT12), .B(KEYINPUT108), .ZN(n543) );
  XOR2_X1 U463 ( .A(KEYINPUT10), .B(n537), .Z(n553) );
  XOR2_X1 U464 ( .A(G122), .B(G104), .Z(n551) );
  XOR2_X1 U465 ( .A(G143), .B(G113), .Z(n547) );
  XNOR2_X1 U466 ( .A(G902), .B(KEYINPUT15), .ZN(n665) );
  INV_X1 U467 ( .A(G107), .ZN(n427) );
  XNOR2_X1 U468 ( .A(n405), .B(G137), .ZN(n513) );
  INV_X1 U469 ( .A(G140), .ZN(n405) );
  NAND2_X1 U470 ( .A1(n711), .A2(n468), .ZN(n467) );
  NAND2_X1 U471 ( .A1(n572), .A2(n696), .ZN(n589) );
  NAND2_X1 U472 ( .A1(G214), .A2(n540), .ZN(n712) );
  INV_X1 U473 ( .A(KEYINPUT79), .ZN(n430) );
  INV_X1 U474 ( .A(n701), .ZN(n469) );
  INV_X1 U475 ( .A(G902), .ZN(n452) );
  NAND2_X1 U476 ( .A1(n457), .A2(G902), .ZN(n454) );
  XNOR2_X1 U477 ( .A(n557), .B(n556), .ZN(n596) );
  XNOR2_X1 U478 ( .A(G110), .B(KEYINPUT76), .ZN(n500) );
  XNOR2_X1 U479 ( .A(G128), .B(G119), .ZN(n496) );
  XNOR2_X1 U480 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n558) );
  XOR2_X1 U481 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n559) );
  XNOR2_X1 U482 ( .A(n434), .B(n535), .ZN(n673) );
  XNOR2_X1 U483 ( .A(n757), .B(n539), .ZN(n434) );
  NAND2_X1 U484 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U485 ( .A1(n719), .A2(KEYINPUT34), .ZN(n377) );
  NAND2_X1 U486 ( .A1(n379), .A2(n622), .ZN(n375) );
  INV_X1 U487 ( .A(KEYINPUT114), .ZN(n456) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n597) );
  INV_X1 U489 ( .A(G478), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n436), .B(n524), .ZN(n674) );
  XNOR2_X1 U491 ( .A(n384), .B(n516), .ZN(n436) );
  NAND2_X1 U492 ( .A1(n412), .A2(n411), .ZN(n473) );
  XNOR2_X1 U493 ( .A(G104), .B(G110), .ZN(n758) );
  XNOR2_X1 U494 ( .A(n746), .B(n488), .ZN(n747) );
  XNOR2_X1 U495 ( .A(n578), .B(n577), .ZN(n789) );
  XNOR2_X1 U496 ( .A(n570), .B(n569), .ZN(n783) );
  AND2_X1 U497 ( .A1(n458), .A2(n461), .ZN(n570) );
  XNOR2_X1 U498 ( .A(n594), .B(n440), .ZN(n595) );
  XNOR2_X1 U499 ( .A(KEYINPUT36), .B(KEYINPUT118), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n634), .B(n635), .ZN(n787) );
  AND2_X1 U501 ( .A1(n622), .A2(n468), .ZN(n429) );
  XNOR2_X1 U502 ( .A(n653), .B(KEYINPUT107), .ZN(n676) );
  XNOR2_X1 U503 ( .A(n398), .B(n397), .ZN(n396) );
  XNOR2_X1 U504 ( .A(n741), .B(n742), .ZN(n743) );
  AND2_X1 U505 ( .A1(n650), .A2(KEYINPUT34), .ZN(n361) );
  XOR2_X1 U506 ( .A(KEYINPUT74), .B(G469), .Z(n362) );
  INV_X1 U507 ( .A(n571), .ZN(n468) );
  NOR2_X2 U508 ( .A1(n597), .A2(n567), .ZN(n687) );
  XOR2_X1 U509 ( .A(KEYINPUT82), .B(KEYINPUT23), .Z(n363) );
  XOR2_X1 U510 ( .A(n406), .B(n513), .Z(n364) );
  XNOR2_X1 U511 ( .A(n598), .B(KEYINPUT115), .ZN(n622) );
  XOR2_X1 U512 ( .A(KEYINPUT92), .B(KEYINPUT39), .Z(n365) );
  XOR2_X1 U513 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n366) );
  AND2_X1 U514 ( .A1(n665), .A2(n482), .ZN(n367) );
  OR2_X1 U515 ( .A1(n665), .A2(n482), .ZN(n368) );
  XOR2_X1 U516 ( .A(n673), .B(n672), .Z(n369) );
  XOR2_X1 U517 ( .A(n357), .B(KEYINPUT62), .Z(n370) );
  XOR2_X1 U518 ( .A(KEYINPUT46), .B(KEYINPUT91), .Z(n371) );
  INV_X1 U519 ( .A(KEYINPUT48), .ZN(n388) );
  XOR2_X1 U520 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n372) );
  NOR2_X1 U521 ( .A1(G952), .A2(n775), .ZN(n756) );
  INV_X1 U522 ( .A(n756), .ZN(n471) );
  OR2_X1 U523 ( .A1(n665), .A2(n731), .ZN(n373) );
  INV_X1 U524 ( .A(G472), .ZN(n457) );
  NOR2_X2 U525 ( .A1(n361), .A2(n375), .ZN(n374) );
  NAND2_X1 U526 ( .A1(n377), .A2(n378), .ZN(n376) );
  INV_X1 U527 ( .A(n650), .ZN(n378) );
  NAND2_X1 U528 ( .A1(n719), .A2(KEYINPUT34), .ZN(n379) );
  XNOR2_X2 U529 ( .A(n380), .B(n623), .ZN(n786) );
  AND2_X2 U530 ( .A1(n448), .A2(n373), .ZN(n447) );
  NAND2_X1 U531 ( .A1(n358), .A2(G217), .ZN(n398) );
  XNOR2_X1 U532 ( .A(n473), .B(n370), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n444), .A2(n445), .ZN(n381) );
  NOR2_X1 U534 ( .A1(n692), .A2(n683), .ZN(n600) );
  XNOR2_X2 U535 ( .A(n381), .B(KEYINPUT81), .ZN(n737) );
  NAND2_X1 U536 ( .A1(n699), .A2(n383), .ZN(n700) );
  XNOR2_X2 U537 ( .A(n383), .B(n456), .ZN(n525) );
  XNOR2_X2 U538 ( .A(n383), .B(n426), .ZN(n658) );
  NOR2_X1 U539 ( .A1(n647), .A2(n383), .ZN(n707) );
  NAND2_X1 U540 ( .A1(n652), .A2(n383), .ZN(n653) );
  XNOR2_X1 U541 ( .A(n474), .B(n384), .ZN(n741) );
  NAND2_X1 U542 ( .A1(n395), .A2(n386), .ZN(n389) );
  NAND2_X1 U543 ( .A1(n389), .A2(n387), .ZN(n391) );
  NAND2_X1 U544 ( .A1(n392), .A2(n395), .ZN(n390) );
  INV_X1 U545 ( .A(n608), .ZN(n394) );
  AND2_X1 U546 ( .A1(n396), .A2(n471), .ZN(G66) );
  INV_X1 U547 ( .A(n755), .ZN(n397) );
  INV_X1 U548 ( .A(n741), .ZN(n401) );
  NAND2_X1 U549 ( .A1(n741), .A2(n362), .ZN(n404) );
  NAND2_X1 U550 ( .A1(n407), .A2(n629), .ZN(n631) );
  NAND2_X1 U551 ( .A1(n707), .A2(n407), .ZN(n648) );
  XNOR2_X2 U552 ( .A(n407), .B(KEYINPUT99), .ZN(n650) );
  XNOR2_X2 U553 ( .A(n620), .B(n619), .ZN(n407) );
  XNOR2_X1 U554 ( .A(n409), .B(n565), .ZN(n752) );
  XNOR2_X2 U555 ( .A(n442), .B(n410), .ZN(n409) );
  INV_X1 U556 ( .A(n447), .ZN(n411) );
  NOR2_X1 U557 ( .A1(n737), .A2(n457), .ZN(n412) );
  NAND2_X1 U558 ( .A1(n414), .A2(n413), .ZN(n748) );
  INV_X1 U559 ( .A(n447), .ZN(n413) );
  NAND2_X1 U560 ( .A1(n415), .A2(n411), .ZN(n477) );
  NOR2_X1 U561 ( .A1(n737), .A2(n416), .ZN(n415) );
  INV_X1 U562 ( .A(G210), .ZN(n416) );
  XNOR2_X1 U563 ( .A(n502), .B(n503), .ZN(n504) );
  NAND2_X1 U564 ( .A1(n562), .A2(G221), .ZN(n501) );
  XNOR2_X2 U565 ( .A(n418), .B(n510), .ZN(n697) );
  NOR2_X2 U566 ( .A1(n755), .A2(G902), .ZN(n418) );
  XNOR2_X2 U567 ( .A(n419), .B(n366), .ZN(n762) );
  NAND2_X1 U568 ( .A1(n422), .A2(n527), .ZN(n528) );
  NAND2_X1 U569 ( .A1(n673), .A2(n665), .ZN(n484) );
  INV_X1 U570 ( .A(n525), .ZN(n637) );
  NOR2_X2 U571 ( .A1(n787), .A2(n680), .ZN(n644) );
  NAND2_X1 U572 ( .A1(n636), .A2(n632), .ZN(n633) );
  NOR2_X2 U573 ( .A1(n647), .A2(n658), .ZN(n621) );
  NOR2_X2 U574 ( .A1(n587), .A2(n573), .ZN(n581) );
  NAND2_X1 U575 ( .A1(n674), .A2(n457), .ZN(n455) );
  NAND2_X1 U576 ( .A1(n462), .A2(n429), .ZN(n599) );
  XNOR2_X2 U577 ( .A(n621), .B(KEYINPUT33), .ZN(n719) );
  XNOR2_X2 U578 ( .A(n431), .B(n430), .ZN(n647) );
  NAND2_X1 U579 ( .A1(n469), .A2(n625), .ZN(n431) );
  NOR2_X1 U580 ( .A1(n752), .A2(G902), .ZN(n433) );
  XNOR2_X2 U581 ( .A(n484), .B(n483), .ZN(n588) );
  BUF_X1 U582 ( .A(n762), .Z(n435) );
  INV_X2 U583 ( .A(n593), .ZN(n612) );
  XNOR2_X1 U584 ( .A(n438), .B(n437), .ZN(n573) );
  XNOR2_X2 U585 ( .A(G107), .B(G116), .ZN(n442) );
  XNOR2_X2 U586 ( .A(n612), .B(KEYINPUT38), .ZN(n711) );
  XNOR2_X1 U587 ( .A(n443), .B(n750), .ZN(G60) );
  XNOR2_X1 U588 ( .A(n576), .B(n575), .ZN(n695) );
  NAND2_X1 U589 ( .A1(n479), .A2(n478), .ZN(n449) );
  XNOR2_X2 U590 ( .A(G143), .B(G128), .ZN(n536) );
  INV_X1 U591 ( .A(n762), .ZN(n444) );
  INV_X1 U592 ( .A(KEYINPUT90), .ZN(n446) );
  NAND2_X1 U593 ( .A1(n449), .A2(n481), .ZN(n448) );
  OR2_X1 U594 ( .A1(n674), .A2(n451), .ZN(n450) );
  NOR2_X1 U595 ( .A1(n464), .A2(n463), .ZN(n458) );
  NAND2_X1 U596 ( .A1(n459), .A2(n461), .ZN(n568) );
  NOR2_X1 U597 ( .A1(n464), .A2(n460), .ZN(n459) );
  INV_X1 U598 ( .A(n466), .ZN(n460) );
  INV_X1 U599 ( .A(n528), .ZN(n462) );
  NAND2_X1 U600 ( .A1(n466), .A2(n687), .ZN(n463) );
  NAND2_X1 U601 ( .A1(n467), .A2(n365), .ZN(n466) );
  XNOR2_X1 U602 ( .A(n477), .B(n369), .ZN(n476) );
  XNOR2_X1 U603 ( .A(n470), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U604 ( .A1(n472), .A2(n471), .ZN(n470) );
  XNOR2_X1 U605 ( .A(n475), .B(n372), .ZN(G51) );
  NAND2_X1 U606 ( .A1(n476), .A2(n471), .ZN(n475) );
  NAND2_X1 U607 ( .A1(n762), .A2(KEYINPUT89), .ZN(n478) );
  NAND2_X1 U608 ( .A1(n480), .A2(n368), .ZN(n479) );
  INV_X1 U609 ( .A(n762), .ZN(n480) );
  INV_X1 U610 ( .A(KEYINPUT89), .ZN(n482) );
  XNOR2_X2 U611 ( .A(n771), .B(n485), .ZN(n516) );
  XOR2_X1 U612 ( .A(n487), .B(n500), .Z(n486) );
  XOR2_X1 U613 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n487) );
  XNOR2_X1 U614 ( .A(KEYINPUT125), .B(KEYINPUT59), .ZN(n488) );
  INV_X1 U615 ( .A(n788), .ZN(n662) );
  NAND2_X1 U616 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n586) );
  XNOR2_X1 U619 ( .A(KEYINPUT77), .B(KEYINPUT22), .ZN(n630) );
  XNOR2_X1 U620 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U621 ( .A(n748), .B(n747), .ZN(n749) );
  INV_X1 U622 ( .A(KEYINPUT42), .ZN(n577) );
  XNOR2_X1 U623 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U624 ( .A1(G234), .A2(G237), .ZN(n489) );
  XNOR2_X1 U625 ( .A(n489), .B(KEYINPUT14), .ZN(n491) );
  NAND2_X1 U626 ( .A1(n491), .A2(G952), .ZN(n490) );
  XNOR2_X1 U627 ( .A(n490), .B(KEYINPUT97), .ZN(n726) );
  NAND2_X1 U628 ( .A1(n726), .A2(n775), .ZN(n615) );
  INV_X1 U629 ( .A(n615), .ZN(n495) );
  NAND2_X1 U630 ( .A1(n491), .A2(G902), .ZN(n492) );
  XOR2_X1 U631 ( .A(KEYINPUT98), .B(n492), .Z(n614) );
  NAND2_X1 U632 ( .A1(n614), .A2(G953), .ZN(n493) );
  NOR2_X1 U633 ( .A1(G900), .A2(n493), .ZN(n494) );
  NOR2_X1 U634 ( .A1(n495), .A2(n494), .ZN(n571) );
  XOR2_X2 U635 ( .A(G146), .B(G125), .Z(n537) );
  XNOR2_X1 U636 ( .A(n553), .B(n513), .ZN(n773) );
  XNOR2_X1 U637 ( .A(n363), .B(n496), .ZN(n497) );
  XOR2_X1 U638 ( .A(KEYINPUT24), .B(n497), .Z(n503) );
  NAND2_X1 U639 ( .A1(G234), .A2(n775), .ZN(n498) );
  XNOR2_X1 U640 ( .A(n501), .B(n486), .ZN(n502) );
  XNOR2_X1 U641 ( .A(n504), .B(n773), .ZN(n755) );
  NAND2_X1 U642 ( .A1(G234), .A2(n665), .ZN(n505) );
  XNOR2_X1 U643 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U644 ( .A(KEYINPUT102), .B(n507), .ZN(n511) );
  NAND2_X1 U645 ( .A1(G217), .A2(n511), .ZN(n509) );
  XNOR2_X1 U646 ( .A(KEYINPUT25), .B(KEYINPUT104), .ZN(n508) );
  NAND2_X1 U647 ( .A1(G221), .A2(n511), .ZN(n512) );
  XNOR2_X1 U648 ( .A(KEYINPUT21), .B(n512), .ZN(n628) );
  INV_X1 U649 ( .A(n628), .ZN(n696) );
  XOR2_X1 U650 ( .A(KEYINPUT73), .B(G131), .Z(n550) );
  NAND2_X1 U651 ( .A1(G227), .A2(n775), .ZN(n514) );
  NOR2_X1 U652 ( .A1(n701), .A2(n587), .ZN(n515) );
  XNOR2_X1 U653 ( .A(n515), .B(KEYINPUT105), .ZN(n649) );
  INV_X1 U654 ( .A(n649), .ZN(n527) );
  XOR2_X1 U655 ( .A(G119), .B(KEYINPUT75), .Z(n518) );
  XNOR2_X1 U656 ( .A(G113), .B(KEYINPUT3), .ZN(n517) );
  XNOR2_X1 U657 ( .A(n518), .B(n517), .ZN(n534) );
  XNOR2_X1 U658 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U659 ( .A(n534), .B(n521), .Z(n523) );
  NAND2_X1 U660 ( .A1(n545), .A2(G210), .ZN(n522) );
  XNOR2_X1 U661 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U662 ( .A1(n712), .A2(n525), .ZN(n526) );
  XOR2_X1 U663 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n530) );
  NAND2_X1 U664 ( .A1(G224), .A2(n775), .ZN(n529) );
  XNOR2_X1 U665 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U666 ( .A(n531), .B(KEYINPUT95), .Z(n532) );
  XNOR2_X1 U667 ( .A(n533), .B(n532), .ZN(n535) );
  INV_X1 U668 ( .A(n536), .ZN(n538) );
  XNOR2_X1 U669 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U670 ( .A1(G210), .A2(n540), .ZN(n541) );
  INV_X1 U671 ( .A(KEYINPUT96), .ZN(n542) );
  XNOR2_X1 U672 ( .A(KEYINPUT13), .B(G475), .ZN(n557) );
  XNOR2_X1 U673 ( .A(n544), .B(n543), .ZN(n549) );
  NAND2_X1 U674 ( .A1(G214), .A2(n545), .ZN(n546) );
  XNOR2_X1 U675 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U676 ( .A(n549), .B(n548), .ZN(n555) );
  XNOR2_X1 U677 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U678 ( .A(n555), .B(n554), .ZN(n746) );
  NOR2_X1 U679 ( .A1(G902), .A2(n746), .ZN(n556) );
  XNOR2_X1 U680 ( .A(n596), .B(KEYINPUT109), .ZN(n567) );
  XNOR2_X1 U681 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U682 ( .A(n561), .B(n560), .Z(n564) );
  NAND2_X1 U683 ( .A1(G217), .A2(n562), .ZN(n563) );
  XNOR2_X1 U684 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U685 ( .A1(n567), .A2(n597), .ZN(n580) );
  NOR2_X1 U686 ( .A1(n568), .A2(n580), .ZN(n566) );
  XOR2_X1 U687 ( .A(KEYINPUT119), .B(n566), .Z(n785) );
  INV_X1 U688 ( .A(n785), .ZN(n666) );
  INV_X1 U689 ( .A(n687), .ZN(n590) );
  XNOR2_X1 U690 ( .A(KEYINPUT116), .B(KEYINPUT40), .ZN(n569) );
  NOR2_X1 U691 ( .A1(n697), .A2(n571), .ZN(n572) );
  NOR2_X1 U692 ( .A1(n596), .A2(n597), .ZN(n574) );
  NAND2_X1 U693 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U694 ( .A1(n581), .A2(n695), .ZN(n578) );
  INV_X1 U695 ( .A(n580), .ZN(n689) );
  NOR2_X1 U696 ( .A1(n689), .A2(n687), .ZN(n716) );
  INV_X1 U697 ( .A(n716), .ZN(n583) );
  NAND2_X1 U698 ( .A1(n360), .A2(n581), .ZN(n602) );
  NOR2_X1 U699 ( .A1(KEYINPUT47), .A2(n602), .ZN(n582) );
  NAND2_X1 U700 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U701 ( .A(n584), .B(KEYINPUT78), .ZN(n609) );
  NAND2_X1 U702 ( .A1(n602), .A2(KEYINPUT47), .ZN(n585) );
  NAND2_X1 U703 ( .A1(n585), .A2(KEYINPUT87), .ZN(n601) );
  NOR2_X1 U704 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U705 ( .A1(n591), .A2(n712), .ZN(n592) );
  NAND2_X1 U706 ( .A1(n593), .A2(n610), .ZN(n594) );
  NOR2_X1 U707 ( .A1(n702), .A2(n595), .ZN(n692) );
  NAND2_X1 U708 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U709 ( .A1(n612), .A2(n599), .ZN(n683) );
  NAND2_X1 U710 ( .A1(n601), .A2(n600), .ZN(n607) );
  NOR2_X1 U711 ( .A1(KEYINPUT87), .A2(n684), .ZN(n603) );
  INV_X1 U712 ( .A(KEYINPUT47), .ZN(n604) );
  NOR2_X1 U713 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U714 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U715 ( .A1(n610), .A2(n702), .ZN(n611) );
  XNOR2_X1 U716 ( .A(KEYINPUT43), .B(n611), .ZN(n613) );
  NAND2_X1 U717 ( .A1(n613), .A2(n612), .ZN(n694) );
  NAND2_X1 U718 ( .A1(n666), .A2(n668), .ZN(n774) );
  NOR2_X1 U719 ( .A1(G898), .A2(n775), .ZN(n761) );
  NAND2_X1 U720 ( .A1(n614), .A2(n761), .ZN(n616) );
  NAND2_X1 U721 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U722 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X1 U723 ( .A(KEYINPUT69), .B(KEYINPUT0), .ZN(n619) );
  NOR2_X1 U724 ( .A1(n786), .A2(KEYINPUT93), .ZN(n624) );
  XNOR2_X1 U725 ( .A(KEYINPUT32), .B(KEYINPUT66), .ZN(n635) );
  NAND2_X1 U726 ( .A1(n441), .A2(n658), .ZN(n626) );
  XNOR2_X1 U727 ( .A(KEYINPUT84), .B(n627), .ZN(n632) );
  XNOR2_X1 U728 ( .A(n633), .B(KEYINPUT83), .ZN(n634) );
  AND2_X1 U729 ( .A1(n636), .A2(n702), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n637), .A2(n660), .ZN(n638) );
  NOR2_X1 U731 ( .A1(n697), .A2(n638), .ZN(n680) );
  NAND2_X1 U732 ( .A1(n639), .A2(n644), .ZN(n640) );
  NAND2_X1 U733 ( .A1(n640), .A2(KEYINPUT44), .ZN(n646) );
  INV_X1 U734 ( .A(KEYINPUT71), .ZN(n641) );
  XNOR2_X1 U735 ( .A(n786), .B(n641), .ZN(n643) );
  INV_X1 U736 ( .A(KEYINPUT44), .ZN(n642) );
  XNOR2_X1 U737 ( .A(n648), .B(KEYINPUT31), .ZN(n690) );
  NOR2_X1 U738 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U739 ( .A(KEYINPUT106), .B(n651), .ZN(n652) );
  NOR2_X1 U740 ( .A1(n690), .A2(n676), .ZN(n654) );
  NOR2_X1 U741 ( .A1(n716), .A2(n654), .ZN(n655) );
  INV_X1 U742 ( .A(n786), .ZN(n656) );
  NAND2_X1 U743 ( .A1(n656), .A2(KEYINPUT44), .ZN(n657) );
  NAND2_X1 U744 ( .A1(n657), .A2(KEYINPUT93), .ZN(n663) );
  AND2_X1 U745 ( .A1(n658), .A2(n697), .ZN(n659) );
  NAND2_X1 U746 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U747 ( .A(KEYINPUT113), .B(n661), .ZN(n788) );
  INV_X1 U748 ( .A(KEYINPUT2), .ZN(n731) );
  AND2_X1 U749 ( .A1(n666), .A2(KEYINPUT2), .ZN(n667) );
  XOR2_X1 U750 ( .A(KEYINPUT94), .B(KEYINPUT85), .Z(n671) );
  XNOR2_X1 U751 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U753 ( .A1(n676), .A2(n687), .ZN(n675) );
  XNOR2_X1 U754 ( .A(n675), .B(G104), .ZN(G6) );
  XOR2_X1 U755 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n678) );
  NAND2_X1 U756 ( .A1(n676), .A2(n689), .ZN(n677) );
  XNOR2_X1 U757 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U758 ( .A(G107), .B(n679), .ZN(G9) );
  XOR2_X1 U759 ( .A(G110), .B(n680), .Z(G12) );
  XOR2_X1 U760 ( .A(G128), .B(KEYINPUT29), .Z(n682) );
  NAND2_X1 U761 ( .A1(n684), .A2(n689), .ZN(n681) );
  XNOR2_X1 U762 ( .A(n682), .B(n681), .ZN(G30) );
  XOR2_X1 U763 ( .A(n683), .B(G143), .Z(G45) );
  NAND2_X1 U764 ( .A1(n684), .A2(n687), .ZN(n685) );
  XNOR2_X1 U765 ( .A(n685), .B(KEYINPUT120), .ZN(n686) );
  XNOR2_X1 U766 ( .A(G146), .B(n686), .ZN(G48) );
  NAND2_X1 U767 ( .A1(n690), .A2(n687), .ZN(n688) );
  XNOR2_X1 U768 ( .A(n688), .B(G113), .ZN(G15) );
  NAND2_X1 U769 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U770 ( .A(n691), .B(G116), .ZN(G18) );
  XNOR2_X1 U771 ( .A(G125), .B(n692), .ZN(n693) );
  XNOR2_X1 U772 ( .A(n693), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U773 ( .A(G140), .B(n694), .ZN(G42) );
  INV_X1 U774 ( .A(n695), .ZN(n710) );
  OR2_X1 U775 ( .A1(n719), .A2(n710), .ZN(n728) );
  NOR2_X1 U776 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U777 ( .A(n698), .B(KEYINPUT49), .ZN(n699) );
  XOR2_X1 U778 ( .A(KEYINPUT121), .B(n700), .Z(n705) );
  NAND2_X1 U779 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U780 ( .A(KEYINPUT50), .B(n703), .Z(n704) );
  NOR2_X1 U781 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U782 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U783 ( .A(KEYINPUT51), .B(n708), .Z(n709) );
  NOR2_X1 U784 ( .A1(n710), .A2(n709), .ZN(n722) );
  NOR2_X1 U785 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U787 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n720) );
  NOR2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U791 ( .A(n723), .B(KEYINPUT122), .Z(n724) );
  XNOR2_X1 U792 ( .A(KEYINPUT52), .B(n724), .ZN(n725) );
  NAND2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U794 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U795 ( .A(n729), .B(KEYINPUT123), .ZN(n730) );
  NAND2_X1 U796 ( .A1(n730), .A2(n775), .ZN(n739) );
  XNOR2_X1 U797 ( .A(KEYINPUT86), .B(n731), .ZN(n733) );
  NAND2_X1 U798 ( .A1(n774), .A2(n733), .ZN(n732) );
  XNOR2_X1 U799 ( .A(n732), .B(KEYINPUT88), .ZN(n735) );
  NAND2_X1 U800 ( .A1(n435), .A2(n733), .ZN(n734) );
  NAND2_X1 U801 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U802 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U803 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U804 ( .A(KEYINPUT53), .B(n740), .ZN(G75) );
  NAND2_X1 U805 ( .A1(n358), .A2(G469), .ZN(n744) );
  XOR2_X1 U806 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n742) );
  NOR2_X1 U807 ( .A1(n756), .A2(n745), .ZN(G54) );
  XNOR2_X1 U808 ( .A(KEYINPUT68), .B(KEYINPUT60), .ZN(n750) );
  NAND2_X1 U809 ( .A1(G478), .A2(n358), .ZN(n751) );
  XNOR2_X1 U810 ( .A(n751), .B(n752), .ZN(n753) );
  NOR2_X1 U811 ( .A1(n756), .A2(n753), .ZN(G63) );
  XNOR2_X1 U812 ( .A(n757), .B(G101), .ZN(n759) );
  XNOR2_X1 U813 ( .A(n759), .B(n758), .ZN(n760) );
  NOR2_X1 U814 ( .A1(n761), .A2(n760), .ZN(n769) );
  NOR2_X1 U815 ( .A1(G953), .A2(n435), .ZN(n763) );
  XOR2_X1 U816 ( .A(KEYINPUT126), .B(n763), .Z(n767) );
  NAND2_X1 U817 ( .A1(G953), .A2(G224), .ZN(n764) );
  XNOR2_X1 U818 ( .A(KEYINPUT61), .B(n764), .ZN(n765) );
  NAND2_X1 U819 ( .A1(n765), .A2(G898), .ZN(n766) );
  NAND2_X1 U820 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U821 ( .A(n769), .B(n768), .ZN(G69) );
  XOR2_X1 U822 ( .A(n770), .B(n771), .Z(n772) );
  XOR2_X1 U823 ( .A(n773), .B(n772), .Z(n777) );
  XNOR2_X1 U824 ( .A(n777), .B(n774), .ZN(n776) );
  NAND2_X1 U825 ( .A1(n776), .A2(n775), .ZN(n782) );
  XNOR2_X1 U826 ( .A(G227), .B(n777), .ZN(n778) );
  NAND2_X1 U827 ( .A1(n778), .A2(G900), .ZN(n779) );
  XOR2_X1 U828 ( .A(KEYINPUT127), .B(n779), .Z(n780) );
  NAND2_X1 U829 ( .A1(G953), .A2(n780), .ZN(n781) );
  NAND2_X1 U830 ( .A1(n782), .A2(n781), .ZN(G72) );
  BUF_X1 U831 ( .A(n783), .Z(n784) );
  XOR2_X1 U832 ( .A(G131), .B(n784), .Z(G33) );
  XOR2_X1 U833 ( .A(G134), .B(n785), .Z(G36) );
  XNOR2_X1 U834 ( .A(n786), .B(G122), .ZN(G24) );
  XOR2_X1 U835 ( .A(n787), .B(G119), .Z(G21) );
  XOR2_X1 U836 ( .A(G101), .B(n788), .Z(G3) );
  XOR2_X1 U837 ( .A(n789), .B(G137), .Z(G39) );
endmodule

