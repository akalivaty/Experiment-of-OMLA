

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813;

  XNOR2_X1 U383 ( .A(n447), .B(n426), .ZN(n602) );
  INV_X1 U384 ( .A(n667), .ZN(n362) );
  XNOR2_X1 U385 ( .A(n617), .B(KEYINPUT1), .ZN(n744) );
  BUF_X1 U386 ( .A(n744), .Z(n418) );
  INV_X1 U387 ( .A(G953), .ZN(n805) );
  NOR2_X2 U388 ( .A1(n599), .A2(n728), .ZN(n603) );
  NOR2_X1 U389 ( .A1(n744), .A2(n745), .ZN(n384) );
  XNOR2_X2 U390 ( .A(n611), .B(KEYINPUT109), .ZN(n728) );
  XNOR2_X2 U391 ( .A(n588), .B(KEYINPUT32), .ZN(n665) );
  OR2_X2 U392 ( .A1(n687), .A2(n442), .ZN(n441) );
  XNOR2_X2 U393 ( .A(n419), .B(n505), .ZN(n687) );
  NOR2_X1 U394 ( .A1(n382), .A2(n467), .ZN(n466) );
  AND2_X1 U395 ( .A1(n784), .A2(n684), .ZN(n415) );
  NOR2_X1 U396 ( .A1(n368), .A2(n401), .ZN(n400) );
  XNOR2_X1 U397 ( .A(n434), .B(n608), .ZN(n732) );
  NOR2_X1 U398 ( .A1(n466), .A2(n464), .ZN(n463) );
  OR2_X1 U399 ( .A1(n658), .A2(KEYINPUT34), .ZN(n467) );
  NOR2_X1 U400 ( .A1(n769), .A2(n382), .ZN(n381) );
  XNOR2_X1 U401 ( .A(n612), .B(KEYINPUT40), .ZN(n386) );
  XNOR2_X1 U402 ( .A(n480), .B(KEYINPUT41), .ZN(n778) );
  NOR2_X1 U403 ( .A1(n474), .A2(n473), .ZN(n627) );
  XNOR2_X1 U404 ( .A(n610), .B(KEYINPUT39), .ZN(n652) );
  XNOR2_X1 U405 ( .A(n384), .B(n385), .ZN(n655) );
  INV_X1 U406 ( .A(n751), .ZN(n361) );
  XNOR2_X1 U407 ( .A(n694), .B(KEYINPUT62), .ZN(n695) );
  XNOR2_X1 U408 ( .A(n796), .B(n562), .ZN(n419) );
  XNOR2_X1 U409 ( .A(n519), .B(KEYINPUT10), .ZN(n803) );
  XNOR2_X1 U410 ( .A(KEYINPUT83), .B(KEYINPUT46), .ZN(n483) );
  BUF_X1 U411 ( .A(n379), .Z(n363) );
  XNOR2_X1 U412 ( .A(n666), .B(KEYINPUT87), .ZN(n676) );
  NOR2_X1 U413 ( .A1(n441), .A2(n440), .ZN(n429) );
  XNOR2_X2 U414 ( .A(n383), .B(n487), .ZN(n802) );
  NOR2_X1 U415 ( .A1(n428), .A2(n429), .ZN(n427) );
  XNOR2_X2 U416 ( .A(G146), .B(G125), .ZN(n519) );
  NAND2_X1 U417 ( .A1(n508), .A2(n684), .ZN(n444) );
  NAND2_X1 U418 ( .A1(n511), .A2(KEYINPUT88), .ZN(n440) );
  INV_X1 U419 ( .A(KEYINPUT15), .ZN(n506) );
  XNOR2_X1 U420 ( .A(n534), .B(n533), .ZN(n638) );
  NOR2_X1 U421 ( .A1(G902), .A2(n699), .ZN(n534) );
  XNOR2_X1 U422 ( .A(G134), .B(G131), .ZN(n561) );
  OR2_X1 U423 ( .A1(n477), .A2(n475), .ZN(n474) );
  XNOR2_X1 U424 ( .A(n670), .B(KEYINPUT81), .ZN(n672) );
  NAND2_X1 U425 ( .A1(n672), .A2(n460), .ZN(n459) );
  NOR2_X1 U426 ( .A1(G237), .A2(G953), .ZN(n527) );
  XNOR2_X1 U427 ( .A(KEYINPUT102), .B(KEYINPUT11), .ZN(n520) );
  XNOR2_X1 U428 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U429 ( .A(G113), .B(G104), .ZN(n522) );
  XOR2_X1 U430 ( .A(G140), .B(G122), .Z(n526) );
  XNOR2_X1 U431 ( .A(n422), .B(G140), .ZN(n578) );
  INV_X1 U432 ( .A(G137), .ZN(n422) );
  OR2_X1 U433 ( .A1(n638), .A2(n637), .ZN(n766) );
  NAND2_X1 U434 ( .A1(n443), .A2(n548), .ZN(n442) );
  INV_X1 U435 ( .A(n508), .ZN(n443) );
  NAND2_X1 U436 ( .A1(n439), .A2(n364), .ZN(n428) );
  INV_X1 U437 ( .A(n440), .ZN(n437) );
  AND2_X1 U438 ( .A1(n602), .A2(n425), .ZN(n615) );
  AND2_X1 U439 ( .A1(n748), .A2(n377), .ZN(n425) );
  OR2_X2 U440 ( .A1(n717), .A2(G902), .ZN(n432) );
  XNOR2_X1 U441 ( .A(n539), .B(G113), .ZN(n491) );
  XNOR2_X1 U442 ( .A(KEYINPUT74), .B(KEYINPUT5), .ZN(n556) );
  XOR2_X1 U443 ( .A(G146), .B(G137), .Z(n557) );
  XNOR2_X1 U444 ( .A(n488), .B(G110), .ZN(n795) );
  XNOR2_X1 U445 ( .A(G104), .B(KEYINPUT91), .ZN(n488) );
  XNOR2_X1 U446 ( .A(n448), .B(n538), .ZN(n567) );
  XNOR2_X1 U447 ( .A(n537), .B(n449), .ZN(n448) );
  INV_X1 U448 ( .A(KEYINPUT66), .ZN(n449) );
  INV_X1 U449 ( .A(KEYINPUT79), .ZN(n498) );
  XNOR2_X1 U450 ( .A(n795), .B(KEYINPUT70), .ZN(n579) );
  XNOR2_X1 U451 ( .A(n472), .B(n471), .ZN(n470) );
  XNOR2_X1 U452 ( .A(G101), .B(G107), .ZN(n471) );
  NAND2_X1 U453 ( .A1(n805), .A2(G227), .ZN(n472) );
  XNOR2_X1 U454 ( .A(KEYINPUT77), .B(G146), .ZN(n469) );
  NAND2_X1 U455 ( .A1(n391), .A2(n635), .ZN(n610) );
  AND2_X1 U456 ( .A1(n634), .A2(n392), .ZN(n391) );
  NOR2_X1 U457 ( .A1(n763), .A2(n393), .ZN(n392) );
  NAND2_X1 U458 ( .A1(n465), .A2(n468), .ZN(n464) );
  XNOR2_X1 U459 ( .A(n424), .B(n423), .ZN(n722) );
  INV_X1 U460 ( .A(KEYINPUT78), .ZN(n423) );
  NAND2_X1 U461 ( .A1(n627), .A2(n626), .ZN(n424) );
  OR2_X1 U462 ( .A1(n672), .A2(n460), .ZN(n457) );
  INV_X1 U463 ( .A(n459), .ZN(n458) );
  NAND2_X1 U464 ( .A1(n665), .A2(n664), .ZN(n666) );
  INV_X1 U465 ( .A(KEYINPUT108), .ZN(n416) );
  XNOR2_X1 U466 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n500) );
  XNOR2_X1 U467 ( .A(n452), .B(KEYINPUT38), .ZN(n763) );
  INV_X1 U468 ( .A(n377), .ZN(n393) );
  INV_X1 U469 ( .A(KEYINPUT73), .ZN(n385) );
  INV_X1 U470 ( .A(n616), .ZN(n478) );
  NAND2_X1 U471 ( .A1(n479), .A2(n476), .ZN(n475) );
  NAND2_X1 U472 ( .A1(n361), .A2(n616), .ZN(n476) );
  XNOR2_X1 U473 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n497) );
  XNOR2_X1 U474 ( .A(G128), .B(KEYINPUT82), .ZN(n568) );
  XOR2_X1 U475 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n569) );
  XNOR2_X1 U476 ( .A(n803), .B(n420), .ZN(n572) );
  XNOR2_X1 U477 ( .A(n578), .B(n421), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n530), .B(n529), .ZN(n699) );
  XNOR2_X1 U479 ( .A(n366), .B(n528), .ZN(n529) );
  XNOR2_X1 U480 ( .A(n524), .B(n523), .ZN(n530) );
  NAND2_X1 U481 ( .A1(n683), .A2(n682), .ZN(n446) );
  NAND2_X1 U482 ( .A1(n427), .A2(n430), .ZN(n620) );
  XNOR2_X1 U483 ( .A(n394), .B(n378), .ZN(n585) );
  XNOR2_X1 U484 ( .A(n390), .B(KEYINPUT30), .ZN(n635) );
  NOR2_X1 U485 ( .A1(n361), .A2(n762), .ZN(n390) );
  INV_X1 U486 ( .A(G478), .ZN(n544) );
  XNOR2_X1 U487 ( .A(n576), .B(n577), .ZN(n426) );
  OR2_X1 U488 ( .A1(n706), .A2(G902), .ZN(n447) );
  XNOR2_X1 U489 ( .A(n591), .B(n590), .ZN(n634) );
  XNOR2_X1 U490 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U491 ( .A(n560), .B(KEYINPUT98), .ZN(n387) );
  XNOR2_X1 U492 ( .A(n542), .B(n451), .ZN(n710) );
  XNOR2_X1 U493 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U494 ( .A(n699), .B(KEYINPUT59), .ZN(n700) );
  XNOR2_X1 U495 ( .A(n802), .B(n485), .ZN(n717) );
  XNOR2_X1 U496 ( .A(n470), .B(n469), .ZN(n486) );
  XNOR2_X1 U497 ( .A(n618), .B(KEYINPUT42), .ZN(n380) );
  INV_X1 U498 ( .A(n722), .ZN(n729) );
  OR2_X1 U499 ( .A1(n511), .A2(KEYINPUT88), .ZN(n364) );
  AND2_X1 U500 ( .A1(n373), .A2(n740), .ZN(n365) );
  XOR2_X1 U501 ( .A(n526), .B(n525), .Z(n366) );
  XNOR2_X1 U502 ( .A(n506), .B(G902), .ZN(n684) );
  AND2_X1 U503 ( .A1(n445), .A2(n444), .ZN(n367) );
  NOR2_X1 U504 ( .A1(n732), .A2(n459), .ZN(n368) );
  XOR2_X1 U505 ( .A(KEYINPUT68), .B(G469), .Z(n369) );
  AND2_X1 U506 ( .A1(KEYINPUT2), .A2(n738), .ZN(n370) );
  AND2_X1 U507 ( .A1(n599), .A2(n587), .ZN(n371) );
  AND2_X1 U508 ( .A1(n813), .A2(n663), .ZN(n372) );
  AND2_X1 U509 ( .A1(n651), .A2(n650), .ZN(n373) );
  NOR2_X1 U510 ( .A1(n766), .A2(n554), .ZN(n374) );
  AND2_X1 U511 ( .A1(n496), .A2(n482), .ZN(n375) );
  AND2_X1 U512 ( .A1(n751), .A2(n478), .ZN(n376) );
  AND2_X1 U513 ( .A1(n601), .A2(n600), .ZN(n377) );
  INV_X1 U514 ( .A(G110), .ZN(n421) );
  INV_X1 U515 ( .A(G116), .ZN(n539) );
  XOR2_X1 U516 ( .A(n555), .B(KEYINPUT22), .Z(n378) );
  INV_X1 U517 ( .A(KEYINPUT0), .ZN(n494) );
  XNOR2_X2 U518 ( .A(n379), .B(n495), .ZN(n796) );
  XNOR2_X1 U519 ( .A(n363), .B(n558), .ZN(n388) );
  XNOR2_X2 U520 ( .A(n492), .B(n491), .ZN(n379) );
  NAND2_X1 U521 ( .A1(n380), .A2(n386), .ZN(n484) );
  XNOR2_X1 U522 ( .A(n380), .B(G137), .ZN(G39) );
  NOR2_X1 U523 ( .A1(n763), .A2(n762), .ZN(n613) );
  NAND2_X1 U524 ( .A1(n367), .A2(n441), .ZN(n452) );
  NAND2_X1 U525 ( .A1(n382), .A2(KEYINPUT34), .ZN(n462) );
  NOR2_X1 U526 ( .A1(n779), .A2(n382), .ZN(n780) );
  XNOR2_X2 U527 ( .A(n657), .B(n656), .ZN(n382) );
  XNOR2_X1 U528 ( .A(n389), .B(n383), .ZN(n694) );
  XNOR2_X2 U529 ( .A(n562), .B(n561), .ZN(n383) );
  XNOR2_X2 U530 ( .A(n432), .B(n369), .ZN(n617) );
  XNOR2_X1 U531 ( .A(n386), .B(G131), .ZN(G33) );
  NAND2_X1 U532 ( .A1(n395), .A2(n374), .ZN(n394) );
  XNOR2_X1 U533 ( .A(n396), .B(KEYINPUT0), .ZN(n395) );
  NOR2_X2 U534 ( .A1(n624), .A2(n518), .ZN(n396) );
  INV_X1 U535 ( .A(n397), .ZN(n410) );
  XNOR2_X2 U536 ( .A(G119), .B(KEYINPUT3), .ZN(n397) );
  NAND2_X1 U537 ( .A1(n397), .A2(n405), .ZN(n412) );
  NAND2_X1 U538 ( .A1(n400), .A2(n398), .ZN(n674) );
  NAND2_X1 U539 ( .A1(n732), .A2(n399), .ZN(n398) );
  AND2_X1 U540 ( .A1(n671), .A2(KEYINPUT106), .ZN(n399) );
  NAND2_X1 U541 ( .A1(n402), .A2(n457), .ZN(n401) );
  NAND2_X1 U542 ( .A1(n403), .A2(n458), .ZN(n402) );
  INV_X1 U543 ( .A(n671), .ZN(n403) );
  NOR2_X2 U544 ( .A1(n658), .A2(n592), .ZN(n593) );
  XNOR2_X2 U545 ( .A(n404), .B(n494), .ZN(n658) );
  NOR2_X1 U546 ( .A1(n624), .A2(n518), .ZN(n404) );
  XNOR2_X2 U547 ( .A(G122), .B(G107), .ZN(n535) );
  XNOR2_X1 U548 ( .A(G101), .B(KEYINPUT69), .ZN(n405) );
  XNOR2_X1 U549 ( .A(G101), .B(KEYINPUT69), .ZN(n493) );
  XNOR2_X1 U550 ( .A(n417), .B(n416), .ZN(n456) );
  XNOR2_X1 U551 ( .A(n484), .B(n483), .ZN(n482) );
  BUF_X1 U552 ( .A(n585), .Z(n406) );
  XNOR2_X1 U553 ( .A(n680), .B(KEYINPUT45), .ZN(n407) );
  BUF_X1 U554 ( .A(n796), .Z(n408) );
  XNOR2_X1 U555 ( .A(n680), .B(KEYINPUT45), .ZN(n739) );
  BUF_X1 U556 ( .A(n620), .Z(n409) );
  INV_X1 U557 ( .A(n617), .ZN(n479) );
  NAND2_X1 U558 ( .A1(n410), .A2(n411), .ZN(n413) );
  NAND2_X1 U559 ( .A1(n413), .A2(n412), .ZN(n492) );
  INV_X1 U560 ( .A(n493), .ZN(n411) );
  AND2_X1 U561 ( .A1(n441), .A2(n512), .ZN(n431) );
  BUF_X1 U562 ( .A(n665), .Z(n414) );
  INV_X1 U563 ( .A(n658), .ZN(n435) );
  BUF_X1 U564 ( .A(n705), .Z(n714) );
  NAND2_X1 U565 ( .A1(n445), .A2(n444), .ZN(n438) );
  NAND2_X1 U566 ( .A1(n674), .A2(n673), .ZN(n417) );
  INV_X1 U567 ( .A(n754), .ZN(n436) );
  XNOR2_X2 U568 ( .A(n620), .B(KEYINPUT19), .ZN(n624) );
  NAND2_X1 U569 ( .A1(n367), .A2(n431), .ZN(n430) );
  XNOR2_X2 U570 ( .A(n433), .B(KEYINPUT4), .ZN(n562) );
  XNOR2_X1 U571 ( .A(n433), .B(n543), .ZN(n451) );
  XNOR2_X2 U572 ( .A(n499), .B(n498), .ZN(n433) );
  NAND2_X1 U573 ( .A1(n436), .A2(n435), .ZN(n434) );
  NAND2_X1 U574 ( .A1(n438), .A2(n437), .ZN(n439) );
  NAND2_X1 U575 ( .A1(n687), .A2(n508), .ZN(n445) );
  AND2_X2 U576 ( .A1(n415), .A2(n446), .ZN(n705) );
  XNOR2_X1 U577 ( .A(n450), .B(n637), .ZN(n670) );
  INV_X1 U578 ( .A(n628), .ZN(n450) );
  NAND2_X1 U579 ( .A1(n585), .A2(n371), .ZN(n588) );
  XNOR2_X2 U580 ( .A(n453), .B(KEYINPUT85), .ZN(n454) );
  NAND2_X1 U581 ( .A1(n455), .A2(n456), .ZN(n453) );
  NAND2_X2 U582 ( .A1(n454), .A2(n679), .ZN(n680) );
  NAND2_X1 U583 ( .A1(n668), .A2(n669), .ZN(n455) );
  INV_X1 U584 ( .A(KEYINPUT106), .ZN(n460) );
  XNOR2_X2 U585 ( .A(n593), .B(n461), .ZN(n671) );
  INV_X1 U586 ( .A(KEYINPUT100), .ZN(n461) );
  NAND2_X1 U587 ( .A1(n463), .A2(n462), .ZN(n661) );
  NAND2_X1 U588 ( .A1(n658), .A2(KEYINPUT34), .ZN(n465) );
  INV_X1 U589 ( .A(n659), .ZN(n468) );
  XNOR2_X1 U590 ( .A(n486), .B(n580), .ZN(n485) );
  NAND2_X1 U591 ( .A1(n759), .A2(n614), .ZN(n480) );
  XNOR2_X1 U592 ( .A(n613), .B(KEYINPUT112), .ZN(n759) );
  NOR2_X1 U593 ( .A1(n615), .A2(n478), .ZN(n473) );
  AND2_X1 U594 ( .A1(n615), .A2(n376), .ZN(n477) );
  NAND2_X1 U595 ( .A1(n778), .A2(n627), .ZN(n618) );
  AND2_X2 U596 ( .A1(n651), .A2(n481), .ZN(n804) );
  AND2_X1 U597 ( .A1(n650), .A2(n738), .ZN(n481) );
  INV_X1 U598 ( .A(n578), .ZN(n487) );
  NAND2_X1 U599 ( .A1(n489), .A2(KEYINPUT64), .ZN(n668) );
  NAND2_X1 U600 ( .A1(n490), .A2(KEYINPUT44), .ZN(n489) );
  NAND2_X1 U601 ( .A1(n676), .A2(n813), .ZN(n490) );
  NAND2_X1 U602 ( .A1(n739), .A2(n365), .ZN(n784) );
  BUF_X1 U603 ( .A(n407), .Z(n789) );
  INV_X1 U604 ( .A(n579), .ZN(n580) );
  XOR2_X1 U605 ( .A(n535), .B(n497), .Z(n495) );
  XOR2_X1 U606 ( .A(KEYINPUT84), .B(n735), .Z(n496) );
  XNOR2_X1 U607 ( .A(KEYINPUT48), .B(KEYINPUT67), .ZN(n648) );
  XNOR2_X1 U608 ( .A(n539), .B(KEYINPUT7), .ZN(n540) );
  INV_X1 U609 ( .A(KEYINPUT2), .ZN(n682) );
  XNOR2_X1 U610 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT104), .B(n638), .Z(n628) );
  XNOR2_X2 U613 ( .A(G143), .B(G128), .ZN(n499) );
  XNOR2_X1 U614 ( .A(n519), .B(n500), .ZN(n503) );
  NAND2_X1 U615 ( .A1(n805), .A2(G224), .ZN(n501) );
  XNOR2_X1 U616 ( .A(n501), .B(KEYINPUT92), .ZN(n502) );
  XNOR2_X1 U617 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U618 ( .A(n579), .B(n504), .ZN(n505) );
  INV_X1 U619 ( .A(G902), .ZN(n563) );
  INV_X1 U620 ( .A(G237), .ZN(n507) );
  NAND2_X1 U621 ( .A1(n563), .A2(n507), .ZN(n509) );
  AND2_X1 U622 ( .A1(n509), .A2(G210), .ZN(n508) );
  NAND2_X1 U623 ( .A1(n509), .A2(G214), .ZN(n510) );
  XNOR2_X1 U624 ( .A(n510), .B(KEYINPUT93), .ZN(n762) );
  INV_X1 U625 ( .A(n762), .ZN(n511) );
  INV_X1 U626 ( .A(KEYINPUT88), .ZN(n512) );
  NAND2_X1 U627 ( .A1(G234), .A2(G237), .ZN(n513) );
  XNOR2_X1 U628 ( .A(n513), .B(KEYINPUT14), .ZN(n773) );
  NOR2_X1 U629 ( .A1(G953), .A2(G952), .ZN(n515) );
  NOR2_X1 U630 ( .A1(G902), .A2(n805), .ZN(n514) );
  NOR2_X1 U631 ( .A1(n515), .A2(n514), .ZN(n516) );
  AND2_X1 U632 ( .A1(n773), .A2(n516), .ZN(n601) );
  NAND2_X1 U633 ( .A1(G953), .A2(G898), .ZN(n517) );
  NAND2_X1 U634 ( .A1(n601), .A2(n517), .ZN(n518) );
  XNOR2_X1 U635 ( .A(n803), .B(n520), .ZN(n524) );
  INV_X1 U636 ( .A(KEYINPUT12), .ZN(n521) );
  XNOR2_X1 U637 ( .A(G143), .B(G131), .ZN(n525) );
  XNOR2_X1 U638 ( .A(n527), .B(KEYINPUT76), .ZN(n559) );
  NAND2_X1 U639 ( .A1(G214), .A2(n559), .ZN(n528) );
  XNOR2_X1 U640 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n532) );
  INV_X1 U641 ( .A(G475), .ZN(n531) );
  XOR2_X1 U642 ( .A(G134), .B(KEYINPUT9), .Z(n536) );
  XNOR2_X1 U643 ( .A(n536), .B(n535), .ZN(n543) );
  XOR2_X1 U644 ( .A(KEYINPUT8), .B(KEYINPUT65), .Z(n538) );
  NAND2_X1 U645 ( .A1(G234), .A2(n805), .ZN(n537) );
  NAND2_X1 U646 ( .A1(n567), .A2(G217), .ZN(n541) );
  NOR2_X1 U647 ( .A1(n710), .A2(G902), .ZN(n545) );
  INV_X1 U648 ( .A(KEYINPUT105), .ZN(n546) );
  XNOR2_X1 U649 ( .A(n547), .B(n546), .ZN(n637) );
  XOR2_X1 U650 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n550) );
  INV_X1 U651 ( .A(n684), .ZN(n548) );
  NAND2_X1 U652 ( .A1(G234), .A2(n548), .ZN(n549) );
  XNOR2_X1 U653 ( .A(n550), .B(n549), .ZN(n575) );
  NAND2_X1 U654 ( .A1(G221), .A2(n575), .ZN(n553) );
  INV_X1 U655 ( .A(KEYINPUT96), .ZN(n551) );
  XNOR2_X1 U656 ( .A(n551), .B(KEYINPUT21), .ZN(n552) );
  XNOR2_X1 U657 ( .A(n553), .B(n552), .ZN(n748) );
  INV_X1 U658 ( .A(n748), .ZN(n554) );
  INV_X1 U659 ( .A(KEYINPUT71), .ZN(n555) );
  XNOR2_X1 U660 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U661 ( .A1(n559), .A2(G210), .ZN(n560) );
  NAND2_X1 U662 ( .A1(n694), .A2(n563), .ZN(n566) );
  INV_X1 U663 ( .A(KEYINPUT99), .ZN(n564) );
  XNOR2_X1 U664 ( .A(n564), .B(G472), .ZN(n565) );
  XNOR2_X2 U665 ( .A(n566), .B(n565), .ZN(n751) );
  XNOR2_X1 U666 ( .A(n751), .B(KEYINPUT6), .ZN(n599) );
  INV_X1 U667 ( .A(n599), .ZN(n654) );
  AND2_X1 U668 ( .A1(n567), .A2(G221), .ZN(n574) );
  XNOR2_X1 U669 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U670 ( .A(n570), .B(G119), .ZN(n571) );
  XNOR2_X1 U671 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U672 ( .A(n574), .B(n573), .ZN(n706) );
  NAND2_X1 U673 ( .A1(G217), .A2(n575), .ZN(n576) );
  XNOR2_X1 U674 ( .A(KEYINPUT94), .B(KEYINPUT25), .ZN(n577) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT107), .ZN(n747) );
  NAND2_X1 U676 ( .A1(n747), .A2(n418), .ZN(n581) );
  NOR2_X1 U677 ( .A1(n654), .A2(n581), .ZN(n582) );
  NAND2_X1 U678 ( .A1(n406), .A2(n582), .ZN(n673) );
  XNOR2_X1 U679 ( .A(n673), .B(G101), .ZN(G3) );
  NAND2_X1 U680 ( .A1(n602), .A2(n418), .ZN(n583) );
  NOR2_X1 U681 ( .A1(n751), .A2(n583), .ZN(n584) );
  NAND2_X1 U682 ( .A1(n406), .A2(n584), .ZN(n664) );
  XNOR2_X1 U683 ( .A(G110), .B(KEYINPUT114), .ZN(n586) );
  XNOR2_X1 U684 ( .A(n664), .B(n586), .ZN(G12) );
  NOR2_X1 U685 ( .A1(n747), .A2(n418), .ZN(n587) );
  XNOR2_X1 U686 ( .A(n414), .B(G119), .ZN(G21) );
  INV_X1 U687 ( .A(KEYINPUT97), .ZN(n591) );
  INV_X1 U688 ( .A(n602), .ZN(n589) );
  NAND2_X1 U689 ( .A1(n589), .A2(n748), .ZN(n745) );
  NOR2_X1 U690 ( .A1(n745), .A2(n617), .ZN(n590) );
  NAND2_X1 U691 ( .A1(n634), .A2(n361), .ZN(n592) );
  AND2_X1 U692 ( .A1(n628), .A2(n637), .ZN(n723) );
  INV_X1 U693 ( .A(n723), .ZN(n731) );
  NOR2_X1 U694 ( .A1(n671), .A2(n731), .ZN(n597) );
  XOR2_X1 U695 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n595) );
  XNOR2_X1 U696 ( .A(G107), .B(KEYINPUT26), .ZN(n594) );
  XNOR2_X1 U697 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U698 ( .A(n597), .B(n596), .ZN(G9) );
  NOR2_X1 U699 ( .A1(n628), .A2(n637), .ZN(n611) );
  NOR2_X1 U700 ( .A1(n728), .A2(n671), .ZN(n598) );
  XOR2_X1 U701 ( .A(G104), .B(n598), .Z(G6) );
  NAND2_X1 U702 ( .A1(G953), .A2(G900), .ZN(n600) );
  NAND2_X1 U703 ( .A1(n603), .A2(n615), .ZN(n619) );
  NOR2_X1 U704 ( .A1(n762), .A2(n619), .ZN(n604) );
  XNOR2_X1 U705 ( .A(n604), .B(KEYINPUT110), .ZN(n605) );
  NAND2_X1 U706 ( .A1(n605), .A2(n418), .ZN(n606) );
  XNOR2_X1 U707 ( .A(n606), .B(KEYINPUT43), .ZN(n607) );
  INV_X1 U708 ( .A(n452), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n607), .A2(n639), .ZN(n650) );
  XNOR2_X1 U710 ( .A(n650), .B(G140), .ZN(G42) );
  NAND2_X1 U711 ( .A1(n655), .A2(n751), .ZN(n754) );
  XNOR2_X1 U712 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n608) );
  NOR2_X1 U713 ( .A1(n728), .A2(n732), .ZN(n609) );
  XOR2_X1 U714 ( .A(G113), .B(n609), .Z(G15) );
  NAND2_X1 U715 ( .A1(n652), .A2(n611), .ZN(n612) );
  INV_X1 U716 ( .A(n766), .ZN(n614) );
  XOR2_X1 U717 ( .A(KEYINPUT28), .B(KEYINPUT111), .Z(n616) );
  INV_X1 U718 ( .A(n619), .ZN(n621) );
  NAND2_X1 U719 ( .A1(n621), .A2(n409), .ZN(n622) );
  XNOR2_X1 U720 ( .A(n622), .B(KEYINPUT36), .ZN(n623) );
  NOR2_X2 U721 ( .A1(n418), .A2(n623), .ZN(n735) );
  INV_X1 U722 ( .A(KEYINPUT47), .ZN(n631) );
  BUF_X1 U723 ( .A(n624), .Z(n625) );
  INV_X1 U724 ( .A(n625), .ZN(n626) );
  NOR2_X1 U725 ( .A1(KEYINPUT81), .A2(n670), .ZN(n629) );
  NAND2_X1 U726 ( .A1(n722), .A2(n629), .ZN(n630) );
  NAND2_X1 U727 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U728 ( .A1(n722), .A2(KEYINPUT47), .ZN(n632) );
  NAND2_X1 U729 ( .A1(n633), .A2(n632), .ZN(n642) );
  AND2_X1 U730 ( .A1(n635), .A2(n634), .ZN(n636) );
  AND2_X1 U731 ( .A1(n377), .A2(n636), .ZN(n641) );
  NAND2_X1 U732 ( .A1(n638), .A2(n637), .ZN(n659) );
  NOR2_X1 U733 ( .A1(n659), .A2(n639), .ZN(n640) );
  NAND2_X1 U734 ( .A1(n641), .A2(n640), .ZN(n727) );
  NAND2_X1 U735 ( .A1(n642), .A2(n727), .ZN(n646) );
  AND2_X1 U736 ( .A1(n722), .A2(KEYINPUT81), .ZN(n643) );
  NOR2_X1 U737 ( .A1(KEYINPUT47), .A2(n643), .ZN(n644) );
  INV_X1 U738 ( .A(n670), .ZN(n760) );
  NOR2_X1 U739 ( .A1(n644), .A2(n760), .ZN(n645) );
  NOR2_X1 U740 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U741 ( .A1(n375), .A2(n647), .ZN(n649) );
  XNOR2_X1 U742 ( .A(n649), .B(n648), .ZN(n651) );
  NAND2_X1 U743 ( .A1(n723), .A2(n652), .ZN(n738) );
  INV_X1 U744 ( .A(KEYINPUT75), .ZN(n653) );
  XNOR2_X1 U745 ( .A(n804), .B(n653), .ZN(n681) );
  NAND2_X1 U746 ( .A1(n655), .A2(n654), .ZN(n657) );
  XOR2_X1 U747 ( .A(KEYINPUT90), .B(KEYINPUT33), .Z(n656) );
  INV_X1 U748 ( .A(KEYINPUT35), .ZN(n660) );
  XNOR2_X2 U749 ( .A(n661), .B(n660), .ZN(n813) );
  INV_X1 U750 ( .A(KEYINPUT44), .ZN(n662) );
  NOR2_X1 U751 ( .A1(n662), .A2(KEYINPUT64), .ZN(n663) );
  INV_X1 U752 ( .A(n676), .ZN(n667) );
  NAND2_X1 U753 ( .A1(n372), .A2(n667), .ZN(n669) );
  INV_X1 U754 ( .A(n813), .ZN(n675) );
  NOR2_X1 U755 ( .A1(n675), .A2(KEYINPUT44), .ZN(n678) );
  XNOR2_X1 U756 ( .A(n362), .B(KEYINPUT86), .ZN(n677) );
  NAND2_X1 U757 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U758 ( .A1(n681), .A2(n407), .ZN(n683) );
  XNOR2_X1 U759 ( .A(KEYINPUT80), .B(n370), .ZN(n740) );
  NAND2_X1 U760 ( .A1(n705), .A2(G210), .ZN(n689) );
  XNOR2_X1 U761 ( .A(KEYINPUT89), .B(KEYINPUT54), .ZN(n685) );
  XOR2_X1 U762 ( .A(n685), .B(KEYINPUT55), .Z(n686) );
  XNOR2_X1 U763 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U764 ( .A(n689), .B(n688), .ZN(n691) );
  INV_X1 U765 ( .A(G952), .ZN(n690) );
  NAND2_X1 U766 ( .A1(n690), .A2(G953), .ZN(n708) );
  NAND2_X1 U767 ( .A1(n691), .A2(n708), .ZN(n693) );
  INV_X1 U768 ( .A(KEYINPUT56), .ZN(n692) );
  XNOR2_X1 U769 ( .A(n693), .B(n692), .ZN(G51) );
  NAND2_X1 U770 ( .A1(n705), .A2(G472), .ZN(n696) );
  XNOR2_X1 U771 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U772 ( .A1(n697), .A2(n708), .ZN(n698) );
  XNOR2_X1 U773 ( .A(n698), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U774 ( .A1(n705), .A2(G475), .ZN(n701) );
  XNOR2_X1 U775 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U776 ( .A1(n702), .A2(n708), .ZN(n704) );
  INV_X1 U777 ( .A(KEYINPUT60), .ZN(n703) );
  XNOR2_X1 U778 ( .A(n704), .B(n703), .ZN(G60) );
  NAND2_X1 U779 ( .A1(n714), .A2(G217), .ZN(n707) );
  XNOR2_X1 U780 ( .A(n707), .B(n706), .ZN(n709) );
  INV_X1 U781 ( .A(n708), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n709), .A2(n720), .ZN(G66) );
  NAND2_X1 U783 ( .A1(n714), .A2(G478), .ZN(n712) );
  XNOR2_X1 U784 ( .A(n710), .B(KEYINPUT124), .ZN(n711) );
  XNOR2_X1 U785 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U786 ( .A1(n713), .A2(n720), .ZN(G63) );
  NAND2_X1 U787 ( .A1(n714), .A2(G469), .ZN(n719) );
  XNOR2_X1 U788 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n715) );
  XNOR2_X1 U789 ( .A(n715), .B(KEYINPUT58), .ZN(n716) );
  XNOR2_X1 U790 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U791 ( .A(n719), .B(n718), .ZN(n721) );
  NOR2_X1 U792 ( .A1(n721), .A2(n720), .ZN(G54) );
  XOR2_X1 U793 ( .A(G128), .B(KEYINPUT29), .Z(n725) );
  NAND2_X1 U794 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U795 ( .A(n725), .B(n724), .ZN(G30) );
  XOR2_X1 U796 ( .A(G143), .B(KEYINPUT115), .Z(n726) );
  XNOR2_X1 U797 ( .A(n727), .B(n726), .ZN(G45) );
  NOR2_X1 U798 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U799 ( .A(G146), .B(n730), .Z(G48) );
  NOR2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U801 ( .A(KEYINPUT116), .B(n733), .Z(n734) );
  XNOR2_X1 U802 ( .A(G116), .B(n734), .ZN(G18) );
  XOR2_X1 U803 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n737) );
  XNOR2_X1 U804 ( .A(G125), .B(n735), .ZN(n736) );
  XNOR2_X1 U805 ( .A(n737), .B(n736), .ZN(G27) );
  XNOR2_X1 U806 ( .A(G134), .B(n738), .ZN(G36) );
  INV_X1 U807 ( .A(n789), .ZN(n743) );
  INV_X1 U808 ( .A(n740), .ZN(n741) );
  NAND2_X1 U809 ( .A1(n804), .A2(n741), .ZN(n742) );
  OR2_X1 U810 ( .A1(n743), .A2(n742), .ZN(n783) );
  NAND2_X1 U811 ( .A1(n745), .A2(n418), .ZN(n746) );
  XNOR2_X1 U812 ( .A(n746), .B(KEYINPUT50), .ZN(n753) );
  NOR2_X1 U813 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U814 ( .A(KEYINPUT49), .B(n749), .Z(n750) );
  NOR2_X1 U815 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U816 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U817 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U818 ( .A(KEYINPUT51), .B(n756), .Z(n757) );
  NAND2_X1 U819 ( .A1(n778), .A2(n757), .ZN(n758) );
  XOR2_X1 U820 ( .A(KEYINPUT118), .B(n758), .Z(n771) );
  NAND2_X1 U821 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U822 ( .A(KEYINPUT120), .B(n761), .Z(n768) );
  NAND2_X1 U823 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U824 ( .A(KEYINPUT119), .B(n764), .ZN(n765) );
  NOR2_X1 U825 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U826 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U827 ( .A(KEYINPUT121), .B(n381), .Z(n770) );
  NOR2_X1 U828 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U829 ( .A(KEYINPUT52), .B(n772), .ZN(n775) );
  NAND2_X1 U830 ( .A1(G952), .A2(n773), .ZN(n774) );
  NOR2_X1 U831 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U832 ( .A(KEYINPUT122), .B(n776), .Z(n777) );
  NAND2_X1 U833 ( .A1(n805), .A2(n777), .ZN(n781) );
  INV_X1 U834 ( .A(n778), .ZN(n779) );
  NOR2_X1 U835 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U836 ( .A1(n783), .A2(n782), .ZN(n787) );
  INV_X1 U837 ( .A(n784), .ZN(n785) );
  NOR2_X1 U838 ( .A1(n785), .A2(n682), .ZN(n786) );
  OR2_X1 U839 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U840 ( .A(KEYINPUT53), .B(n788), .Z(G75) );
  NAND2_X1 U841 ( .A1(n789), .A2(n805), .ZN(n793) );
  NAND2_X1 U842 ( .A1(G953), .A2(G224), .ZN(n790) );
  XNOR2_X1 U843 ( .A(KEYINPUT61), .B(n790), .ZN(n791) );
  NAND2_X1 U844 ( .A1(n791), .A2(G898), .ZN(n792) );
  NAND2_X1 U845 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U846 ( .A(n794), .B(KEYINPUT126), .ZN(n801) );
  XNOR2_X1 U847 ( .A(n408), .B(n795), .ZN(n798) );
  NOR2_X1 U848 ( .A1(G898), .A2(n805), .ZN(n797) );
  NOR2_X1 U849 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U850 ( .A(n799), .B(KEYINPUT125), .Z(n800) );
  XNOR2_X1 U851 ( .A(n801), .B(n800), .ZN(G69) );
  XNOR2_X1 U852 ( .A(n802), .B(n803), .ZN(n807) );
  XNOR2_X1 U853 ( .A(n807), .B(n804), .ZN(n806) );
  NAND2_X1 U854 ( .A1(n806), .A2(n805), .ZN(n812) );
  XNOR2_X1 U855 ( .A(n807), .B(G227), .ZN(n808) );
  XNOR2_X1 U856 ( .A(n808), .B(KEYINPUT127), .ZN(n809) );
  NAND2_X1 U857 ( .A1(n809), .A2(G900), .ZN(n810) );
  NAND2_X1 U858 ( .A1(n810), .A2(G953), .ZN(n811) );
  NAND2_X1 U859 ( .A1(n812), .A2(n811), .ZN(G72) );
  XNOR2_X1 U860 ( .A(n813), .B(G122), .ZN(G24) );
endmodule

