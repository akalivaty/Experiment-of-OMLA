//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT74), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT74), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n189), .A3(G104), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT75), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n196), .A2(new_n189), .A3(KEYINPUT75), .A4(G104), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n192), .A2(new_n195), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n189), .A2(G104), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  INV_X1    g017(.A(new_n202), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(new_n190), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n201), .A2(new_n203), .B1(G101), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G116), .ZN(new_n208));
  OAI21_X1  g022(.A(G113), .B1(new_n208), .B2(KEYINPUT5), .ZN(new_n209));
  XNOR2_X1  g023(.A(G116), .B(G119), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(KEYINPUT5), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n210), .A3(KEYINPUT67), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n211), .A2(new_n212), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n210), .A2(KEYINPUT5), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT79), .B1(new_n226), .B2(new_n209), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n206), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G101), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(new_n201), .B2(new_n204), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n195), .A2(new_n192), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n199), .A2(new_n200), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n203), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n224), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT67), .B1(new_n223), .B2(new_n210), .ZN(new_n237));
  OAI22_X1  g051(.A1(new_n236), .A2(new_n237), .B1(new_n210), .B2(new_n223), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n232), .A3(new_n204), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n229), .A2(KEYINPUT4), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n228), .B1(new_n235), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G110), .B(G122), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT80), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n228), .B(new_n244), .C1(new_n235), .C2(new_n242), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT6), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(KEYINPUT6), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n238), .B(new_n241), .C1(new_n230), .C2(new_n234), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n244), .B1(new_n251), .B2(new_n228), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n243), .A2(new_n254), .A3(new_n245), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT80), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n249), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT0), .A4(G128), .ZN(new_n262));
  XNOR2_X1  g076(.A(G143), .B(G146), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT0), .B(G128), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G125), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n259), .A2(new_n261), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT66), .B(G128), .Z(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(G143), .B2(new_n258), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n259), .A3(new_n261), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n266), .B1(new_n275), .B2(G125), .ZN(new_n276));
  INV_X1    g090(.A(G224), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n277), .A2(G953), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n257), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G210), .B1(G237), .B2(G902), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(KEYINPUT7), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n276), .B(new_n284), .Z(new_n285));
  NAND2_X1  g099(.A1(new_n205), .A2(G101), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n233), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n225), .A2(new_n287), .A3(new_n227), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n210), .A2(KEYINPUT5), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n209), .B1(new_n289), .B2(KEYINPUT81), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(KEYINPUT81), .B2(new_n289), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n237), .B2(new_n236), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n206), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n244), .B(KEYINPUT8), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n285), .B1(new_n288), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n248), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n283), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n281), .A2(new_n282), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n282), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT80), .B(new_n255), .C1(new_n250), .C2(new_n252), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n279), .B1(new_n302), .B2(new_n249), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n303), .B2(new_n298), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n188), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n265), .B1(new_n239), .B2(new_n240), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n230), .B2(new_n234), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT64), .B1(new_n308), .B2(G137), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n309), .A2(KEYINPUT11), .B1(new_n308), .B2(G137), .ZN(new_n310));
  INV_X1    g124(.A(G131), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT11), .ZN(new_n312));
  OAI211_X1 g126(.A(KEYINPUT64), .B(new_n312), .C1(new_n308), .C2(G137), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n311), .B1(new_n310), .B2(new_n313), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n274), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n267), .B1(new_n270), .B2(new_n272), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n263), .A2(KEYINPUT76), .A3(new_n273), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n233), .A3(new_n286), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT10), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n271), .B2(new_n274), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n206), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n307), .A2(new_n316), .A3(new_n324), .A4(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT68), .B(G953), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G227), .ZN(new_n330));
  XOR2_X1   g144(.A(G110), .B(G140), .Z(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n328), .A2(KEYINPUT78), .A3(new_n333), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n307), .A2(new_n324), .A3(new_n327), .ZN(new_n338));
  INV_X1    g152(.A(new_n316), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT12), .ZN(new_n342));
  INV_X1    g156(.A(new_n275), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n287), .A2(new_n343), .ZN(new_n344));
  AOI211_X1 g158(.A(new_n342), .B(new_n316), .C1(new_n344), .C2(new_n322), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n322), .B1(new_n206), .B2(new_n275), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT12), .B1(new_n346), .B2(new_n339), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n328), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n332), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n341), .A2(G469), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G469), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n348), .A2(new_n334), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n333), .B1(new_n340), .B2(new_n328), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n352), .B(new_n283), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n352), .A2(new_n283), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n351), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT9), .B(G234), .ZN(new_n359));
  OAI21_X1  g173(.A(G221), .B1(new_n359), .B2(G902), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G237), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n329), .A2(G214), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n260), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n329), .A2(G143), .A3(G214), .A4(new_n362), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n311), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT17), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n311), .A3(new_n365), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G140), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G125), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(KEYINPUT16), .ZN(new_n373));
  XNOR2_X1  g187(.A(G125), .B(G140), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(KEYINPUT16), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(G146), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n258), .B(new_n373), .C1(KEYINPUT16), .C2(new_n374), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n366), .A2(new_n379), .A3(KEYINPUT17), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n366), .B2(KEYINPUT17), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n370), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT83), .B1(new_n374), .B2(new_n258), .ZN(new_n383));
  INV_X1    g197(.A(G125), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n372), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G146), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n383), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT18), .A3(G131), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n364), .B2(new_n365), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n364), .A2(new_n365), .A3(new_n390), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n382), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n193), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT86), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n382), .A2(KEYINPUT86), .A3(new_n398), .A4(new_n394), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n283), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G475), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n374), .B(KEYINPUT19), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n377), .B1(new_n258), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n369), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n366), .B2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n394), .A2(new_n408), .A3(new_n398), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n395), .B2(new_n397), .ZN(new_n410));
  NOR2_X1   g224(.A1(G475), .A2(G902), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT85), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n404), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n398), .B1(new_n382), .B2(new_n394), .ZN(new_n415));
  NOR4_X1   g229(.A1(new_n415), .A2(new_n409), .A3(KEYINPUT20), .A4(new_n412), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n403), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G217), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n359), .A2(new_n418), .A3(G953), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(KEYINPUT89), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n260), .A2(G128), .ZN(new_n424));
  OR2_X1    g238(.A1(KEYINPUT66), .A2(G128), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT66), .A2(G128), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(G143), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT87), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n427), .A2(KEYINPUT87), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n308), .B(new_n424), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G116), .B(G122), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(new_n189), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n268), .A2(new_n435), .A3(G143), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n428), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT13), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n424), .B(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT88), .A3(G134), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n439), .B1(new_n436), .B2(new_n428), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(new_n308), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n434), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n214), .A2(G122), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n189), .B1(new_n447), .B2(KEYINPUT14), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n432), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n308), .B1(new_n437), .B2(new_n424), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n452), .B2(new_n431), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n422), .B(new_n423), .C1(new_n446), .C2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n431), .A2(new_n433), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT88), .B1(new_n441), .B2(G134), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n444), .A2(new_n443), .A3(new_n308), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n431), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n449), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n458), .A2(new_n460), .A3(new_n421), .A4(new_n420), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n461), .A3(new_n283), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT15), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n463), .A3(G478), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(G478), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n454), .A2(new_n461), .A3(new_n283), .A4(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n283), .B(new_n329), .C1(G234), .C2(G237), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(G898), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G952), .ZN(new_n470));
  AOI211_X1 g284(.A(G953), .B(new_n470), .C1(G234), .C2(G237), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n464), .A2(new_n466), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n417), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n305), .A2(new_n361), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n418), .B1(G234), .B2(new_n283), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT23), .B1(new_n272), .B2(G119), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n272), .A2(G119), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n425), .A2(KEYINPUT23), .A3(G119), .A4(new_n426), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G110), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT24), .B(G110), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n481), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n425), .A2(new_n426), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n487), .B(new_n488), .C1(new_n207), .C2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n485), .B(new_n490), .C1(new_n376), .C2(new_n377), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n488), .B1(new_n489), .B2(new_n207), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n486), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(G110), .B2(new_n484), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n386), .A2(G146), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n375), .B2(G146), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT22), .B(G137), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n329), .A2(G221), .A3(G234), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n498), .B(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT25), .B1(new_n504), .B2(new_n283), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT73), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n479), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n498), .A2(new_n503), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n498), .A2(new_n503), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n508), .B1(new_n511), .B2(G902), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n504), .A2(KEYINPUT25), .A3(new_n283), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT73), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n478), .A2(G902), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n507), .A2(new_n514), .B1(new_n504), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(G472), .A2(G902), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n265), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n314), .B2(new_n315), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n308), .A2(G137), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n308), .A2(G137), .ZN(new_n525));
  OAI21_X1  g339(.A(G131), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n275), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n521), .A2(new_n527), .A3(KEYINPUT30), .ZN(new_n528));
  INV_X1    g342(.A(new_n527), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n521), .A2(KEYINPUT65), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n309), .A2(KEYINPUT11), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n313), .A3(new_n523), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G131), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n265), .B1(new_n533), .B2(new_n522), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT65), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n529), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n528), .B(new_n238), .C1(new_n537), .C2(KEYINPUT30), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n218), .A2(new_n224), .B1(new_n216), .B2(new_n217), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n521), .A2(new_n527), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n329), .A2(G210), .A3(new_n362), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT27), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(G101), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n538), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n538), .A2(KEYINPUT31), .A3(new_n540), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT28), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n540), .A2(KEYINPUT69), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT69), .B1(new_n540), .B2(new_n550), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n540), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n534), .A2(new_n535), .ZN(new_n555));
  AOI211_X1 g369(.A(KEYINPUT65), .B(new_n265), .C1(new_n533), .C2(new_n522), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n527), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n554), .B1(new_n557), .B2(new_n238), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n553), .B1(new_n558), .B2(new_n550), .ZN(new_n559));
  INV_X1    g373(.A(new_n544), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n519), .B1(new_n549), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n538), .A2(new_n540), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n560), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT29), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n553), .B(new_n544), .C1(new_n558), .C2(new_n550), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n521), .A2(new_n527), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n238), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(KEYINPUT71), .A3(new_n540), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT71), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n571), .A3(new_n238), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(KEYINPUT28), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n560), .A2(new_n565), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n553), .A3(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n575), .A2(new_n283), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n562), .A2(KEYINPUT32), .B1(new_n577), .B2(G472), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n579));
  AOI22_X1  g393(.A1(new_n547), .A2(new_n548), .B1(new_n559), .B2(new_n560), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n519), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n517), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n477), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(new_n301), .C1(new_n303), .C2(new_n298), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n586), .A2(new_n187), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n300), .A2(KEYINPUT90), .A3(new_n304), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n587), .A2(new_n473), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G472), .B1(new_n580), .B2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n549), .A2(new_n561), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n518), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n516), .A2(new_n360), .A3(new_n358), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n394), .A2(new_n408), .A3(new_n398), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n392), .A2(new_n393), .ZN(new_n597));
  INV_X1    g411(.A(new_n378), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n407), .A2(new_n366), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n599), .B2(new_n368), .ZN(new_n600));
  INV_X1    g414(.A(new_n381), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n366), .A2(new_n379), .A3(KEYINPUT17), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n597), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n596), .B(new_n413), .C1(new_n604), .C2(new_n398), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT20), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n410), .A2(new_n404), .A3(new_n413), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n606), .A2(new_n607), .B1(new_n402), .B2(G475), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n454), .A2(new_n461), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT91), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT91), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n454), .A2(new_n461), .A3(new_n612), .A4(new_n609), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT92), .B1(new_n446), .B2(new_n453), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n615), .A2(new_n419), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n609), .B1(new_n615), .B2(new_n419), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n614), .A2(G478), .A3(new_n283), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT93), .B(G478), .Z(new_n620));
  NAND2_X1  g434(.A1(new_n462), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n608), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n589), .A2(new_n595), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT94), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  NAND2_X1  g440(.A1(new_n587), .A2(new_n588), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n606), .A2(new_n607), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT95), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n464), .A2(new_n466), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n473), .B(KEYINPUT96), .Z(new_n635));
  NAND2_X1  g449(.A1(new_n403), .A2(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n627), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n595), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  INV_X1    g454(.A(KEYINPUT36), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n503), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n498), .ZN(new_n643));
  INV_X1    g457(.A(new_n515), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n507), .B2(new_n514), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n305), .A2(new_n361), .A3(new_n475), .A4(new_n647), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n648), .A2(new_n593), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  AOI21_X1  g465(.A(new_n646), .B1(new_n578), .B2(new_n581), .ZN(new_n652));
  INV_X1    g466(.A(new_n627), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n464), .A2(new_n466), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n467), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT97), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(KEYINPUT97), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n657), .A2(new_n472), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n403), .A2(new_n660), .ZN(new_n661));
  AOI211_X1 g475(.A(new_n654), .B(new_n661), .C1(new_n630), .C2(new_n631), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n652), .A2(new_n653), .A3(new_n361), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  NAND3_X1  g478(.A1(new_n591), .A2(KEYINPUT32), .A3(new_n518), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n570), .A2(new_n572), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n283), .B1(new_n666), .B2(new_n544), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n560), .B1(new_n538), .B2(new_n540), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n665), .A2(new_n581), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n659), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n361), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n300), .A2(new_n304), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT38), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n608), .A2(new_n654), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n678), .A2(new_n187), .A3(new_n646), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n672), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n260), .ZN(G45));
  NAND2_X1  g496(.A1(new_n283), .A2(G478), .ZN(new_n683));
  AOI221_X4 g497(.A(new_n683), .B1(new_n616), .B2(new_n617), .C1(new_n611), .C2(new_n613), .ZN(new_n684));
  INV_X1    g498(.A(new_n621), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n417), .B(new_n660), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n652), .A2(new_n653), .A3(new_n687), .A4(new_n361), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NAND2_X1  g503(.A1(new_n577), .A2(G472), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n665), .A2(new_n581), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n352), .A2(KEYINPUT99), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n340), .A2(new_n328), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n332), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n333), .B(new_n328), .C1(new_n345), .C2(new_n347), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n693), .B1(new_n697), .B2(new_n283), .ZN(new_n698));
  AOI211_X1 g512(.A(G902), .B(new_n692), .C1(new_n695), .C2(new_n696), .ZN(new_n699));
  INV_X1    g513(.A(new_n360), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n691), .A2(new_n516), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n622), .A2(new_n587), .A3(new_n473), .A4(new_n588), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT41), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n219), .ZN(G15));
  NOR4_X1   g520(.A1(new_n702), .A2(new_n627), .A3(new_n634), .A4(new_n636), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n214), .ZN(G18));
  AND3_X1   g522(.A1(new_n587), .A2(new_n588), .A3(new_n701), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n652), .A2(new_n709), .A3(new_n475), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  AND3_X1   g525(.A1(new_n587), .A2(new_n588), .A3(new_n678), .ZN(new_n712));
  INV_X1    g526(.A(new_n549), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n544), .B1(new_n573), .B2(new_n553), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n518), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n590), .ZN(new_n716));
  INV_X1    g530(.A(new_n635), .ZN(new_n717));
  NOR4_X1   g531(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n712), .A2(new_n516), .A3(new_n716), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT100), .B(G122), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G24));
  NAND2_X1  g535(.A1(new_n686), .A2(KEYINPUT101), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n715), .A2(new_n647), .A3(new_n590), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT101), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n622), .A2(new_n724), .A3(new_n660), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n709), .A2(new_n722), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  NAND3_X1  g541(.A1(new_n300), .A2(new_n187), .A3(new_n304), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT103), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n300), .A2(new_n304), .A3(new_n730), .A4(new_n187), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n358), .A2(new_n360), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n358), .A2(KEYINPUT102), .A3(new_n360), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n729), .A2(new_n731), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n358), .A2(KEYINPUT102), .A3(new_n360), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT102), .B1(new_n358), .B2(new_n360), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(KEYINPUT104), .A3(new_n731), .A4(new_n729), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n722), .A2(new_n725), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT32), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n592), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n578), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n516), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n743), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n691), .A2(new_n516), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n738), .B2(new_n742), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n744), .A2(KEYINPUT42), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n751), .A2(KEYINPUT42), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  NAND3_X1  g570(.A1(new_n743), .A2(new_n582), .A3(new_n662), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NOR2_X1   g572(.A1(new_n684), .A2(new_n685), .ZN(new_n759));
  OR3_X1    g573(.A1(new_n759), .A2(KEYINPUT43), .A3(new_n417), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT43), .B1(new_n759), .B2(new_n417), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n646), .B1(new_n590), .B2(new_n592), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n760), .A2(new_n762), .A3(KEYINPUT44), .A4(new_n761), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n731), .A3(new_n729), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n341), .A2(new_n350), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n341), .A2(KEYINPUT45), .A3(new_n350), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(G469), .A3(new_n771), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT105), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT105), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n356), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n355), .B1(new_n775), .B2(KEYINPUT46), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n360), .B(new_n673), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n767), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(G137), .Z(G39));
  OAI21_X1  g594(.A(new_n360), .B1(new_n776), .B2(new_n777), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT106), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(KEYINPUT47), .ZN(new_n783));
  XNOR2_X1  g597(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n360), .B(new_n785), .C1(new_n776), .C2(new_n777), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n729), .A2(new_n731), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n787), .A2(new_n691), .A3(new_n516), .A4(new_n686), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n783), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n783), .A2(KEYINPUT107), .A3(new_n786), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NAND3_X1  g608(.A1(new_n516), .A2(new_n360), .A3(new_n187), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT108), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n796), .A2(new_n677), .A3(new_n417), .A4(new_n759), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n698), .A2(new_n699), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT109), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT49), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n672), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n760), .A2(new_n471), .A3(new_n761), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n716), .A2(new_n516), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n701), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n677), .A2(new_n187), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT50), .ZN(new_n808));
  INV_X1    g622(.A(new_n802), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n787), .A2(new_n805), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n723), .A3(new_n810), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n787), .A2(new_n517), .A3(new_n472), .A4(new_n805), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n672), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n759), .A2(new_n608), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n808), .A2(new_n816), .A3(KEYINPUT51), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n802), .A2(new_n803), .A3(new_n787), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n799), .A2(new_n700), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT114), .Z(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n783), .B2(new_n786), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n817), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n783), .A2(new_n786), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n819), .B1(new_n824), .B2(new_n820), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n808), .A3(new_n816), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n809), .A2(new_n750), .A3(new_n810), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT48), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n829), .A2(KEYINPUT115), .A3(new_n830), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n470), .B(G953), .C1(new_n804), .C2(new_n709), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n813), .A2(new_n622), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n831), .B(new_n834), .C1(new_n829), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n743), .A2(new_n745), .A3(new_n723), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n646), .A2(new_n661), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n633), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT110), .B1(new_n464), .B2(new_n466), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n841), .A2(new_n845), .A3(new_n361), .A4(new_n632), .ZN(new_n846));
  INV_X1    g660(.A(new_n691), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n787), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n839), .A2(new_n757), .A3(new_n840), .A4(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n753), .B2(new_n662), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n839), .B1(new_n851), .B2(new_n840), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n582), .A2(new_n589), .A3(new_n622), .A4(new_n701), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(new_n649), .A3(new_n719), .A4(new_n583), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT111), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n676), .A2(new_n187), .A3(new_n635), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n608), .B1(new_n843), .B2(new_n844), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n654), .A2(KEYINPUT110), .ZN(new_n861));
  INV_X1    g675(.A(new_n844), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n417), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n305), .A3(KEYINPUT111), .A4(new_n635), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n864), .A3(new_n595), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n595), .A2(new_n305), .A3(new_n622), .A4(new_n635), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n710), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n856), .A2(new_n867), .A3(new_n707), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n663), .A2(new_n688), .A3(new_n726), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n587), .A2(new_n588), .A3(new_n678), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n670), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n361), .A2(KEYINPUT113), .A3(new_n646), .A4(new_n660), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n646), .A2(new_n660), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n732), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT52), .B1(new_n869), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(new_n871), .B2(new_n876), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n663), .A3(new_n688), .A4(new_n726), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n755), .A2(new_n868), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n853), .A2(new_n854), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n743), .A2(new_n582), .A3(new_n754), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n749), .B(new_n744), .C1(new_n738), .C2(new_n742), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT42), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n881), .B(new_n884), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n663), .A2(new_n688), .A3(new_n726), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n877), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n718), .A2(new_n587), .A3(new_n588), .A4(new_n678), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n803), .A2(new_n891), .B1(new_n648), .B2(new_n593), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n752), .A2(new_n476), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n704), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n865), .A2(new_n710), .A3(new_n866), .ZN(new_n895));
  INV_X1    g709(.A(new_n707), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n887), .A2(new_n890), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n757), .A2(new_n840), .A3(new_n849), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT112), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n851), .A2(new_n839), .A3(new_n840), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT53), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n838), .B1(new_n883), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n854), .B1(new_n853), .B2(new_n882), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n898), .A2(new_n902), .A3(KEYINPUT53), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(KEYINPUT54), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n837), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(G952), .A2(G953), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n801), .B1(new_n908), .B2(new_n909), .ZN(G75));
  AOI21_X1  g724(.A(new_n283), .B1(new_n905), .B2(new_n906), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(G210), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n257), .A2(new_n280), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n303), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT55), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n912), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n912), .B2(new_n913), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n329), .A2(G952), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G51));
  XNOR2_X1  g734(.A(new_n356), .B(KEYINPUT57), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n904), .A2(new_n907), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT116), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n904), .A2(KEYINPUT116), .A3(new_n907), .A4(new_n921), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n697), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n773), .A2(new_n774), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n911), .A2(KEYINPUT117), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT117), .B1(new_n911), .B2(new_n928), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n919), .B1(new_n926), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n415), .B2(new_n409), .ZN(new_n934));
  INV_X1    g748(.A(new_n919), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .A4(new_n410), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G60));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT59), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n904), .A2(new_n907), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n614), .A2(new_n618), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n940), .A2(new_n942), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n944), .A3(new_n919), .ZN(G63));
  XNOR2_X1  g759(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n418), .A2(new_n283), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n905), .B2(new_n906), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(new_n504), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n643), .B(KEYINPUT119), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n935), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n951), .A2(new_n953), .A3(KEYINPUT61), .A4(new_n935), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  OAI21_X1  g772(.A(G953), .B1(new_n468), .B2(new_n277), .ZN(new_n959));
  INV_X1    g773(.A(new_n329), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n868), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n302), .B(new_n249), .C1(G898), .C2(new_n329), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT120), .Z(new_n963));
  XNOR2_X1  g777(.A(new_n961), .B(new_n963), .ZN(G69));
  OAI21_X1  g778(.A(new_n528), .B1(new_n537), .B2(KEYINPUT30), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(new_n405), .Z(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT121), .Z(new_n967));
  INV_X1    g781(.A(new_n779), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n863), .A2(new_n622), .ZN(new_n969));
  NOR4_X1   g783(.A1(new_n752), .A2(new_n787), .A3(new_n969), .A4(new_n674), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT122), .Z(new_n971));
  OAI21_X1  g785(.A(KEYINPUT62), .B1(new_n681), .B2(new_n869), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n681), .A2(KEYINPUT62), .A3(new_n869), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(new_n793), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n967), .B1(new_n976), .B2(new_n960), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n960), .A2(G900), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n968), .A2(KEYINPUT123), .A3(new_n889), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT123), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n779), .B2(new_n869), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n755), .A2(new_n757), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n778), .A2(new_n870), .A3(new_n749), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n982), .A2(new_n793), .A3(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n978), .B(new_n966), .C1(new_n986), .C2(new_n960), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n977), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n329), .B1(G227), .B2(G900), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT124), .Z(new_n990));
  XNOR2_X1  g804(.A(new_n988), .B(new_n990), .ZN(G72));
  NOR2_X1   g805(.A1(new_n563), .A2(new_n544), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT125), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n982), .A2(new_n793), .A3(new_n868), .A4(new_n985), .ZN(new_n995));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT63), .Z(new_n997));
  AOI21_X1  g811(.A(new_n994), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT126), .B1(new_n998), .B2(new_n919), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n975), .A2(new_n793), .A3(new_n868), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n997), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n905), .A2(new_n906), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n997), .B1(new_n564), .B2(KEYINPUT127), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n545), .A2(KEYINPUT127), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n564), .B2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g819(.A1(new_n1001), .A2(new_n668), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n998), .A2(KEYINPUT126), .A3(new_n919), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(G57));
endmodule


