

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U550 ( .A1(n694), .A2(n693), .ZN(n729) );
  AND2_X2 U551 ( .A1(n685), .A2(n684), .ZN(n692) );
  NOR2_X1 U552 ( .A1(G164), .A2(G1384), .ZN(n580) );
  NOR2_X1 U553 ( .A1(n683), .A2(n687), .ZN(n515) );
  BUF_X1 U554 ( .A(n614), .Z(n604) );
  XNOR2_X1 U555 ( .A(n591), .B(KEYINPUT31), .ZN(n662) );
  NAND2_X1 U556 ( .A1(G8), .A2(n614), .ZN(n687) );
  XNOR2_X1 U557 ( .A(n580), .B(KEYINPUT64), .ZN(n715) );
  NOR2_X1 U558 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XOR2_X1 U560 ( .A(KEYINPUT1), .B(n531), .Z(n796) );
  XOR2_X2 U561 ( .A(KEYINPUT17), .B(n516), .Z(n886) );
  NAND2_X1 U562 ( .A1(G138), .A2(n886), .ZN(n519) );
  INV_X1 U563 ( .A(G2105), .ZN(n520) );
  NAND2_X1 U564 ( .A1(n520), .A2(G2104), .ZN(n517) );
  XNOR2_X2 U565 ( .A(n517), .B(KEYINPUT65), .ZN(n887) );
  NAND2_X1 U566 ( .A1(G102), .A2(n887), .ZN(n518) );
  NAND2_X1 U567 ( .A1(n519), .A2(n518), .ZN(n525) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n520), .ZN(n882) );
  NAND2_X1 U569 ( .A1(G126), .A2(n882), .ZN(n523) );
  NAND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XOR2_X2 U571 ( .A(KEYINPUT66), .B(n521), .Z(n883) );
  NAND2_X1 U572 ( .A1(G114), .A2(n883), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U574 ( .A1(n525), .A2(n524), .ZN(G164) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n792) );
  NAND2_X1 U576 ( .A1(n792), .A2(G89), .ZN(n526) );
  XNOR2_X1 U577 ( .A(n526), .B(KEYINPUT4), .ZN(n528) );
  XOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .Z(n570) );
  INV_X1 U579 ( .A(G651), .ZN(n530) );
  NOR2_X1 U580 ( .A1(n570), .A2(n530), .ZN(n789) );
  NAND2_X1 U581 ( .A1(G76), .A2(n789), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U583 ( .A(n529), .B(KEYINPUT5), .ZN(n536) );
  NOR2_X2 U584 ( .A1(G651), .A2(n570), .ZN(n788) );
  NAND2_X1 U585 ( .A1(G51), .A2(n788), .ZN(n533) );
  NOR2_X1 U586 ( .A1(G543), .A2(n530), .ZN(n531) );
  NAND2_X1 U587 ( .A1(G63), .A2(n796), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U589 ( .A(KEYINPUT6), .B(n534), .Z(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U591 ( .A(n537), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U592 ( .A1(G137), .A2(n886), .ZN(n539) );
  NAND2_X1 U593 ( .A1(G125), .A2(n882), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n544) );
  NAND2_X1 U595 ( .A1(G101), .A2(n887), .ZN(n540) );
  XOR2_X1 U596 ( .A(KEYINPUT23), .B(n540), .Z(n542) );
  NAND2_X1 U597 ( .A1(G113), .A2(n883), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U599 ( .A1(n544), .A2(n543), .ZN(G160) );
  NAND2_X1 U600 ( .A1(G52), .A2(n788), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G64), .A2(n796), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G90), .A2(n792), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G77), .A2(n789), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  XNOR2_X1 U607 ( .A(KEYINPUT68), .B(n550), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n552), .A2(n551), .ZN(G171) );
  NAND2_X1 U609 ( .A1(G88), .A2(n792), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G75), .A2(n789), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U612 ( .A1(G50), .A2(n788), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G62), .A2(n796), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U615 ( .A1(n558), .A2(n557), .ZN(G166) );
  INV_X1 U616 ( .A(G166), .ZN(G303) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U618 ( .A1(G86), .A2(n792), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G61), .A2(n796), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U621 ( .A(KEYINPUT80), .B(n561), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n789), .A2(G73), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT2), .B(n562), .Z(n563) );
  NOR2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n788), .A2(G48), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(G305) );
  NAND2_X1 U627 ( .A1(G49), .A2(n788), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G74), .A2(G651), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U630 ( .A1(n796), .A2(n569), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n570), .A2(G87), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U633 ( .A1(G85), .A2(n792), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G72), .A2(n789), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G47), .A2(n788), .ZN(n575) );
  XNOR2_X1 U637 ( .A(KEYINPUT67), .B(n575), .ZN(n576) );
  NOR2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n796), .A2(G60), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(G290) );
  NAND2_X1 U641 ( .A1(G160), .A2(G40), .ZN(n716) );
  INV_X1 U642 ( .A(n715), .ZN(n581) );
  NOR2_X2 U643 ( .A1(n716), .A2(n581), .ZN(n586) );
  INV_X1 U644 ( .A(n586), .ZN(n614) );
  NOR2_X1 U645 ( .A1(G1966), .A2(n687), .ZN(n668) );
  NOR2_X1 U646 ( .A1(G2084), .A2(n604), .ZN(n664) );
  NOR2_X1 U647 ( .A1(n668), .A2(n664), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT94), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n583), .A2(G8), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n584), .B(KEYINPUT30), .ZN(n585) );
  NOR2_X1 U651 ( .A1(G168), .A2(n585), .ZN(n590) );
  INV_X1 U652 ( .A(G1961), .ZN(n989) );
  NAND2_X1 U653 ( .A1(n604), .A2(n989), .ZN(n588) );
  BUF_X2 U654 ( .A(n586), .Z(n611) );
  XNOR2_X1 U655 ( .A(G2078), .B(KEYINPUT25), .ZN(n911) );
  NAND2_X1 U656 ( .A1(n611), .A2(n911), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n596) );
  NOR2_X1 U658 ( .A1(G171), .A2(n596), .ZN(n589) );
  OR2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U660 ( .A1(G1971), .A2(n687), .ZN(n593) );
  NOR2_X1 U661 ( .A1(G2090), .A2(n604), .ZN(n592) );
  NOR2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n594), .A2(G303), .ZN(n595) );
  XNOR2_X1 U664 ( .A(n595), .B(KEYINPUT96), .ZN(n655) );
  AND2_X1 U665 ( .A1(n662), .A2(n655), .ZN(n654) );
  NAND2_X1 U666 ( .A1(n596), .A2(G171), .ZN(n653) );
  NAND2_X1 U667 ( .A1(G53), .A2(n788), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G65), .A2(n796), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G91), .A2(n792), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G78), .A2(n789), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n1000) );
  NAND2_X1 U674 ( .A1(n611), .A2(G2072), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT27), .ZN(n606) );
  AND2_X1 U676 ( .A1(G1956), .A2(n604), .ZN(n605) );
  NOR2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n646) );
  NOR2_X1 U678 ( .A1(n1000), .A2(n646), .ZN(n607) );
  XOR2_X1 U679 ( .A(n607), .B(KEYINPUT28), .Z(n650) );
  NAND2_X1 U680 ( .A1(G1348), .A2(n614), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G2067), .A2(n611), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U683 ( .A(KEYINPUT92), .B(n610), .Z(n640) );
  XOR2_X1 U684 ( .A(KEYINPUT26), .B(KEYINPUT90), .Z(n613) );
  NAND2_X1 U685 ( .A1(n611), .A2(G1996), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n613), .B(n612), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G1341), .A2(n614), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(KEYINPUT91), .ZN(n616) );
  NOR2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n642) );
  NAND2_X1 U690 ( .A1(G92), .A2(n792), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G66), .A2(n796), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n624) );
  NAND2_X1 U693 ( .A1(G54), .A2(n788), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G79), .A2(n789), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U696 ( .A(KEYINPUT74), .B(n622), .ZN(n623) );
  NOR2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n625), .B(KEYINPUT15), .ZN(n1008) );
  INV_X1 U699 ( .A(n1008), .ZN(n799) );
  NAND2_X1 U700 ( .A1(n788), .A2(G43), .ZN(n626) );
  XNOR2_X1 U701 ( .A(KEYINPUT71), .B(n626), .ZN(n637) );
  NAND2_X1 U702 ( .A1(n792), .A2(G81), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n627), .B(KEYINPUT12), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G68), .A2(n789), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U706 ( .A(n630), .B(KEYINPUT70), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT13), .ZN(n635) );
  XOR2_X1 U708 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n633) );
  NAND2_X1 U709 ( .A1(G56), .A2(n796), .ZN(n632) );
  XNOR2_X1 U710 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n991) );
  AND2_X1 U713 ( .A1(n799), .A2(n991), .ZN(n638) );
  AND2_X1 U714 ( .A1(n642), .A2(n638), .ZN(n639) );
  NOR2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U716 ( .A(KEYINPUT93), .B(n641), .ZN(n645) );
  NAND2_X1 U717 ( .A1(n991), .A2(n642), .ZN(n643) );
  NAND2_X1 U718 ( .A1(n1008), .A2(n643), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n1000), .A2(n646), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U723 ( .A(KEYINPUT29), .B(n651), .Z(n652) );
  NAND2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n663) );
  NAND2_X1 U725 ( .A1(n654), .A2(n663), .ZN(n658) );
  INV_X1 U726 ( .A(n655), .ZN(n656) );
  OR2_X1 U727 ( .A1(n656), .A2(G286), .ZN(n657) );
  AND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n659), .A2(G8), .ZN(n661) );
  XOR2_X1 U730 ( .A(KEYINPUT32), .B(KEYINPUT97), .Z(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n671) );
  NAND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U733 ( .A1(G8), .A2(n664), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U736 ( .A(KEYINPUT95), .B(n669), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n682) );
  NOR2_X1 U738 ( .A1(G2090), .A2(G303), .ZN(n672) );
  NAND2_X1 U739 ( .A1(G8), .A2(n672), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n682), .A2(n673), .ZN(n674) );
  AND2_X1 U741 ( .A1(n674), .A2(n687), .ZN(n678) );
  NOR2_X1 U742 ( .A1(G1981), .A2(G305), .ZN(n675) );
  XOR2_X1 U743 ( .A(n675), .B(KEYINPUT24), .Z(n676) );
  NOR2_X1 U744 ( .A1(n687), .A2(n676), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n694) );
  NOR2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n686) );
  NOR2_X1 U747 ( .A1(G1971), .A2(G303), .ZN(n679) );
  NOR2_X1 U748 ( .A1(n686), .A2(n679), .ZN(n996) );
  INV_X1 U749 ( .A(KEYINPUT33), .ZN(n680) );
  AND2_X1 U750 ( .A1(n996), .A2(n680), .ZN(n681) );
  NAND2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n995) );
  INV_X1 U753 ( .A(n995), .ZN(n683) );
  OR2_X1 U754 ( .A1(KEYINPUT33), .A2(n515), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n686), .A2(KEYINPUT33), .ZN(n688) );
  NOR2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n690) );
  XOR2_X1 U757 ( .A(G1981), .B(G305), .Z(n1011) );
  INV_X1 U758 ( .A(n1011), .ZN(n689) );
  NOR2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U761 ( .A1(G129), .A2(n882), .ZN(n696) );
  NAND2_X1 U762 ( .A1(G117), .A2(n883), .ZN(n695) );
  NAND2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n697), .B(KEYINPUT87), .ZN(n699) );
  NAND2_X1 U765 ( .A1(G141), .A2(n886), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U767 ( .A1(n887), .A2(G105), .ZN(n700) );
  XOR2_X1 U768 ( .A(KEYINPUT38), .B(n700), .Z(n701) );
  NOR2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U770 ( .A(KEYINPUT88), .B(n703), .Z(n876) );
  NAND2_X1 U771 ( .A1(G1996), .A2(n876), .ZN(n713) );
  NAND2_X1 U772 ( .A1(n883), .A2(G107), .ZN(n704) );
  XNOR2_X1 U773 ( .A(n704), .B(KEYINPUT86), .ZN(n711) );
  NAND2_X1 U774 ( .A1(G131), .A2(n886), .ZN(n706) );
  NAND2_X1 U775 ( .A1(G95), .A2(n887), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U777 ( .A1(G119), .A2(n882), .ZN(n707) );
  XNOR2_X1 U778 ( .A(KEYINPUT85), .B(n707), .ZN(n708) );
  NOR2_X1 U779 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n893) );
  NAND2_X1 U781 ( .A1(G1991), .A2(n893), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U783 ( .A(KEYINPUT89), .B(n714), .ZN(n978) );
  INV_X1 U784 ( .A(n978), .ZN(n717) );
  NOR2_X1 U785 ( .A1(n716), .A2(n715), .ZN(n746) );
  NAND2_X1 U786 ( .A1(n717), .A2(n746), .ZN(n733) );
  NAND2_X1 U787 ( .A1(G140), .A2(n886), .ZN(n719) );
  NAND2_X1 U788 ( .A1(G104), .A2(n887), .ZN(n718) );
  NAND2_X1 U789 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U790 ( .A(KEYINPUT34), .B(n720), .ZN(n725) );
  NAND2_X1 U791 ( .A1(G128), .A2(n882), .ZN(n722) );
  NAND2_X1 U792 ( .A1(G116), .A2(n883), .ZN(n721) );
  NAND2_X1 U793 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U794 ( .A(n723), .B(KEYINPUT35), .Z(n724) );
  NOR2_X1 U795 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U796 ( .A(KEYINPUT36), .B(n726), .Z(n727) );
  XOR2_X1 U797 ( .A(KEYINPUT84), .B(n727), .Z(n877) );
  XNOR2_X1 U798 ( .A(G2067), .B(KEYINPUT37), .ZN(n744) );
  NOR2_X1 U799 ( .A1(n877), .A2(n744), .ZN(n972) );
  NAND2_X1 U800 ( .A1(n746), .A2(n972), .ZN(n742) );
  NAND2_X1 U801 ( .A1(n733), .A2(n742), .ZN(n728) );
  XNOR2_X1 U802 ( .A(n730), .B(KEYINPUT98), .ZN(n732) );
  XNOR2_X1 U803 ( .A(G1986), .B(G290), .ZN(n1004) );
  NAND2_X1 U804 ( .A1(n1004), .A2(n746), .ZN(n731) );
  NAND2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n749) );
  XOR2_X1 U806 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n741) );
  NOR2_X1 U807 ( .A1(G1996), .A2(n876), .ZN(n960) );
  INV_X1 U808 ( .A(n733), .ZN(n737) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n735) );
  NOR2_X1 U810 ( .A1(G1991), .A2(n893), .ZN(n734) );
  XOR2_X1 U811 ( .A(KEYINPUT99), .B(n734), .Z(n976) );
  NOR2_X1 U812 ( .A1(n735), .A2(n976), .ZN(n736) );
  NOR2_X1 U813 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U814 ( .A(n738), .B(KEYINPUT100), .ZN(n739) );
  NOR2_X1 U815 ( .A1(n960), .A2(n739), .ZN(n740) );
  XNOR2_X1 U816 ( .A(n741), .B(n740), .ZN(n743) );
  NAND2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n877), .A2(n744), .ZN(n973) );
  NAND2_X1 U819 ( .A1(n745), .A2(n973), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n751) );
  XNOR2_X1 U822 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n750) );
  XNOR2_X1 U823 ( .A(n751), .B(n750), .ZN(G329) );
  XNOR2_X1 U824 ( .A(G2451), .B(G2443), .ZN(n761) );
  XOR2_X1 U825 ( .A(G2446), .B(KEYINPUT103), .Z(n753) );
  XNOR2_X1 U826 ( .A(KEYINPUT104), .B(G2438), .ZN(n752) );
  XNOR2_X1 U827 ( .A(n753), .B(n752), .ZN(n757) );
  XOR2_X1 U828 ( .A(G2435), .B(G2454), .Z(n755) );
  XNOR2_X1 U829 ( .A(G1341), .B(G1348), .ZN(n754) );
  XNOR2_X1 U830 ( .A(n755), .B(n754), .ZN(n756) );
  XOR2_X1 U831 ( .A(n757), .B(n756), .Z(n759) );
  XNOR2_X1 U832 ( .A(G2430), .B(G2427), .ZN(n758) );
  XNOR2_X1 U833 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n761), .B(n760), .ZN(n762) );
  AND2_X1 U835 ( .A1(n762), .A2(G14), .ZN(G401) );
  AND2_X1 U836 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U837 ( .A(G860), .B(KEYINPUT72), .Z(n769) );
  INV_X1 U838 ( .A(n991), .ZN(n800) );
  OR2_X1 U839 ( .A1(n769), .A2(n800), .ZN(G153) );
  INV_X1 U840 ( .A(G57), .ZN(G237) );
  NAND2_X1 U841 ( .A1(G7), .A2(G661), .ZN(n763) );
  XNOR2_X1 U842 ( .A(n763), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U843 ( .A(G223), .ZN(n829) );
  NAND2_X1 U844 ( .A1(n829), .A2(G567), .ZN(n764) );
  XOR2_X1 U845 ( .A(KEYINPUT11), .B(n764), .Z(G234) );
  XNOR2_X1 U846 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U847 ( .A1(G868), .A2(G301), .ZN(n766) );
  INV_X1 U848 ( .A(G868), .ZN(n812) );
  NAND2_X1 U849 ( .A1(n1008), .A2(n812), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n766), .A2(n765), .ZN(G284) );
  INV_X1 U851 ( .A(n1000), .ZN(G299) );
  NOR2_X1 U852 ( .A1(G868), .A2(G299), .ZN(n768) );
  NOR2_X1 U853 ( .A1(G286), .A2(n812), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n768), .A2(n767), .ZN(G297) );
  NAND2_X1 U855 ( .A1(G559), .A2(n769), .ZN(n770) );
  XOR2_X1 U856 ( .A(KEYINPUT75), .B(n770), .Z(n771) );
  NAND2_X1 U857 ( .A1(n771), .A2(n799), .ZN(n772) );
  XNOR2_X1 U858 ( .A(n772), .B(KEYINPUT16), .ZN(n773) );
  XNOR2_X1 U859 ( .A(KEYINPUT76), .B(n773), .ZN(G148) );
  NAND2_X1 U860 ( .A1(n799), .A2(G868), .ZN(n774) );
  NOR2_X1 U861 ( .A1(G559), .A2(n774), .ZN(n776) );
  NOR2_X1 U862 ( .A1(G868), .A2(n800), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n776), .A2(n775), .ZN(G282) );
  NAND2_X1 U864 ( .A1(G123), .A2(n882), .ZN(n777) );
  XOR2_X1 U865 ( .A(KEYINPUT18), .B(n777), .Z(n782) );
  NAND2_X1 U866 ( .A1(n887), .A2(G99), .ZN(n779) );
  NAND2_X1 U867 ( .A1(G111), .A2(n883), .ZN(n778) );
  NAND2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U869 ( .A(KEYINPUT77), .B(n780), .Z(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n886), .A2(G135), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n969) );
  XOR2_X1 U873 ( .A(G2096), .B(KEYINPUT78), .Z(n785) );
  XNOR2_X1 U874 ( .A(n969), .B(n785), .ZN(n787) );
  INV_X1 U875 ( .A(G2100), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(G156) );
  NAND2_X1 U877 ( .A1(G55), .A2(n788), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G80), .A2(n789), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U880 ( .A1(G93), .A2(n792), .ZN(n793) );
  XNOR2_X1 U881 ( .A(KEYINPUT79), .B(n793), .ZN(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U883 ( .A1(n796), .A2(G67), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n813) );
  NAND2_X1 U885 ( .A1(G559), .A2(n799), .ZN(n801) );
  XNOR2_X1 U886 ( .A(n801), .B(n800), .ZN(n810) );
  NOR2_X1 U887 ( .A1(G860), .A2(n810), .ZN(n802) );
  XOR2_X1 U888 ( .A(n813), .B(n802), .Z(G145) );
  XNOR2_X1 U889 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n804) );
  XNOR2_X1 U890 ( .A(G288), .B(KEYINPUT19), .ZN(n803) );
  XNOR2_X1 U891 ( .A(n804), .B(n803), .ZN(n805) );
  XNOR2_X1 U892 ( .A(G305), .B(n805), .ZN(n807) );
  XNOR2_X1 U893 ( .A(n1000), .B(G166), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n807), .B(n806), .ZN(n808) );
  XNOR2_X1 U895 ( .A(n808), .B(G290), .ZN(n809) );
  XNOR2_X1 U896 ( .A(n809), .B(n813), .ZN(n901) );
  XNOR2_X1 U897 ( .A(n901), .B(n810), .ZN(n811) );
  NOR2_X1 U898 ( .A1(n812), .A2(n811), .ZN(n815) );
  NOR2_X1 U899 ( .A1(G868), .A2(n813), .ZN(n814) );
  NOR2_X1 U900 ( .A1(n815), .A2(n814), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n816) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n816), .Z(n817) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U907 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n821) );
  NAND2_X1 U908 ( .A1(G132), .A2(G82), .ZN(n820) );
  XNOR2_X1 U909 ( .A(n821), .B(n820), .ZN(n822) );
  NOR2_X1 U910 ( .A1(n822), .A2(G218), .ZN(n823) );
  NAND2_X1 U911 ( .A1(G96), .A2(n823), .ZN(n834) );
  NAND2_X1 U912 ( .A1(n834), .A2(G2106), .ZN(n827) );
  NAND2_X1 U913 ( .A1(G69), .A2(G120), .ZN(n824) );
  NOR2_X1 U914 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(G108), .A2(n825), .ZN(n835) );
  NAND2_X1 U916 ( .A1(n835), .A2(G567), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(n836) );
  NAND2_X1 U918 ( .A1(G483), .A2(G661), .ZN(n828) );
  NOR2_X1 U919 ( .A1(n836), .A2(n828), .ZN(n833) );
  NAND2_X1 U920 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n829), .ZN(G217) );
  NAND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n830) );
  XNOR2_X1 U923 ( .A(KEYINPUT105), .B(n830), .ZN(n831) );
  NAND2_X1 U924 ( .A1(n831), .A2(G661), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G82), .ZN(G220) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n836), .ZN(G319) );
  XOR2_X1 U936 ( .A(G2096), .B(G2678), .Z(n838) );
  XNOR2_X1 U937 ( .A(G2067), .B(KEYINPUT43), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U939 ( .A(n839), .B(KEYINPUT42), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2072), .B(G2090), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U942 ( .A(KEYINPUT106), .B(G2100), .Z(n843) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1961), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n848), .B(G2474), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1981), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U952 ( .A(KEYINPUT41), .B(G1956), .Z(n852) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G124), .A2(n882), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n855), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U958 ( .A1(n887), .A2(G100), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G112), .A2(n883), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U961 ( .A(KEYINPUT108), .B(n858), .Z(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G136), .A2(n886), .ZN(n861) );
  XNOR2_X1 U964 ( .A(KEYINPUT107), .B(n861), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(G162) );
  XNOR2_X1 U966 ( .A(G162), .B(n969), .ZN(n881) );
  XOR2_X1 U967 ( .A(KEYINPUT110), .B(KEYINPUT48), .Z(n872) );
  NAND2_X1 U968 ( .A1(G139), .A2(n886), .ZN(n865) );
  NAND2_X1 U969 ( .A1(G103), .A2(n887), .ZN(n864) );
  NAND2_X1 U970 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G127), .A2(n882), .ZN(n867) );
  NAND2_X1 U972 ( .A1(G115), .A2(n883), .ZN(n866) );
  NAND2_X1 U973 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n963) );
  XNOR2_X1 U976 ( .A(n963), .B(KEYINPUT109), .ZN(n871) );
  XNOR2_X1 U977 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U978 ( .A(n873), .B(KEYINPUT46), .Z(n875) );
  XNOR2_X1 U979 ( .A(G164), .B(KEYINPUT111), .ZN(n874) );
  XNOR2_X1 U980 ( .A(n875), .B(n874), .ZN(n879) );
  XOR2_X1 U981 ( .A(n877), .B(n876), .Z(n878) );
  XNOR2_X1 U982 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n881), .B(n880), .ZN(n897) );
  NAND2_X1 U984 ( .A1(G130), .A2(n882), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G118), .A2(n883), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n892) );
  NAND2_X1 U987 ( .A1(G142), .A2(n886), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G106), .A2(n887), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U990 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U993 ( .A(G160), .B(n895), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U995 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U996 ( .A(KEYINPUT112), .B(n991), .Z(n900) );
  XNOR2_X1 U997 ( .A(G286), .B(G171), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n1008), .B(n901), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n904), .ZN(G397) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n905), .B(KEYINPUT49), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G401), .A2(n906), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n907), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT113), .B(n908), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1011 ( .A(G1991), .B(G25), .ZN(n920) );
  XNOR2_X1 U1012 ( .A(G27), .B(n911), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(G2067), .B(G26), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(G33), .B(G2072), .ZN(n912) );
  NOR2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G32), .B(G1996), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(KEYINPUT117), .B(n918), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(G28), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n922), .B(KEYINPUT53), .ZN(n925) );
  XOR2_X1 U1023 ( .A(G2084), .B(G34), .Z(n923) );
  XNOR2_X1 U1024 ( .A(KEYINPUT54), .B(n923), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(G35), .B(G2090), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(KEYINPUT55), .B(n928), .ZN(n930) );
  INV_X1 U1029 ( .A(G29), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1031 ( .A1(n931), .A2(G11), .ZN(n988) );
  XNOR2_X1 U1032 ( .A(G1971), .B(G22), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(G23), .B(G1976), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n935) );
  XOR2_X1 U1035 ( .A(G1986), .B(G24), .Z(n934) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n937) );
  XOR2_X1 U1037 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n936) );
  XNOR2_X1 U1038 ( .A(n937), .B(n936), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(G1961), .B(G5), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n938) );
  NOR2_X1 U1041 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G1956), .B(G20), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n942) );
  NOR2_X1 U1046 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1047 ( .A(KEYINPUT123), .B(n944), .ZN(n945) );
  NOR2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1049 ( .A(KEYINPUT124), .B(n947), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(G1348), .B(KEYINPUT59), .ZN(n948) );
  XNOR2_X1 U1051 ( .A(n948), .B(G4), .ZN(n949) );
  NAND2_X1 U1052 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1053 ( .A(n951), .B(KEYINPUT60), .ZN(n952) );
  XOR2_X1 U1054 ( .A(KEYINPUT125), .B(n952), .Z(n953) );
  NOR2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1056 ( .A(KEYINPUT61), .B(n955), .Z(n956) );
  NOR2_X1 U1057 ( .A1(G16), .A2(n956), .ZN(n957) );
  XNOR2_X1 U1058 ( .A(KEYINPUT127), .B(n957), .ZN(n986) );
  XOR2_X1 U1059 ( .A(G2090), .B(G162), .Z(n958) );
  XNOR2_X1 U1060 ( .A(KEYINPUT114), .B(n958), .ZN(n959) );
  NOR2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n962) );
  XOR2_X1 U1062 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n961) );
  XOR2_X1 U1063 ( .A(n962), .B(n961), .Z(n968) );
  XOR2_X1 U1064 ( .A(G2072), .B(n963), .Z(n965) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n964) );
  NOR2_X1 U1066 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1067 ( .A(KEYINPUT50), .B(n966), .ZN(n967) );
  NAND2_X1 U1068 ( .A1(n968), .A2(n967), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G160), .B(G2084), .ZN(n970) );
  NAND2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1076 ( .A(KEYINPUT52), .B(n981), .Z(n982) );
  NOR2_X1 U1077 ( .A1(KEYINPUT55), .A2(n982), .ZN(n983) );
  XOR2_X1 U1078 ( .A(KEYINPUT116), .B(n983), .Z(n984) );
  NAND2_X1 U1079 ( .A1(n984), .A2(G29), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n1021) );
  XNOR2_X1 U1082 ( .A(KEYINPUT56), .B(G16), .ZN(n1019) );
  XNOR2_X1 U1083 ( .A(G171), .B(KEYINPUT120), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(n990), .B(n989), .ZN(n993) );
  XOR2_X1 U1085 ( .A(n991), .B(G1341), .Z(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n1007) );
  INV_X1 U1087 ( .A(G1971), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(G166), .A2(n994), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1091 ( .A(KEYINPUT121), .B(n999), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(n1000), .B(G1956), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1005), .B(KEYINPUT122), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G1348), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(G168), .B(G1966), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(n1013), .B(KEYINPUT57), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n1014) );
  XNOR2_X1 U1103 ( .A(n1015), .B(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

