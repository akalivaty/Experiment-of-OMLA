//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n558, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n466), .A2(KEYINPUT64), .B1(G113), .B2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n469), .A3(G125), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n461), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n462), .A2(KEYINPUT65), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT66), .A2(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(G2104), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n475), .A2(new_n479), .A3(G137), .A4(new_n461), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n472), .B2(new_n474), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n471), .A2(new_n483), .ZN(G160));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n475), .A2(new_n479), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(new_n461), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n475), .A2(new_n479), .A3(KEYINPUT67), .A4(G2105), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT68), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT69), .Z(new_n494));
  NOR2_X1   g069(.A1(new_n486), .A2(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(G136), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n491), .A2(new_n496), .ZN(G162));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n475), .A2(new_n479), .A3(new_n499), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n500), .A2(KEYINPUT4), .B1(new_n468), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n475), .A2(new_n479), .A3(G126), .A4(G2105), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT70), .A2(G114), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT70), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2105), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(G102), .A2(G2105), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(G2104), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n503), .A2(KEYINPUT71), .A3(new_n508), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n502), .B1(new_n511), .B2(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT5), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(G543), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n524), .A2(G88), .B1(new_n525), .B2(G50), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n522), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT74), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n524), .A2(G89), .B1(new_n525), .B2(G51), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT73), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n521), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n519), .A2(new_n523), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT75), .B(G90), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n523), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n537), .A2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n516), .A2(new_n518), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n521), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n549), .B1(new_n548), .B2(new_n547), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n524), .A2(G81), .B1(new_n525), .B2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT78), .Z(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT79), .Z(G188));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(KEYINPUT80), .B2(KEYINPUT9), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n525), .B(new_n563), .C1(KEYINPUT80), .C2(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n524), .A2(G91), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n566), .B(new_n567), .C1(new_n540), .C2(new_n562), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n564), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n521), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND2_X1  g149(.A1(new_n522), .A2(new_n526), .ZN(G303));
  NAND2_X1  g150(.A1(new_n524), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n525), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n545), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n525), .ZN(new_n583));
  AND3_X1   g158(.A1(new_n519), .A2(G86), .A3(new_n523), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT81), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT81), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n524), .A2(G85), .B1(new_n525), .B2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n521), .B2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n519), .A2(G66), .ZN(new_n592));
  INV_X1    g167(.A(G79), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT83), .B1(new_n593), .B2(new_n515), .ZN(new_n594));
  OR3_X1    g169(.A1(new_n593), .A2(new_n515), .A3(KEYINPUT83), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n525), .A2(KEYINPUT82), .ZN(new_n597));
  INV_X1    g172(.A(G54), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n598), .B1(new_n540), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(G651), .A2(new_n596), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n519), .A2(G92), .A3(new_n523), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n591), .B1(new_n606), .B2(G868), .ZN(G321));
  XOR2_X1   g182(.A(G321), .B(KEYINPUT84), .Z(G284));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G299), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NOR2_X1   g189(.A1(new_n605), .A2(G559), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  MUX2_X1   g192(.A(new_n552), .B(new_n617), .S(G868), .Z(G323));
  XOR2_X1   g193(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n619));
  XNOR2_X1  g194(.A(G323), .B(new_n619), .ZN(G282));
  NAND2_X1  g195(.A1(new_n489), .A2(G123), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n461), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n495), .A2(G135), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n481), .A2(new_n468), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n628), .A2(new_n629), .A3(new_n634), .ZN(G156));
  INV_X1    g210(.A(G14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n636), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n650), .A2(KEYINPUT88), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(KEYINPUT88), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n653), .A2(KEYINPUT89), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(KEYINPUT89), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT90), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT18), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n658), .B(KEYINPUT17), .ZN(new_n663));
  INV_X1    g238(.A(new_n657), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n663), .A2(new_n659), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT92), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n664), .B1(new_n658), .B2(new_n659), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  AOI22_X1  g243(.A1(new_n668), .A2(KEYINPUT91), .B1(new_n659), .B2(new_n663), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(KEYINPUT91), .B2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n662), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT93), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n679), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n682), .A2(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(KEYINPUT20), .ZN(new_n684));
  OAI221_X1 g259(.A(new_n681), .B1(new_n679), .B2(new_n677), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n689), .ZN(new_n692));
  AND3_X1   g267(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n691), .B1(new_n690), .B2(new_n692), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(G229));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G22), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1971), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT32), .B(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT94), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(G6), .ZN(new_n703));
  INV_X1    g278(.A(G305), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n696), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n699), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n702), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n709));
  NAND2_X1  g284(.A1(G288), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n576), .A2(new_n578), .A3(KEYINPUT95), .A4(new_n577), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n708), .B1(new_n712), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n706), .A2(new_n707), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n489), .A2(G119), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n461), .A2(G107), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n495), .A2(G131), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G25), .B2(G29), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  AND2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  MUX2_X1   g306(.A(G24), .B(G290), .S(G16), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1986), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n718), .A2(new_n719), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n719), .B1(new_n718), .B2(new_n734), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G2090), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n740), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(KEYINPUT29), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n740), .A2(G32), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT101), .B(KEYINPUT26), .Z(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n481), .A2(G105), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G141), .B2(new_n495), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n489), .A2(G129), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n746), .B1(new_n755), .B2(new_n740), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n696), .A2(G20), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT23), .ZN(new_n760));
  INV_X1    g335(.A(G299), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(new_n696), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G168), .A2(new_n696), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n696), .B2(G21), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n740), .B1(new_n768), .B2(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n768), .B2(G34), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G160), .B2(G29), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n766), .A2(new_n767), .B1(G2084), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n766), .A2(new_n767), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n740), .A2(G33), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(new_n461), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT100), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n495), .A2(G139), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n774), .B1(new_n782), .B2(new_n740), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n783), .A2(G2072), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n773), .A2(new_n784), .ZN(new_n785));
  OAI22_X1  g360(.A1(new_n783), .A2(G2072), .B1(G2084), .B2(new_n771), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n627), .A2(new_n740), .ZN(new_n787));
  NOR2_X1   g362(.A1(G171), .A2(new_n696), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n696), .A2(G5), .ZN(new_n789));
  OAI21_X1  g364(.A(G1961), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G11), .ZN(new_n791));
  INV_X1    g366(.A(G28), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(KEYINPUT30), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n740), .B1(new_n794), .B2(G28), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n790), .B(new_n791), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n788), .A2(G1961), .A3(new_n789), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n786), .A2(new_n787), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n764), .A2(new_n772), .A3(new_n785), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n740), .A2(G27), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n740), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2078), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n745), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n696), .A2(G4), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n606), .B2(new_n696), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT96), .B(G1348), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT97), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n805), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n696), .A2(G19), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n553), .B2(new_n696), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(G1341), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(G1341), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n808), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n740), .A2(G26), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT28), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n489), .A2(G128), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n461), .A2(G116), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n495), .A2(G140), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(G29), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT98), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(G2067), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(G2067), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n813), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n743), .A2(new_n739), .A3(new_n744), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n743), .A2(KEYINPUT102), .A3(new_n739), .A4(new_n744), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n803), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n738), .A2(new_n834), .ZN(G311));
  OAI21_X1  g410(.A(KEYINPUT103), .B1(new_n738), .B2(new_n834), .ZN(new_n836));
  INV_X1    g411(.A(new_n834), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n838));
  INV_X1    g413(.A(new_n737), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n735), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n836), .A2(new_n841), .ZN(G150));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  INV_X1    g418(.A(G67), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n545), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n521), .B1(new_n845), .B2(KEYINPUT104), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(KEYINPUT104), .B2(new_n845), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n524), .A2(G93), .B1(new_n525), .B2(G55), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n605), .A2(new_n613), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n552), .A2(new_n849), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n550), .A2(new_n847), .A3(new_n551), .A4(new_n848), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n853), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT105), .ZN(new_n861));
  INV_X1    g436(.A(G860), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n858), .B2(new_n859), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n851), .B1(new_n861), .B2(new_n863), .ZN(G145));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n489), .A2(G130), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G118), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n867), .A2(new_n868), .B1(new_n870), .B2(G2105), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n495), .A2(G142), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n754), .A2(new_n821), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n754), .A2(new_n821), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n873), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n725), .B(new_n632), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n502), .A2(new_n509), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n878), .A2(new_n880), .A3(new_n882), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n884), .B2(new_n887), .ZN(new_n890));
  OAI22_X1  g465(.A1(new_n889), .A2(new_n890), .B1(new_n781), .B2(new_n777), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n782), .A3(new_n888), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n626), .B(G160), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G162), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n895), .B1(new_n891), .B2(new_n893), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n865), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n901), .A2(new_n896), .A3(KEYINPUT40), .A4(new_n897), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(G395));
  XNOR2_X1  g478(.A(new_n712), .B(G290), .ZN(new_n904));
  NAND2_X1  g479(.A1(G166), .A2(KEYINPUT107), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n906));
  NAND2_X1  g481(.A1(G303), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n905), .A2(G305), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G305), .B1(new_n905), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n710), .A2(new_n711), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(G290), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n617), .B(new_n857), .ZN(new_n916));
  NAND2_X1  g491(.A1(G299), .A2(new_n605), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(G299), .A2(new_n605), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n918), .B2(new_n919), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n761), .A2(new_n606), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n917), .A3(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n916), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n921), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n922), .B1(new_n921), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n915), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n921), .A2(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n910), .A2(new_n914), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n921), .A2(new_n922), .A3(new_n928), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n936), .A3(G868), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT108), .B1(new_n849), .B2(new_n609), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n931), .A2(new_n936), .A3(KEYINPUT108), .A4(G868), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(G295));
  AND2_X1   g516(.A1(new_n939), .A2(new_n940), .ZN(G331));
  NAND2_X1  g517(.A1(G168), .A2(G171), .ZN(new_n943));
  OAI21_X1  g518(.A(G301), .B1(new_n532), .B2(new_n534), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n856), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n854), .A2(new_n944), .A3(new_n855), .A4(new_n943), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n920), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n856), .B2(new_n945), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n856), .A2(new_n945), .A3(new_n950), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n934), .B(new_n948), .C1(new_n954), .C2(new_n927), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n897), .ZN(new_n956));
  INV_X1    g531(.A(new_n953), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n947), .B1(new_n957), .B2(new_n951), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(new_n924), .A3(new_n926), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n934), .B1(new_n959), .B2(new_n948), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT43), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n920), .A2(new_n947), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n952), .B2(new_n953), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n927), .B1(new_n947), .B2(new_n946), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n915), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n955), .A2(new_n967), .A3(new_n968), .A4(new_n897), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n956), .C2(new_n960), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n970), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n963), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n956), .A2(new_n960), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n977), .B2(new_n968), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n955), .A2(new_n967), .A3(new_n897), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT112), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n955), .A2(new_n967), .A3(new_n981), .A4(new_n897), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(KEYINPUT43), .A3(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n978), .A2(new_n983), .A3(KEYINPUT113), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT113), .B1(new_n978), .B2(new_n983), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n976), .B1(new_n984), .B2(new_n985), .ZN(G397));
  INV_X1    g561(.A(G1996), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n754), .B(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G2067), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n821), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n726), .A2(new_n729), .ZN(new_n992));
  OAI22_X1  g567(.A1(new_n991), .A2(new_n992), .B1(G2067), .B2(new_n821), .ZN(new_n993));
  INV_X1    g568(.A(new_n509), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n468), .A2(new_n501), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n466), .A2(KEYINPUT64), .ZN(new_n999));
  NAND2_X1  g574(.A1(G113), .A2(G2104), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n470), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G2105), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n480), .A2(new_n482), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(G40), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n998), .A2(new_n1004), .A3(KEYINPUT45), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n993), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1005), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1007), .A2(G1986), .A3(G290), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n1008), .B(KEYINPUT127), .Z(new_n1009));
  INV_X1    g584(.A(KEYINPUT48), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(new_n725), .B(new_n729), .Z(new_n1012));
  NOR2_X1   g587(.A1(new_n991), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT46), .B1(new_n1005), .B2(new_n987), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n990), .A2(new_n755), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(new_n1005), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1005), .A2(KEYINPUT46), .A3(new_n987), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1020), .A2(KEYINPUT126), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(KEYINPUT126), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1014), .A2(new_n1015), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g599(.A(new_n1006), .B(new_n1024), .C1(new_n1016), .C2(new_n1023), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g601(.A(G1384), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1026), .B(new_n1027), .C1(new_n502), .C2(new_n509), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1004), .A2(G2084), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n511), .A2(new_n512), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1030), .B2(new_n997), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1028), .B(new_n1029), .C1(new_n1031), .C2(new_n1026), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  NOR3_X1   g610(.A1(G164), .A2(new_n1035), .A3(G1384), .ZN(new_n1036));
  INV_X1    g611(.A(G40), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n471), .A2(new_n483), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n767), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1041), .A2(KEYINPUT117), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1034), .A2(G168), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(G8), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1027), .B1(new_n502), .B2(new_n509), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1004), .B1(new_n1035), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n503), .A2(KEYINPUT71), .A3(new_n508), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT71), .B1(new_n503), .B2(new_n508), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n997), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(KEYINPUT45), .A3(new_n1027), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1966), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1026), .B1(new_n1049), .B2(new_n1027), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1028), .ZN(new_n1053));
  INV_X1    g628(.A(G2084), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1038), .A2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1051), .B1(new_n1056), .B2(KEYINPUT117), .ZN(new_n1057));
  AOI21_X1  g632(.A(G168), .B1(new_n1057), .B2(new_n1034), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT51), .B1(new_n1044), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1043), .A2(new_n1060), .A3(G8), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT62), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1059), .A2(new_n1064), .A3(new_n1061), .ZN(new_n1065));
  INV_X1    g640(.A(G8), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G166), .A2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n1068));
  OR2_X1    g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(KEYINPUT114), .B2(KEYINPUT55), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1041), .A2(new_n1028), .A3(new_n1038), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(G2090), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1049), .A2(new_n1027), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1035), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1004), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1971), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(G8), .B(new_n1071), .C1(new_n1073), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT115), .B(G1981), .Z(new_n1080));
  NOR2_X1   g655(.A1(G305), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1981), .ZN(new_n1082));
  INV_X1    g657(.A(new_n584), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n583), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1084), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1086), .B(KEYINPUT49), .C1(G305), .C2(new_n1080), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1066), .B1(new_n998), .B2(new_n1038), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1976), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT52), .B1(G288), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1088), .B(new_n1091), .C1(new_n1090), .C2(new_n912), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1088), .B1(new_n1090), .B2(new_n912), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1089), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1038), .B1(new_n998), .B2(new_n1026), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1096), .A2(KEYINPUT116), .B1(new_n1031), .B2(new_n1026), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1004), .B1(KEYINPUT50), .B2(new_n1045), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n739), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1077), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1066), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1078), .B(new_n1095), .C1(new_n1103), .C2(new_n1071), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(G2078), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT123), .B(G1961), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1072), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1105), .A2(G2078), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1046), .A2(new_n1050), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G171), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1104), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1063), .A2(new_n1065), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(G288), .A2(G1976), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1089), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1088), .B1(new_n1117), .B2(new_n1081), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1095), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n1078), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G286), .A2(new_n1066), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1053), .B1(new_n1074), .B2(KEYINPUT50), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT117), .B1(new_n1125), .B2(new_n1029), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1122), .B(new_n1123), .C1(new_n1124), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1034), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1122), .B1(new_n1129), .B2(new_n1123), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1121), .B1(new_n1131), .B2(new_n1104), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1095), .A2(new_n1078), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n1134));
  OAI21_X1  g709(.A(G8), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1071), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1133), .B(new_n1137), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1120), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1038), .B1(new_n1045), .B2(new_n1035), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1035), .B2(new_n1074), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(G2072), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(G299), .B(KEYINPUT57), .Z(new_n1145));
  INV_X1    g720(.A(new_n1100), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n1098), .A2(new_n1099), .B1(new_n1074), .B2(KEYINPUT50), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1144), .B(new_n1145), .C1(new_n1148), .C2(G1956), .ZN(new_n1149));
  INV_X1    g724(.A(G1348), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n998), .A2(new_n1038), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(G2067), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1004), .A2(new_n1045), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(KEYINPUT121), .A3(new_n989), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1072), .A2(new_n1150), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(new_n605), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1149), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(G1956), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1161), .A2(KEYINPUT122), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1145), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1161), .B2(KEYINPUT122), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1158), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT61), .B1(new_n1166), .B2(new_n1149), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n605), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n605), .A2(new_n1168), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1169), .B1(new_n1156), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1072), .A2(new_n1150), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1173));
  AND4_X1   g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1170), .A4(new_n1169), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1106), .A2(G1996), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT58), .B(G1341), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1154), .A2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g753(.A(KEYINPUT59), .B(new_n553), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT59), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1141), .B2(new_n987), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(new_n552), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1167), .A2(new_n1175), .A3(new_n1183), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1149), .A2(KEYINPUT61), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1165), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  OR2_X1    g762(.A1(new_n1112), .A2(G171), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT54), .ZN(new_n1189));
  AOI211_X1 g764(.A(new_n1105), .B(G2078), .C1(new_n998), .C2(KEYINPUT45), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1046), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1107), .A2(new_n1109), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1189), .B1(new_n1192), .B2(G171), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1104), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(G171), .B1(new_n1190), .B2(new_n1046), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1107), .A2(new_n1109), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(KEYINPUT124), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1113), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1196), .A2(KEYINPUT124), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1189), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1194), .A2(new_n1200), .A3(new_n1062), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1115), .B(new_n1139), .C1(new_n1187), .C2(new_n1201), .ZN(new_n1202));
  XOR2_X1   g777(.A(G290), .B(G1986), .Z(new_n1203));
  NAND2_X1  g778(.A1(new_n1013), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1005), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1202), .A2(KEYINPUT125), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(KEYINPUT125), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1025), .B1(new_n1206), .B2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g783(.A1(new_n901), .A2(new_n897), .A3(new_n896), .ZN(new_n1210));
  NOR2_X1   g784(.A1(G227), .A2(new_n459), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n1211), .B1(new_n693), .B2(new_n694), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1212), .B1(new_n654), .B2(new_n655), .ZN(new_n1213));
  NAND3_X1  g787(.A1(new_n1210), .A2(new_n974), .A3(new_n1213), .ZN(G225));
  INV_X1    g788(.A(G225), .ZN(G308));
endmodule


