

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579;

  XOR2_X1 U322 ( .A(n382), .B(KEYINPUT41), .Z(n553) );
  XOR2_X1 U323 ( .A(G71GAT), .B(G120GAT), .Z(n361) );
  XNOR2_X1 U324 ( .A(n394), .B(n368), .ZN(n369) );
  INV_X1 U325 ( .A(KEYINPUT121), .ZN(n448) );
  XNOR2_X1 U326 ( .A(n370), .B(n369), .ZN(n374) );
  XNOR2_X1 U327 ( .A(n448), .B(KEYINPUT55), .ZN(n449) );
  XNOR2_X1 U328 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U329 ( .A(KEYINPUT28), .B(n465), .Z(n527) );
  XNOR2_X1 U330 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n291) );
  XNOR2_X1 U333 ( .A(G134GAT), .B(G106GAT), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n300) );
  XOR2_X1 U335 ( .A(G36GAT), .B(G190GAT), .Z(n397) );
  XOR2_X1 U336 ( .A(G29GAT), .B(G43GAT), .Z(n293) );
  XNOR2_X1 U337 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n355) );
  XOR2_X1 U339 ( .A(n397), .B(n355), .Z(n295) );
  NAND2_X1 U340 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U342 ( .A(n296), .B(KEYINPUT11), .Z(n298) );
  XOR2_X1 U343 ( .A(G50GAT), .B(G162GAT), .Z(n441) );
  XNOR2_X1 U344 ( .A(G218GAT), .B(n441), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U347 ( .A(KEYINPUT72), .B(G85GAT), .Z(n302) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G92GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U350 ( .A(KEYINPUT73), .B(n303), .Z(n372) );
  XOR2_X1 U351 ( .A(n304), .B(n372), .Z(n549) );
  XOR2_X1 U352 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n306) );
  XNOR2_X1 U353 ( .A(KEYINPUT82), .B(KEYINPUT81), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U355 ( .A(G183GAT), .B(KEYINPUT19), .Z(n307) );
  XOR2_X1 U356 ( .A(n308), .B(n307), .Z(n399) );
  XOR2_X1 U357 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n310) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(G176GAT), .ZN(n309) );
  XOR2_X1 U359 ( .A(n310), .B(n309), .Z(n323) );
  XOR2_X1 U360 ( .A(G99GAT), .B(G190GAT), .Z(n312) );
  XNOR2_X1 U361 ( .A(G43GAT), .B(G15GAT), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U363 ( .A(n361), .B(n313), .Z(n315) );
  NAND2_X1 U364 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n317) );
  INV_X1 U366 ( .A(KEYINPUT20), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U368 ( .A(KEYINPUT0), .B(G127GAT), .Z(n319) );
  XNOR2_X1 U369 ( .A(G113GAT), .B(G134GAT), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n422) );
  XNOR2_X1 U371 ( .A(n422), .B(KEYINPUT83), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U373 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X2 U374 ( .A(n399), .B(n324), .Z(n517) );
  XOR2_X1 U375 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n326) );
  XNOR2_X1 U376 ( .A(G183GAT), .B(G64GAT), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U378 ( .A(G211GAT), .B(KEYINPUT76), .Z(n328) );
  XNOR2_X1 U379 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n341) );
  XOR2_X1 U382 ( .A(KEYINPUT13), .B(G57GAT), .Z(n360) );
  XOR2_X1 U383 ( .A(G78GAT), .B(G71GAT), .Z(n332) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(G22GAT), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U386 ( .A(n360), .B(n333), .Z(n335) );
  NAND2_X1 U387 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U389 ( .A(n336), .B(G155GAT), .Z(n339) );
  XNOR2_X1 U390 ( .A(G1GAT), .B(KEYINPUT68), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n337), .B(G15GAT), .ZN(n354) );
  XNOR2_X1 U392 ( .A(n354), .B(G127GAT), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U394 ( .A(n341), .B(n340), .Z(n469) );
  INV_X1 U395 ( .A(n469), .ZN(n572) );
  XOR2_X1 U396 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n343) );
  XNOR2_X1 U397 ( .A(KEYINPUT29), .B(G197GAT), .ZN(n342) );
  XOR2_X1 U398 ( .A(n343), .B(n342), .Z(n347) );
  XOR2_X1 U399 ( .A(G50GAT), .B(G36GAT), .Z(n345) );
  XOR2_X1 U400 ( .A(G169GAT), .B(G8GAT), .Z(n400) );
  XOR2_X1 U401 ( .A(G22GAT), .B(G141GAT), .Z(n442) );
  XNOR2_X1 U402 ( .A(n400), .B(n442), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n349) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U407 ( .A(KEYINPUT65), .B(G113GAT), .Z(n351) );
  XNOR2_X1 U408 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U410 ( .A(n353), .B(n352), .Z(n357) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U412 ( .A(n357), .B(n356), .Z(n498) );
  INV_X1 U413 ( .A(n498), .ZN(n566) );
  XOR2_X1 U414 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n359) );
  XNOR2_X1 U415 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n358) );
  XOR2_X1 U416 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U417 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n363) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U421 ( .A(G204GAT), .B(KEYINPUT74), .Z(n367) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(G64GAT), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n394) );
  NAND2_X1 U424 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(G106GAT), .B(G78GAT), .ZN(n371) );
  XNOR2_X1 U426 ( .A(n371), .B(G148GAT), .ZN(n436) );
  XOR2_X1 U427 ( .A(n372), .B(n436), .Z(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n382) );
  NAND2_X1 U429 ( .A1(n566), .A2(n553), .ZN(n375) );
  XOR2_X1 U430 ( .A(n375), .B(KEYINPUT46), .Z(n376) );
  NOR2_X1 U431 ( .A1(n572), .A2(n376), .ZN(n377) );
  XOR2_X1 U432 ( .A(KEYINPUT114), .B(n377), .Z(n378) );
  NOR2_X1 U433 ( .A1(n549), .A2(n378), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n379), .B(KEYINPUT47), .ZN(n386) );
  XOR2_X1 U435 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n381) );
  XNOR2_X1 U436 ( .A(KEYINPUT36), .B(n549), .ZN(n576) );
  NAND2_X1 U437 ( .A1(n572), .A2(n576), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n384) );
  NOR2_X1 U439 ( .A1(n566), .A2(n382), .ZN(n383) );
  NAND2_X1 U440 ( .A1(n384), .A2(n383), .ZN(n385) );
  NAND2_X1 U441 ( .A1(n386), .A2(n385), .ZN(n388) );
  XOR2_X1 U442 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n525) );
  XOR2_X1 U444 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n390) );
  NAND2_X1 U445 ( .A1(G226GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n393) );
  XOR2_X1 U447 ( .A(KEYINPUT21), .B(G211GAT), .Z(n392) );
  XNOR2_X1 U448 ( .A(G197GAT), .B(G218GAT), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n435) );
  XOR2_X1 U450 ( .A(n393), .B(n435), .Z(n396) );
  XNOR2_X1 U451 ( .A(G92GAT), .B(n394), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U453 ( .A(n398), .B(n397), .Z(n402) );
  XNOR2_X1 U454 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U455 ( .A(n402), .B(n401), .Z(n515) );
  INV_X1 U456 ( .A(n515), .ZN(n454) );
  NAND2_X1 U457 ( .A1(n525), .A2(n454), .ZN(n404) );
  XOR2_X1 U458 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n563) );
  XOR2_X1 U460 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n406) );
  XNOR2_X1 U461 ( .A(G155GAT), .B(KEYINPUT85), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n439) );
  XOR2_X1 U463 ( .A(n439), .B(G162GAT), .Z(n408) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U466 ( .A(G29GAT), .B(n409), .ZN(n429) );
  XOR2_X1 U467 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n411) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(G120GAT), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U470 ( .A(G57GAT), .B(G148GAT), .Z(n413) );
  XNOR2_X1 U471 ( .A(G1GAT), .B(G85GAT), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n427) );
  XOR2_X1 U474 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n417) );
  XNOR2_X1 U475 ( .A(KEYINPUT88), .B(KEYINPUT92), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U477 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n419) );
  XNOR2_X1 U478 ( .A(KEYINPUT4), .B(KEYINPUT90), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U481 ( .A(n422), .B(KEYINPUT89), .Z(n423) );
  XNOR2_X1 U482 ( .A(KEYINPUT6), .B(n423), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U485 ( .A(n429), .B(n428), .Z(n463) );
  XOR2_X1 U486 ( .A(KEYINPUT84), .B(KEYINPUT22), .Z(n431) );
  XNOR2_X1 U487 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n446) );
  XOR2_X1 U489 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n433) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U492 ( .A(n434), .B(KEYINPUT23), .Z(n438) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n465) );
  NOR2_X1 U499 ( .A1(n463), .A2(n465), .ZN(n447) );
  AND2_X1 U500 ( .A1(n563), .A2(n447), .ZN(n450) );
  NOR2_X1 U501 ( .A1(n517), .A2(n451), .ZN(n558) );
  NAND2_X1 U502 ( .A1(n549), .A2(n558), .ZN(n453) );
  INV_X1 U503 ( .A(n463), .ZN(n562) );
  NOR2_X1 U504 ( .A1(n382), .A2(n498), .ZN(n486) );
  INV_X1 U505 ( .A(n517), .ZN(n528) );
  NAND2_X1 U506 ( .A1(n454), .A2(n528), .ZN(n455) );
  XOR2_X1 U507 ( .A(KEYINPUT98), .B(n455), .Z(n456) );
  NOR2_X1 U508 ( .A1(n465), .A2(n456), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(KEYINPUT99), .ZN(n458) );
  XNOR2_X1 U510 ( .A(n458), .B(KEYINPUT25), .ZN(n461) );
  NAND2_X1 U511 ( .A1(n465), .A2(n517), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n459), .B(KEYINPUT26), .ZN(n565) );
  XNOR2_X1 U513 ( .A(n515), .B(KEYINPUT27), .ZN(n464) );
  NOR2_X1 U514 ( .A1(n565), .A2(n464), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n461), .A2(n460), .ZN(n462) );
  NOR2_X1 U516 ( .A1(n463), .A2(n462), .ZN(n468) );
  NOR2_X1 U517 ( .A1(n464), .A2(n562), .ZN(n526) );
  NAND2_X1 U518 ( .A1(n526), .A2(n527), .ZN(n466) );
  NOR2_X1 U519 ( .A1(n466), .A2(n528), .ZN(n467) );
  NOR2_X1 U520 ( .A1(n468), .A2(n467), .ZN(n483) );
  NOR2_X1 U521 ( .A1(n549), .A2(n469), .ZN(n470) );
  XOR2_X1 U522 ( .A(KEYINPUT78), .B(n470), .Z(n471) );
  XNOR2_X1 U523 ( .A(n471), .B(KEYINPUT16), .ZN(n472) );
  NOR2_X1 U524 ( .A1(n483), .A2(n472), .ZN(n500) );
  NAND2_X1 U525 ( .A1(n486), .A2(n500), .ZN(n480) );
  NOR2_X1 U526 ( .A1(n562), .A2(n480), .ZN(n474) );
  XNOR2_X1 U527 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n473) );
  XNOR2_X1 U528 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U529 ( .A(G1GAT), .B(n475), .Z(G1324GAT) );
  NOR2_X1 U530 ( .A1(n515), .A2(n480), .ZN(n476) );
  XOR2_X1 U531 ( .A(G8GAT), .B(n476), .Z(G1325GAT) );
  NOR2_X1 U532 ( .A1(n517), .A2(n480), .ZN(n478) );
  XNOR2_X1 U533 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U535 ( .A(G15GAT), .B(n479), .Z(G1326GAT) );
  NOR2_X1 U536 ( .A1(n527), .A2(n480), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT102), .B(n481), .Z(n482) );
  XNOR2_X1 U538 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  NOR2_X1 U539 ( .A1(n572), .A2(n483), .ZN(n484) );
  NAND2_X1 U540 ( .A1(n576), .A2(n484), .ZN(n485) );
  XNOR2_X1 U541 ( .A(KEYINPUT37), .B(n485), .ZN(n513) );
  NAND2_X1 U542 ( .A1(n486), .A2(n513), .ZN(n487) );
  XNOR2_X1 U543 ( .A(n487), .B(KEYINPUT104), .ZN(n488) );
  XNOR2_X1 U544 ( .A(n488), .B(KEYINPUT38), .ZN(n496) );
  NOR2_X1 U545 ( .A1(n562), .A2(n496), .ZN(n491) );
  XOR2_X1 U546 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(n489), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U549 ( .A1(n515), .A2(n496), .ZN(n492) );
  XOR2_X1 U550 ( .A(G36GAT), .B(n492), .Z(G1329GAT) );
  NOR2_X1 U551 ( .A1(n517), .A2(n496), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U555 ( .A1(n527), .A2(n496), .ZN(n497) );
  XOR2_X1 U556 ( .A(G50GAT), .B(n497), .Z(G1331GAT) );
  NAND2_X1 U557 ( .A1(n498), .A2(n553), .ZN(n499) );
  XOR2_X1 U558 ( .A(KEYINPUT106), .B(n499), .Z(n512) );
  NAND2_X1 U559 ( .A1(n500), .A2(n512), .ZN(n508) );
  NOR2_X1 U560 ( .A1(n562), .A2(n508), .ZN(n501) );
  XOR2_X1 U561 ( .A(G57GAT), .B(n501), .Z(n502) );
  XNOR2_X1 U562 ( .A(KEYINPUT42), .B(n502), .ZN(G1332GAT) );
  NOR2_X1 U563 ( .A1(n515), .A2(n508), .ZN(n504) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1333GAT) );
  NOR2_X1 U566 ( .A1(n517), .A2(n508), .ZN(n506) );
  XNOR2_X1 U567 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  NOR2_X1 U570 ( .A1(n527), .A2(n508), .ZN(n510) );
  XNOR2_X1 U571 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U574 ( .A1(n513), .A2(n512), .ZN(n522) );
  NOR2_X1 U575 ( .A1(n562), .A2(n522), .ZN(n514) );
  XOR2_X1 U576 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U577 ( .A1(n515), .A2(n522), .ZN(n516) );
  XOR2_X1 U578 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U579 ( .A1(n517), .A2(n522), .ZN(n519) );
  XNOR2_X1 U580 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n519), .B(n518), .ZN(G1338GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n521) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n524) );
  NOR2_X1 U585 ( .A1(n527), .A2(n522), .ZN(n523) );
  XOR2_X1 U586 ( .A(n524), .B(n523), .Z(G1339GAT) );
  NAND2_X1 U587 ( .A1(n525), .A2(n526), .ZN(n540) );
  NAND2_X1 U588 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U589 ( .A1(n540), .A2(n529), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n536), .A2(n566), .ZN(n530) );
  XNOR2_X1 U591 ( .A(n530), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U593 ( .A1(n536), .A2(n553), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  NAND2_X1 U596 ( .A1(n536), .A2(n572), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n538) );
  NAND2_X1 U600 ( .A1(n536), .A2(n549), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U602 ( .A(G134GAT), .B(n539), .Z(G1343GAT) );
  NOR2_X1 U603 ( .A1(n565), .A2(n540), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n566), .A2(n548), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n541), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n543) );
  NAND2_X1 U607 ( .A1(n548), .A2(n553), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(n544), .ZN(G1345GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n546) );
  NAND2_X1 U611 ( .A1(n548), .A2(n572), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U616 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n566), .A2(n558), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1348GAT) );
  NAND2_X1 U619 ( .A1(n558), .A2(n553), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT123), .Z(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n572), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U626 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT60), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT59), .B(n561), .Z(n568) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n577) );
  NAND2_X1 U631 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n577), .A2(n382), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(G204GAT), .B(n571), .Z(G1353GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n574) );
  NAND2_X1 U638 ( .A1(n577), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

