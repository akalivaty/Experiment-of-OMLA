//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n454));
  XOR2_X1   g029(.A(new_n453), .B(new_n454), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(new_n456), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT67), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n473), .A3(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(G101), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n473), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(G2105), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n469), .A2(new_n477), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT68), .ZN(G160));
  NOR2_X1   g060(.A1(new_n479), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(new_n468), .B2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n479), .B2(new_n468), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n466), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(G124), .B2(new_n494), .ZN(G162));
  NAND3_X1  g070(.A1(new_n471), .A2(new_n473), .A3(G126), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n470), .A2(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G102), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n468), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n466), .A2(KEYINPUT4), .A3(G138), .A4(new_n468), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n499), .A2(new_n501), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n513), .A2(new_n515), .A3(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(G50), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n513), .A2(new_n515), .A3(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(G166));
  NAND2_X1  g098(.A1(new_n513), .A2(new_n515), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n511), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n510), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(new_n531), .A3(new_n508), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT71), .B1(new_n509), .B2(new_n510), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(new_n533), .A3(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n529), .A2(new_n536), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AOI22_X1  g115(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT72), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT73), .B(G52), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n524), .A2(new_n511), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n535), .A2(new_n544), .B1(G90), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  XOR2_X1   g122(.A(KEYINPUT74), .B(G81), .Z(new_n548));
  NOR3_X1   g123(.A1(new_n511), .A2(new_n548), .A3(new_n524), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n525), .A2(G56), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n519), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI211_X1 g127(.A(new_n549), .B(new_n552), .C1(G43), .C2(new_n535), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  AOI22_X1  g134(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n519), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n545), .A2(G91), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n535), .A2(KEYINPUT9), .A3(G53), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n534), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(new_n543), .A2(new_n546), .ZN(G301));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n545), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n534), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT75), .Z(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n524), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(G48), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n524), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(new_n526), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n545), .A2(G85), .ZN(new_n585));
  XNOR2_X1  g160(.A(KEYINPUT76), .B(G47), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI221_X1 g162(.A(new_n585), .B1(new_n534), .B2(new_n586), .C1(new_n587), .C2(new_n519), .ZN(G290));
  NAND2_X1  g163(.A1(new_n545), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  NAND2_X1  g165(.A1(new_n535), .A2(G54), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n519), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G171), .B2(new_n595), .ZN(G284));
  OAI21_X1  g172(.A(new_n596), .B1(G171), .B2(new_n595), .ZN(G321));
  OR3_X1    g173(.A1(G168), .A2(KEYINPUT77), .A3(new_n595), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT77), .B1(G168), .B2(new_n595), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(G868), .C2(new_n601), .ZN(G297));
  OAI211_X1 g177(.A(new_n599), .B(new_n600), .C1(G868), .C2(new_n601), .ZN(G280));
  INV_X1    g178(.A(new_n594), .ZN(new_n604));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G860), .ZN(G148));
  INV_X1    g181(.A(new_n553), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n595), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n594), .A2(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g186(.A1(new_n468), .A2(G111), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n470), .B1(new_n612), .B2(KEYINPUT78), .ZN(new_n613));
  OAI221_X1 g188(.A(new_n613), .B1(KEYINPUT78), .B2(new_n612), .C1(G99), .C2(G2105), .ZN(new_n614));
  INV_X1    g189(.A(G135), .ZN(new_n615));
  INV_X1    g190(.A(new_n486), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(G123), .B2(new_n494), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n466), .A2(new_n500), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT79), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2430), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT80), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT16), .B(G2443), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2446), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n635), .B(new_n637), .Z(new_n638));
  AND2_X1   g213(.A1(new_n638), .A2(G14), .ZN(G401));
  XOR2_X1   g214(.A(G2067), .B(G2678), .Z(new_n640));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  AND2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n640), .B2(new_n641), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n646), .ZN(new_n648));
  INV_X1    g223(.A(new_n640), .ZN(new_n649));
  INV_X1    g224(.A(new_n641), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n650), .A3(new_n644), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT82), .B(G2096), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n658), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  AOI22_X1  g239(.A1(new_n662), .A2(KEYINPUT20), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n658), .A3(new_n661), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n665), .B(new_n667), .C1(KEYINPUT20), .C2(new_n662), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1986), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1991), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(G229));
  MUX2_X1   g249(.A(G23), .B(new_n573), .S(G16), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT33), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G6), .ZN(new_n680));
  INV_X1    g255(.A(G305), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT32), .B(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(G22), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n679), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT87), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n684), .B1(new_n688), .B2(G1971), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n678), .B(new_n689), .C1(G1971), .C2(new_n688), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT34), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n679), .A2(G24), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G290), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(G1986), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(KEYINPUT34), .ZN(new_n696));
  AND2_X1   g271(.A1(KEYINPUT83), .A2(G29), .ZN(new_n697));
  NOR2_X1   g272(.A1(KEYINPUT83), .A2(G29), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n486), .A2(G131), .ZN(new_n701));
  NOR2_X1   g276(.A1(G95), .A2(G2105), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(new_n468), .B2(G107), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G119), .B2(new_n494), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT84), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(new_n699), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT35), .B(G1991), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT85), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n711));
  OAI22_X1  g286(.A1(new_n693), .A2(new_n694), .B1(KEYINPUT88), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n691), .A2(new_n695), .A3(new_n696), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(KEYINPUT88), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT89), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n696), .A2(new_n713), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n719), .A2(new_n695), .A3(new_n691), .A4(new_n716), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n699), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G2078), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n679), .A2(G4), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n604), .B2(new_n679), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1348), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n494), .A2(G129), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT26), .Z(new_n731));
  AOI22_X1  g306(.A1(new_n486), .A2(G141), .B1(G105), .B2(new_n500), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G29), .B2(G32), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G21), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G168), .B2(G16), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n736), .A2(new_n737), .B1(new_n739), .B2(G1966), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n736), .B2(new_n737), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n728), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(G29), .A2(G33), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n500), .A2(G103), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT25), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n486), .A2(G139), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n745), .B(new_n746), .C1(new_n468), .C2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2072), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT92), .B(G28), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT30), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n618), .A2(new_n699), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n750), .A2(new_n751), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n752), .A2(new_n755), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n722), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n722), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT29), .B(G2090), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n739), .A2(G1966), .B1(G2078), .B2(new_n724), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n758), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n679), .A2(G5), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G171), .B2(new_n679), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT93), .Z(new_n767));
  INV_X1    g342(.A(G1961), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n742), .B(new_n764), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  OAI21_X1  g345(.A(KEYINPUT23), .B1(new_n601), .B2(new_n679), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n679), .A2(G20), .ZN(new_n772));
  MUX2_X1   g347(.A(KEYINPUT23), .B(new_n771), .S(new_n772), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n679), .A2(G19), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n553), .B2(new_n679), .ZN(new_n776));
  MUX2_X1   g351(.A(new_n775), .B(new_n776), .S(KEYINPUT90), .Z(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(G1341), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT24), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G34), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(G34), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI22_X1  g357(.A1(G160), .A2(G29), .B1(new_n722), .B2(new_n782), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n777), .A2(G1341), .B1(G2084), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n722), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n494), .A2(G128), .ZN(new_n787));
  OR2_X1    g362(.A1(G104), .A2(G2105), .ZN(new_n788));
  INV_X1    g363(.A(G116), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n470), .B1(new_n789), .B2(G2105), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n486), .A2(G140), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G29), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n793), .A2(KEYINPUT91), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(KEYINPUT91), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n786), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n783), .A2(G2084), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n778), .A2(new_n784), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n769), .A2(new_n770), .A3(new_n774), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n721), .A2(new_n725), .A3(new_n801), .ZN(G150));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n803));
  NAND2_X1  g378(.A1(G150), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n721), .A2(KEYINPUT94), .A3(new_n725), .A4(new_n801), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(G311));
  NAND2_X1  g381(.A1(new_n545), .A2(G93), .ZN(new_n807));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  OAI221_X1 g384(.A(new_n807), .B1(new_n534), .B2(new_n808), .C1(new_n809), .C2(new_n519), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT95), .Z(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  NOR2_X1   g389(.A1(new_n594), .A2(new_n605), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n811), .A2(new_n607), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n553), .A2(new_n810), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n817), .B(new_n820), .Z(new_n821));
  OAI21_X1  g396(.A(new_n814), .B1(new_n821), .B2(G860), .ZN(G145));
  XNOR2_X1  g397(.A(G160), .B(new_n618), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G162), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n748), .B(new_n792), .Z(new_n825));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n504), .A2(new_n505), .ZN(new_n827));
  INV_X1    g402(.A(new_n501), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n498), .B2(G2105), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n497), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n466), .B2(G126), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n501), .B1(new_n832), .B2(new_n468), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n504), .A2(new_n505), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT96), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n825), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n733), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n825), .A2(new_n836), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n825), .A2(new_n836), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n734), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n486), .A2(G142), .ZN(new_n843));
  NOR2_X1   g418(.A1(G106), .A2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(new_n468), .B2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G130), .B2(new_n494), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n621), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n705), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n838), .A2(new_n851), .A3(new_n841), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n824), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT97), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n850), .A2(KEYINPUT99), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(KEYINPUT99), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n855), .A2(new_n824), .A3(new_n852), .A4(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT98), .B(G37), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n859), .B(new_n861), .ZN(G395));
  XNOR2_X1  g437(.A(new_n573), .B(G166), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G305), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G290), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n820), .A2(new_n609), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n820), .A2(new_n609), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n594), .B(G299), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT101), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n870), .B(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n874), .A2(new_n868), .A3(new_n867), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n872), .B2(new_n875), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n866), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n872), .A2(new_n875), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n865), .A3(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G868), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n811), .A2(G868), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(G295));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n885), .B2(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n595), .B1(new_n880), .B2(new_n883), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n891), .A2(KEYINPUT102), .A3(new_n886), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(G331));
  INV_X1    g468(.A(new_n874), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  NOR2_X1   g470(.A1(G171), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(G168), .B1(G301), .B2(KEYINPUT103), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n818), .A3(new_n819), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n818), .B2(new_n819), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G286), .B1(G171), .B2(new_n895), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n820), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n896), .A3(new_n899), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n894), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n871), .B1(new_n902), .B2(new_n905), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n871), .ZN(new_n910));
  INV_X1    g485(.A(new_n905), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n896), .B1(new_n904), .B2(new_n899), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n908), .B(new_n910), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n865), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n911), .A2(new_n912), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n866), .B(new_n906), .C1(new_n916), .C2(new_n870), .ZN(new_n917));
  AND4_X1   g492(.A1(KEYINPUT43), .A2(new_n915), .A3(new_n858), .A4(new_n917), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n911), .A2(new_n912), .A3(new_n874), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n870), .B1(new_n902), .B2(new_n905), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n865), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n917), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n915), .A2(new_n924), .A3(new_n858), .A4(new_n917), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n931), .ZN(G397));
  OAI21_X1  g507(.A(KEYINPUT96), .B1(new_n833), .B2(new_n834), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n829), .A2(new_n826), .A3(new_n504), .A4(new_n505), .ZN(new_n934));
  AOI21_X1  g509(.A(G1384), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n935), .A2(KEYINPUT45), .ZN(new_n936));
  INV_X1    g511(.A(G40), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n476), .B2(new_n468), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n469), .A2(new_n483), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(G1996), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n734), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT105), .Z(new_n943));
  INV_X1    g518(.A(new_n940), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n792), .B(new_n797), .ZN(new_n945));
  INV_X1    g520(.A(G1996), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n946), .B2(new_n734), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n709), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n706), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n787), .A2(new_n797), .A3(new_n791), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n940), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n705), .B(new_n949), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n944), .A2(new_n953), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n940), .A2(G1986), .A3(G290), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT48), .Z(new_n956));
  AND3_X1   g531(.A1(new_n948), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n941), .A2(KEYINPUT46), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n941), .A2(KEYINPUT46), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n940), .B1(new_n734), .B2(new_n945), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n952), .A2(new_n957), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n965), .B(new_n966), .C1(new_n833), .C2(new_n834), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n827), .B2(new_n829), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n939), .B(new_n967), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1348), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n939), .A2(new_n973), .A3(new_n968), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n965), .B1(new_n833), .B2(new_n834), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n469), .A2(new_n483), .A3(new_n938), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT117), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n977), .A3(new_n797), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n978), .A3(KEYINPUT60), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT119), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n972), .A2(new_n978), .A3(KEYINPUT119), .A4(KEYINPUT60), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT60), .B1(new_n972), .B2(new_n978), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(new_n594), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n981), .B(new_n982), .C1(new_n594), .C2(new_n984), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT45), .B1(new_n506), .B2(new_n965), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n976), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT45), .B(new_n965), .C1(new_n830), .C2(new_n835), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n975), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT106), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT118), .B(G1996), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n990), .A2(new_n991), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n974), .A2(new_n977), .ZN(new_n997));
  XOR2_X1   g572(.A(KEYINPUT58), .B(G1341), .Z(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n553), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT59), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1000), .A2(new_n1003), .A3(new_n553), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n986), .A2(new_n987), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT56), .B(G2072), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT115), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n990), .A2(new_n991), .A3(new_n994), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT116), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n968), .A2(new_n969), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1010), .B(new_n939), .C1(new_n968), .C2(new_n966), .ZN(new_n1011));
  INV_X1    g586(.A(G1956), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n935), .A2(KEYINPUT45), .B1(new_n993), .B2(KEYINPUT106), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n990), .A4(new_n1007), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1009), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n563), .A2(KEYINPUT113), .A3(new_n566), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1023));
  OAI21_X1  g598(.A(G299), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1023), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(new_n601), .A3(new_n1021), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1017), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT61), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1030), .A2(new_n1009), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1005), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n972), .A2(new_n978), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1028), .B1(new_n594), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1031), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1971), .B1(new_n1014), .B2(new_n990), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1011), .A2(G2090), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G166), .A2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT108), .B(KEYINPUT55), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(KEYINPUT108), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1042), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n574), .A2(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1043), .B1(new_n939), .B2(new_n968), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(new_n573), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1053), .A2(KEYINPUT52), .A3(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT111), .B(G1981), .Z(new_n1058));
  NAND2_X1  g633(.A1(new_n681), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n681), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT49), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1059), .B(KEYINPUT49), .C1(new_n1060), .C2(new_n681), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1054), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1056), .A2(KEYINPUT52), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1057), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n990), .A2(new_n991), .A3(new_n994), .ZN(new_n1069));
  INV_X1    g644(.A(G1971), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n970), .A2(G2090), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1043), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT109), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1046), .B(KEYINPUT109), .C1(new_n1044), .C2(new_n1049), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT110), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1072), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n1082));
  NOR4_X1   g657(.A1(new_n1081), .A2(new_n1078), .A3(new_n1082), .A4(new_n1043), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1052), .B(new_n1068), .C1(new_n1080), .C2(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n970), .A2(G2084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n968), .A2(KEYINPUT45), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n993), .A3(new_n939), .ZN(new_n1087));
  INV_X1    g662(.A(G1966), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT51), .B1(new_n1091), .B2(G168), .ZN(new_n1092));
  OAI21_X1  g667(.A(G8), .B1(new_n1090), .B2(G286), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(KEYINPUT51), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1084), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1069), .B2(G2078), .ZN(new_n1099));
  INV_X1    g674(.A(new_n936), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n481), .A2(G2105), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n938), .A2(KEYINPUT122), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G2078), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(KEYINPUT53), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT122), .B1(new_n938), .B2(new_n1101), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1100), .A2(new_n991), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n970), .A2(new_n768), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1099), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT124), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1099), .A2(new_n1107), .A3(new_n1111), .A4(new_n1108), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(G171), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1103), .A2(KEYINPUT53), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1087), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1099), .A2(new_n1116), .A3(new_n1108), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1117), .B2(G301), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(G171), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT121), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1117), .A2(new_n1122), .A3(G171), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1099), .A2(new_n1107), .A3(G301), .A4(new_n1108), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1121), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1114), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1119), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1039), .A2(new_n1097), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n1131));
  OAI21_X1  g706(.A(G8), .B1(new_n1040), .B2(new_n1072), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1082), .B1(new_n1132), .B2(new_n1078), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1074), .A2(KEYINPUT110), .A3(new_n1079), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n1068), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1065), .A2(new_n1055), .A3(new_n574), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1136), .A2(new_n1059), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1054), .B(KEYINPUT112), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1057), .A2(new_n1067), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1132), .B2(new_n1051), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1141), .A2(G168), .A3(new_n1094), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1094), .A2(G168), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1084), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1139), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1130), .A2(new_n1131), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1131), .B1(new_n1130), .B2(new_n1147), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1095), .A2(KEYINPUT62), .A3(new_n1096), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT62), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1141), .A2(new_n1154), .A3(new_n1052), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1150), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1084), .B1(new_n1123), .B2(new_n1121), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1157), .B(KEYINPUT126), .C1(new_n1152), .C2(new_n1151), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1148), .A2(new_n1149), .A3(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(G290), .B(new_n694), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n948), .B(new_n954), .C1(new_n940), .C2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n964), .B1(new_n1160), .B2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g738(.A1(G229), .A2(new_n464), .ZN(new_n1165));
  NOR2_X1   g739(.A1(G401), .A2(G227), .ZN(new_n1166));
  NAND4_X1  g740(.A1(new_n929), .A2(new_n859), .A3(new_n1165), .A4(new_n1166), .ZN(G225));
  INV_X1    g741(.A(G225), .ZN(G308));
endmodule


