

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581;

  XNOR2_X2 U323 ( .A(n457), .B(n456), .ZN(n534) );
  NOR2_X1 U324 ( .A1(n558), .A2(n557), .ZN(n560) );
  NOR2_X1 U325 ( .A1(n385), .A2(n384), .ZN(n386) );
  NOR2_X1 U326 ( .A1(n578), .A2(n409), .ZN(n410) );
  XNOR2_X1 U327 ( .A(n391), .B(n390), .ZN(n471) );
  XOR2_X1 U328 ( .A(n407), .B(n406), .Z(n573) );
  XOR2_X1 U329 ( .A(KEYINPUT38), .B(n442), .Z(n488) );
  AND2_X1 U330 ( .A1(G231GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U331 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n292) );
  XOR2_X1 U332 ( .A(n320), .B(n319), .Z(n293) );
  XOR2_X1 U333 ( .A(n431), .B(KEYINPUT31), .Z(n294) );
  XNOR2_X1 U334 ( .A(G99GAT), .B(G85GAT), .ZN(n298) );
  NOR2_X1 U335 ( .A1(n452), .A2(n451), .ZN(n453) );
  XNOR2_X1 U336 ( .A(n399), .B(n291), .ZN(n400) );
  INV_X1 U337 ( .A(KEYINPUT94), .ZN(n390) );
  XNOR2_X1 U338 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U339 ( .A(n441), .B(n440), .ZN(n569) );
  INV_X1 U340 ( .A(KEYINPUT120), .ZN(n465) );
  XNOR2_X1 U341 ( .A(n465), .B(G169GAT), .ZN(n466) );
  XNOR2_X1 U342 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U343 ( .A(n467), .B(n466), .ZN(G1348GAT) );
  XNOR2_X1 U344 ( .A(n446), .B(n445), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(G29GAT), .B(G43GAT), .Z(n296) );
  XNOR2_X1 U346 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n424) );
  XNOR2_X1 U348 ( .A(G36GAT), .B(G190GAT), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n297), .B(G218GAT), .ZN(n353) );
  XNOR2_X1 U350 ( .A(n424), .B(n353), .ZN(n311) );
  XOR2_X1 U351 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n300) );
  XOR2_X1 U352 ( .A(G50GAT), .B(G162GAT), .Z(n333) );
  XNOR2_X1 U353 ( .A(n298), .B(KEYINPUT72), .ZN(n431) );
  XNOR2_X1 U354 ( .A(n333), .B(n431), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U356 ( .A(G92GAT), .B(KEYINPUT74), .Z(n302) );
  NAND2_X1 U357 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U359 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U360 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n306) );
  XNOR2_X1 U361 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U363 ( .A(G134GAT), .B(n307), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n558) );
  XNOR2_X1 U366 ( .A(KEYINPUT36), .B(n558), .ZN(n578) );
  XNOR2_X1 U367 ( .A(G127GAT), .B(KEYINPUT81), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n312), .B(KEYINPUT82), .ZN(n313) );
  XOR2_X1 U369 ( .A(n313), .B(KEYINPUT0), .Z(n315) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(G134GAT), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n373) );
  XOR2_X1 U372 ( .A(KEYINPUT83), .B(G99GAT), .Z(n317) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(G190GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n320) );
  XNOR2_X1 U375 ( .A(G15GAT), .B(KEYINPUT65), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n292), .B(n318), .ZN(n319) );
  XOR2_X1 U377 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XOR2_X1 U378 ( .A(G183GAT), .B(G176GAT), .Z(n322) );
  NAND2_X1 U379 ( .A1(G227GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n434), .B(n323), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n293), .B(n324), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n373), .B(n325), .ZN(n329) );
  XOR2_X1 U384 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n327) );
  XNOR2_X1 U385 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U387 ( .A(G169GAT), .B(n328), .ZN(n359) );
  XNOR2_X2 U388 ( .A(n329), .B(n359), .ZN(n518) );
  XOR2_X1 U389 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n331) );
  XNOR2_X1 U390 ( .A(G218GAT), .B(KEYINPUT23), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U392 ( .A(n333), .B(n332), .Z(n335) );
  NAND2_X1 U393 ( .A1(G228GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n349) );
  XOR2_X1 U395 ( .A(KEYINPUT88), .B(KEYINPUT24), .Z(n337) );
  XNOR2_X1 U396 ( .A(G22GAT), .B(KEYINPUT86), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n340) );
  XOR2_X1 U398 ( .A(G211GAT), .B(KEYINPUT89), .Z(n339) );
  XNOR2_X1 U399 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n356) );
  XOR2_X1 U401 ( .A(n340), .B(n356), .Z(n347) );
  XOR2_X1 U402 ( .A(G148GAT), .B(G106GAT), .Z(n342) );
  XNOR2_X1 U403 ( .A(G204GAT), .B(G78GAT), .ZN(n341) );
  XNOR2_X1 U404 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U405 ( .A(KEYINPUT71), .B(n343), .Z(n439) );
  XOR2_X1 U406 ( .A(G155GAT), .B(KEYINPUT2), .Z(n345) );
  XNOR2_X1 U407 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n369) );
  XNOR2_X1 U409 ( .A(n439), .B(n369), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U411 ( .A(n349), .B(n348), .Z(n462) );
  XNOR2_X1 U412 ( .A(n462), .B(KEYINPUT28), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n350), .B(KEYINPUT66), .ZN(n481) );
  XOR2_X1 U414 ( .A(G8GAT), .B(G183GAT), .Z(n394) );
  XOR2_X1 U415 ( .A(n394), .B(G204GAT), .Z(n352) );
  NAND2_X1 U416 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U418 ( .A(n354), .B(n353), .Z(n358) );
  XNOR2_X1 U419 ( .A(G176GAT), .B(G92GAT), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n355), .B(G64GAT), .ZN(n429) );
  XNOR2_X1 U421 ( .A(n356), .B(n429), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n508) );
  XNOR2_X1 U424 ( .A(n508), .B(KEYINPUT27), .ZN(n380) );
  XOR2_X1 U425 ( .A(KEYINPUT91), .B(KEYINPUT4), .Z(n362) );
  XNOR2_X1 U426 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n362), .B(n361), .ZN(n377) );
  XOR2_X1 U428 ( .A(G85GAT), .B(G162GAT), .Z(n364) );
  XNOR2_X1 U429 ( .A(G29GAT), .B(G148GAT), .ZN(n363) );
  XNOR2_X1 U430 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U431 ( .A(KEYINPUT90), .B(G57GAT), .Z(n366) );
  XNOR2_X1 U432 ( .A(G1GAT), .B(G120GAT), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U434 ( .A(n368), .B(n367), .Z(n375) );
  XOR2_X1 U435 ( .A(n369), .B(KEYINPUT6), .Z(n371) );
  NAND2_X1 U436 ( .A1(G225GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U440 ( .A(n377), .B(n376), .Z(n505) );
  NAND2_X1 U441 ( .A1(n380), .A2(n505), .ZN(n378) );
  XOR2_X1 U442 ( .A(KEYINPUT92), .B(n378), .Z(n533) );
  NAND2_X1 U443 ( .A1(n481), .A2(n533), .ZN(n520) );
  NOR2_X1 U444 ( .A1(n518), .A2(n520), .ZN(n389) );
  NOR2_X1 U445 ( .A1(n462), .A2(n518), .ZN(n379) );
  XOR2_X1 U446 ( .A(KEYINPUT26), .B(n379), .Z(n563) );
  INV_X1 U447 ( .A(n380), .ZN(n381) );
  NOR2_X1 U448 ( .A1(n563), .A2(n381), .ZN(n385) );
  NAND2_X1 U449 ( .A1(n508), .A2(n518), .ZN(n382) );
  NAND2_X1 U450 ( .A1(n462), .A2(n382), .ZN(n383) );
  XNOR2_X1 U451 ( .A(n383), .B(KEYINPUT25), .ZN(n384) );
  NOR2_X1 U452 ( .A1(n505), .A2(n386), .ZN(n387) );
  XOR2_X1 U453 ( .A(KEYINPUT93), .B(n387), .Z(n388) );
  NOR2_X1 U454 ( .A1(n389), .A2(n388), .ZN(n391) );
  XOR2_X1 U455 ( .A(G64GAT), .B(G211GAT), .Z(n393) );
  XNOR2_X1 U456 ( .A(G127GAT), .B(G71GAT), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n407) );
  XOR2_X1 U458 ( .A(KEYINPUT13), .B(G57GAT), .Z(n430) );
  XOR2_X1 U459 ( .A(n394), .B(n430), .Z(n396) );
  XNOR2_X1 U460 ( .A(G78GAT), .B(G155GAT), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n401) );
  XOR2_X1 U462 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n398) );
  XNOR2_X1 U463 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U465 ( .A(n402), .B(KEYINPUT77), .Z(n405) );
  XNOR2_X1 U466 ( .A(G22GAT), .B(G15GAT), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n403), .B(G1GAT), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n411), .B(KEYINPUT14), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n406) );
  NAND2_X1 U470 ( .A1(n471), .A2(n573), .ZN(n408) );
  XOR2_X1 U471 ( .A(KEYINPUT99), .B(n408), .Z(n409) );
  XOR2_X1 U472 ( .A(KEYINPUT37), .B(n410), .Z(n502) );
  XOR2_X1 U473 ( .A(G36GAT), .B(n411), .Z(n413) );
  NAND2_X1 U474 ( .A1(G229GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U476 ( .A(n414), .B(G50GAT), .Z(n422) );
  XOR2_X1 U477 ( .A(G113GAT), .B(G197GAT), .Z(n416) );
  XNOR2_X1 U478 ( .A(G169GAT), .B(G141GAT), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U480 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n418) );
  XNOR2_X1 U481 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U485 ( .A(n423), .B(G8GAT), .Z(n426) );
  XNOR2_X1 U486 ( .A(n424), .B(KEYINPUT29), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n565) );
  XOR2_X1 U488 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n428) );
  XNOR2_X1 U489 ( .A(KEYINPUT73), .B(KEYINPUT70), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n438) );
  XOR2_X1 U491 ( .A(n430), .B(n429), .Z(n436) );
  NAND2_X1 U492 ( .A1(G230GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n294), .B(n432), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n441) );
  INV_X1 U497 ( .A(n439), .ZN(n440) );
  NOR2_X1 U498 ( .A1(n565), .A2(n569), .ZN(n472) );
  NAND2_X1 U499 ( .A1(n502), .A2(n472), .ZN(n442) );
  NAND2_X1 U500 ( .A1(n488), .A2(n518), .ZN(n446) );
  XOR2_X1 U501 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n444) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n443) );
  XNOR2_X1 U503 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n457) );
  NOR2_X1 U504 ( .A1(n573), .A2(n578), .ZN(n447) );
  XOR2_X1 U505 ( .A(KEYINPUT45), .B(n447), .Z(n448) );
  NOR2_X1 U506 ( .A1(n569), .A2(n448), .ZN(n449) );
  NAND2_X1 U507 ( .A1(n449), .A2(n565), .ZN(n455) );
  NAND2_X1 U508 ( .A1(n558), .A2(n573), .ZN(n452) );
  XNOR2_X1 U509 ( .A(KEYINPUT41), .B(n569), .ZN(n539) );
  NOR2_X1 U510 ( .A1(n565), .A2(n539), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n450), .B(KEYINPUT46), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n453), .B(KEYINPUT47), .ZN(n454) );
  NAND2_X1 U513 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n534), .A2(n508), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT54), .B(KEYINPUT119), .Z(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n460) );
  NOR2_X1 U517 ( .A1(n460), .A2(n505), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(KEYINPUT64), .ZN(n562) );
  NAND2_X1 U519 ( .A1(n462), .A2(n562), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n463), .B(KEYINPUT55), .ZN(n464) );
  NAND2_X1 U521 ( .A1(n464), .A2(n518), .ZN(n557) );
  NOR2_X1 U522 ( .A1(n565), .A2(n557), .ZN(n467) );
  XOR2_X1 U523 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n474) );
  XOR2_X1 U524 ( .A(KEYINPUT80), .B(KEYINPUT16), .Z(n469) );
  INV_X1 U525 ( .A(n573), .ZN(n544) );
  NAND2_X1 U526 ( .A1(n558), .A2(n544), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n470) );
  AND2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n491) );
  AND2_X1 U529 ( .A1(n472), .A2(n491), .ZN(n482) );
  NAND2_X1 U530 ( .A1(n482), .A2(n505), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U533 ( .A1(n482), .A2(n508), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(KEYINPUT96), .ZN(n477) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n479) );
  NAND2_X1 U537 ( .A1(n482), .A2(n518), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U539 ( .A(G15GAT), .B(n480), .Z(G1326GAT) );
  INV_X1 U540 ( .A(n481), .ZN(n512) );
  NAND2_X1 U541 ( .A1(n512), .A2(n482), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n483), .B(KEYINPUT98), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(n484), .ZN(G1327GAT) );
  XOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT39), .Z(n486) );
  NAND2_X1 U545 ( .A1(n505), .A2(n488), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NAND2_X1 U547 ( .A1(n488), .A2(n508), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U549 ( .A1(n512), .A2(n488), .ZN(n489) );
  XNOR2_X1 U550 ( .A(G50GAT), .B(n489), .ZN(G1331GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n494) );
  INV_X1 U552 ( .A(n565), .ZN(n537) );
  XOR2_X1 U553 ( .A(n539), .B(KEYINPUT103), .Z(n550) );
  NOR2_X1 U554 ( .A1(n537), .A2(n550), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n490), .B(KEYINPUT104), .ZN(n503) );
  NAND2_X1 U556 ( .A1(n503), .A2(n491), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n492), .B(KEYINPUT105), .ZN(n499) );
  NAND2_X1 U558 ( .A1(n499), .A2(n505), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U560 ( .A(G57GAT), .B(n495), .Z(G1332GAT) );
  NAND2_X1 U561 ( .A1(n499), .A2(n508), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n496), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U563 ( .A1(n518), .A2(n499), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n497), .B(KEYINPUT106), .ZN(n498) );
  XNOR2_X1 U565 ( .A(G71GAT), .B(n498), .ZN(G1334GAT) );
  XOR2_X1 U566 ( .A(G78GAT), .B(KEYINPUT43), .Z(n501) );
  NAND2_X1 U567 ( .A1(n499), .A2(n512), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n501), .B(n500), .ZN(G1335GAT) );
  XNOR2_X1 U569 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n504), .B(KEYINPUT107), .ZN(n513) );
  NAND2_X1 U572 ( .A1(n505), .A2(n513), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1336GAT) );
  NAND2_X1 U574 ( .A1(n513), .A2(n508), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U576 ( .A(G99GAT), .B(KEYINPUT109), .Z(n511) );
  NAND2_X1 U577 ( .A1(n513), .A2(n518), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1338GAT) );
  XNOR2_X1 U579 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n517) );
  XOR2_X1 U580 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n515) );
  NAND2_X1 U581 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1339GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n534), .ZN(n519) );
  NOR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n525) );
  NAND2_X1 U586 ( .A1(n537), .A2(n525), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(G113GAT), .ZN(G1340GAT) );
  INV_X1 U588 ( .A(n525), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n550), .A2(n530), .ZN(n523) );
  XNOR2_X1 U590 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U592 ( .A(G120GAT), .B(n524), .Z(G1341GAT) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n527) );
  NAND2_X1 U595 ( .A1(n525), .A2(n544), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(G1342GAT) );
  NOR2_X1 U598 ( .A1(n558), .A2(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(G1343GAT) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n535), .A2(n563), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT116), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n537), .A2(n545), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n538), .ZN(G1344GAT) );
  INV_X1 U606 ( .A(n545), .ZN(n547) );
  NOR2_X1 U607 ( .A1(n547), .A2(n539), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n541) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n558), .A2(n547), .ZN(n548) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(n548), .Z(n549) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n549), .ZN(G1347GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n557), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n552) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(KEYINPUT121), .B(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  NOR2_X1 U623 ( .A1(n573), .A2(n557), .ZN(n556) );
  XOR2_X1 U624 ( .A(G183GAT), .B(n556), .Z(G1350GAT) );
  XNOR2_X1 U625 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(n561), .ZN(G1351GAT) );
  INV_X1 U628 ( .A(n562), .ZN(n564) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n570) );
  INV_X1 U630 ( .A(n570), .ZN(n577) );
  NOR2_X1 U631 ( .A1(n565), .A2(n577), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n577), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G218GAT), .B(n581), .Z(G1355GAT) );
endmodule

