

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  XNOR2_X1 U324 ( .A(n373), .B(n335), .ZN(n336) );
  XNOR2_X1 U325 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n448) );
  XNOR2_X1 U327 ( .A(n341), .B(n340), .ZN(n347) );
  XOR2_X1 U328 ( .A(n333), .B(n332), .Z(n530) );
  AND2_X1 U329 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U330 ( .A(n338), .B(n337), .Z(n293) );
  XOR2_X1 U331 ( .A(G211GAT), .B(KEYINPUT21), .Z(n294) );
  XNOR2_X1 U332 ( .A(n422), .B(n292), .ZN(n335) );
  INV_X1 U333 ( .A(KEYINPUT77), .ZN(n398) );
  XNOR2_X1 U334 ( .A(n339), .B(n293), .ZN(n340) );
  INV_X1 U335 ( .A(KEYINPUT100), .ZN(n471) );
  XNOR2_X1 U336 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U337 ( .A(n466), .B(n465), .ZN(n572) );
  NOR2_X1 U338 ( .A1(n587), .A2(n492), .ZN(n493) );
  XNOR2_X1 U339 ( .A(n472), .B(n471), .ZN(n479) );
  XNOR2_X1 U340 ( .A(n425), .B(n400), .ZN(n404) );
  NAND2_X1 U341 ( .A1(n479), .A2(n478), .ZN(n490) );
  XNOR2_X1 U342 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U343 ( .A(n412), .B(n411), .ZN(n579) );
  NOR2_X1 U344 ( .A1(n539), .A2(n452), .ZN(n570) );
  XOR2_X1 U345 ( .A(KEYINPUT38), .B(n495), .Z(n505) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n295), .B(G29GAT), .ZN(n296) );
  XOR2_X1 U348 ( .A(n296), .B(KEYINPUT72), .Z(n298) );
  XNOR2_X1 U349 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n297) );
  XOR2_X1 U350 ( .A(n298), .B(n297), .Z(n426) );
  XOR2_X1 U351 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n300) );
  XNOR2_X1 U352 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n314) );
  XOR2_X1 U354 ( .A(G197GAT), .B(G22GAT), .Z(n302) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(G141GAT), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U357 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n304) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(G8GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U360 ( .A(n306), .B(n305), .Z(n312) );
  XNOR2_X1 U361 ( .A(G15GAT), .B(G1GAT), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n307), .B(KEYINPUT73), .ZN(n383) );
  XOR2_X1 U363 ( .A(G50GAT), .B(n383), .Z(n309) );
  NAND2_X1 U364 ( .A1(G229GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U366 ( .A(G36GAT), .B(n310), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U368 ( .A(n314), .B(n313), .Z(n315) );
  XOR2_X1 U369 ( .A(n426), .B(n315), .Z(n555) );
  XOR2_X1 U370 ( .A(G120GAT), .B(G71GAT), .Z(n408) );
  XOR2_X1 U371 ( .A(G99GAT), .B(G190GAT), .Z(n317) );
  XNOR2_X1 U372 ( .A(G43GAT), .B(G15GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U374 ( .A(n408), .B(n318), .Z(n320) );
  NAND2_X1 U375 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U377 ( .A(KEYINPUT88), .B(KEYINPUT65), .Z(n322) );
  XNOR2_X1 U378 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U380 ( .A(n324), .B(n323), .Z(n333) );
  XNOR2_X1 U381 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n325), .B(KEYINPUT87), .ZN(n326) );
  XOR2_X1 U383 ( .A(n326), .B(KEYINPUT18), .Z(n328) );
  XNOR2_X1 U384 ( .A(G169GAT), .B(G183GAT), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n374) );
  XOR2_X1 U386 ( .A(KEYINPUT0), .B(G134GAT), .Z(n330) );
  XNOR2_X1 U387 ( .A(KEYINPUT86), .B(G127GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U389 ( .A(G113GAT), .B(n331), .Z(n351) );
  XNOR2_X1 U390 ( .A(n374), .B(n351), .ZN(n332) );
  INV_X1 U391 ( .A(n530), .ZN(n539) );
  XNOR2_X1 U392 ( .A(G197GAT), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n294), .B(n334), .ZN(n373) );
  XOR2_X1 U394 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XOR2_X1 U395 ( .A(n336), .B(G204GAT), .Z(n341) );
  XNOR2_X1 U396 ( .A(G22GAT), .B(G155GAT), .ZN(n391) );
  XOR2_X1 U397 ( .A(n391), .B(KEYINPUT89), .Z(n339) );
  XOR2_X1 U398 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n338) );
  XNOR2_X1 U399 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n337) );
  XOR2_X1 U400 ( .A(G78GAT), .B(G148GAT), .Z(n343) );
  XNOR2_X1 U401 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n406) );
  XOR2_X1 U403 ( .A(KEYINPUT3), .B(KEYINPUT90), .Z(n345) );
  XNOR2_X1 U404 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n406), .B(n350), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n475) );
  XOR2_X1 U408 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n349) );
  XNOR2_X1 U409 ( .A(G57GAT), .B(KEYINPUT94), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n355) );
  XOR2_X1 U411 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n353) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n367) );
  NAND2_X1 U415 ( .A1(G225GAT), .A2(G233GAT), .ZN(n361) );
  XOR2_X1 U416 ( .A(G85GAT), .B(G155GAT), .Z(n357) );
  XNOR2_X1 U417 ( .A(G120GAT), .B(G148GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n359) );
  XOR2_X1 U419 ( .A(G29GAT), .B(G162GAT), .Z(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U422 ( .A(KEYINPUT95), .B(KEYINPUT4), .Z(n363) );
  XNOR2_X1 U423 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n524) );
  XOR2_X1 U427 ( .A(G64GAT), .B(G92GAT), .Z(n369) );
  XNOR2_X1 U428 ( .A(G176GAT), .B(G204GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n405) );
  XOR2_X1 U430 ( .A(G36GAT), .B(G190GAT), .Z(n421) );
  XOR2_X1 U431 ( .A(n405), .B(n421), .Z(n371) );
  NAND2_X1 U432 ( .A1(G226GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U434 ( .A(G8GAT), .B(KEYINPUT83), .Z(n386) );
  XOR2_X1 U435 ( .A(n372), .B(n386), .Z(n376) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U437 ( .A(n376), .B(n375), .Z(n527) );
  XOR2_X1 U438 ( .A(KEYINPUT121), .B(n527), .Z(n447) );
  XOR2_X1 U439 ( .A(G64GAT), .B(G71GAT), .Z(n378) );
  XNOR2_X1 U440 ( .A(G183GAT), .B(G127GAT), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U442 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n380) );
  XNOR2_X1 U443 ( .A(KEYINPUT85), .B(KEYINPUT12), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n395) );
  XOR2_X1 U446 ( .A(n383), .B(KEYINPUT14), .Z(n385) );
  NAND2_X1 U447 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U449 ( .A(G57GAT), .B(KEYINPUT13), .Z(n407) );
  XOR2_X1 U450 ( .A(n407), .B(n386), .Z(n388) );
  XNOR2_X1 U451 ( .A(G78GAT), .B(G211GAT), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n393) );
  INV_X1 U454 ( .A(n391), .ZN(n392) );
  XOR2_X1 U455 ( .A(n393), .B(n392), .Z(n394) );
  XOR2_X1 U456 ( .A(n395), .B(n394), .Z(n491) );
  INV_X1 U457 ( .A(n491), .ZN(n582) );
  XOR2_X1 U458 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n397) );
  XNOR2_X1 U459 ( .A(G99GAT), .B(G85GAT), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n425) );
  NAND2_X1 U461 ( .A1(G230GAT), .A2(G233GAT), .ZN(n399) );
  XOR2_X1 U462 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n402) );
  XNOR2_X1 U463 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U465 ( .A(n404), .B(n403), .Z(n412) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U468 ( .A(n579), .B(KEYINPUT41), .Z(n565) );
  AND2_X1 U469 ( .A1(n555), .A2(n565), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n413), .B(KEYINPUT46), .ZN(n414) );
  NOR2_X1 U471 ( .A1(n582), .A2(n414), .ZN(n435) );
  XOR2_X1 U472 ( .A(KEYINPUT80), .B(KEYINPUT9), .Z(n416) );
  XNOR2_X1 U473 ( .A(KEYINPUT79), .B(KEYINPUT64), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U475 ( .A(G92GAT), .B(KEYINPUT10), .Z(n418) );
  XNOR2_X1 U476 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n434) );
  XOR2_X1 U479 ( .A(KEYINPUT81), .B(n421), .Z(n424) );
  XNOR2_X1 U480 ( .A(n422), .B(G218GAT), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U482 ( .A(n425), .B(KEYINPUT82), .Z(n428) );
  XOR2_X1 U483 ( .A(n426), .B(G134GAT), .Z(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U485 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U486 ( .A1(G232GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n438) );
  INV_X1 U489 ( .A(n438), .ZN(n456) );
  NAND2_X1 U490 ( .A1(n435), .A2(n456), .ZN(n437) );
  XOR2_X1 U491 ( .A(KEYINPUT114), .B(KEYINPUT47), .Z(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n445) );
  INV_X1 U493 ( .A(KEYINPUT36), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n489) );
  NOR2_X1 U495 ( .A1(n489), .A2(n491), .ZN(n441) );
  XOR2_X1 U496 ( .A(KEYINPUT45), .B(KEYINPUT115), .Z(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n443) );
  NOR2_X1 U498 ( .A1(n579), .A2(n555), .ZN(n442) );
  NAND2_X1 U499 ( .A1(n443), .A2(n442), .ZN(n444) );
  NAND2_X1 U500 ( .A1(n445), .A2(n444), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n446), .B(KEYINPUT48), .ZN(n552) );
  NAND2_X1 U502 ( .A1(n447), .A2(n552), .ZN(n449) );
  NOR2_X1 U503 ( .A1(n524), .A2(n450), .ZN(n574) );
  AND2_X1 U504 ( .A1(n475), .A2(n574), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  NAND2_X1 U506 ( .A1(n555), .A2(n570), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n453), .B(KEYINPUT124), .ZN(n455) );
  XOR2_X1 U508 ( .A(G169GAT), .B(KEYINPUT123), .Z(n454) );
  XNOR2_X1 U509 ( .A(n455), .B(n454), .ZN(G1348GAT) );
  INV_X1 U510 ( .A(G190GAT), .ZN(n460) );
  INV_X1 U511 ( .A(n456), .ZN(n562) );
  NAND2_X1 U512 ( .A1(n570), .A2(n562), .ZN(n458) );
  XOR2_X1 U513 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n457) );
  XNOR2_X1 U514 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  INV_X1 U516 ( .A(n555), .ZN(n575) );
  NOR2_X1 U517 ( .A1(n575), .A2(n579), .ZN(n494) );
  INV_X1 U518 ( .A(n494), .ZN(n481) );
  NOR2_X1 U519 ( .A1(n491), .A2(n562), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT16), .ZN(n480) );
  NAND2_X1 U521 ( .A1(n530), .A2(n527), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n462), .A2(n475), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n463), .B(KEYINPUT25), .ZN(n464) );
  XOR2_X1 U524 ( .A(KEYINPUT99), .B(n464), .Z(n469) );
  NOR2_X1 U525 ( .A1(n475), .A2(n530), .ZN(n466) );
  XNOR2_X1 U526 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n465) );
  XOR2_X1 U527 ( .A(n527), .B(KEYINPUT27), .Z(n473) );
  NOR2_X1 U528 ( .A1(n572), .A2(n473), .ZN(n467) );
  XNOR2_X1 U529 ( .A(KEYINPUT98), .B(n467), .ZN(n468) );
  NOR2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U531 ( .A1(n524), .A2(n470), .ZN(n472) );
  INV_X1 U532 ( .A(n473), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n524), .A2(n474), .ZN(n551) );
  XOR2_X1 U534 ( .A(n475), .B(KEYINPUT66), .Z(n476) );
  XNOR2_X1 U535 ( .A(KEYINPUT28), .B(n476), .ZN(n532) );
  NOR2_X1 U536 ( .A1(n551), .A2(n532), .ZN(n537) );
  XNOR2_X1 U537 ( .A(n537), .B(KEYINPUT96), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n477), .A2(n539), .ZN(n478) );
  NAND2_X1 U539 ( .A1(n480), .A2(n490), .ZN(n508) );
  NOR2_X1 U540 ( .A1(n481), .A2(n508), .ZN(n487) );
  NAND2_X1 U541 ( .A1(n487), .A2(n524), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n482), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U544 ( .A1(n527), .A2(n487), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U547 ( .A1(n487), .A2(n530), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U549 ( .A1(n532), .A2(n487), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  BUF_X1 U551 ( .A(n489), .Z(n587) );
  NAND2_X1 U552 ( .A1(n491), .A2(n490), .ZN(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n493), .Z(n521) );
  NAND2_X1 U554 ( .A1(n521), .A2(n494), .ZN(n495) );
  NAND2_X1 U555 ( .A1(n505), .A2(n524), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n500) );
  NAND2_X1 U560 ( .A1(n505), .A2(n527), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n503) );
  NAND2_X1 U564 ( .A1(n505), .A2(n530), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U566 ( .A(G43GAT), .B(n504), .Z(G1330GAT) );
  NAND2_X1 U567 ( .A1(n505), .A2(n532), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U569 ( .A1(n565), .A2(n575), .ZN(n507) );
  XOR2_X1 U570 ( .A(n507), .B(KEYINPUT105), .Z(n520) );
  NOR2_X1 U571 ( .A1(n520), .A2(n508), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n524), .A2(n517), .ZN(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(n509), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n512) );
  NAND2_X1 U576 ( .A1(n517), .A2(n527), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n515) );
  NAND2_X1 U580 ( .A1(n517), .A2(n530), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G71GAT), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U584 ( .A1(n517), .A2(n532), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  INV_X1 U586 ( .A(n520), .ZN(n522) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U588 ( .A(KEYINPUT110), .B(n523), .Z(n533) );
  NAND2_X1 U589 ( .A1(n533), .A2(n524), .ZN(n525) );
  XOR2_X1 U590 ( .A(KEYINPUT111), .B(n525), .Z(n526) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(KEYINPUT112), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n533), .A2(n530), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n535) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n552), .A2(n537), .ZN(n538) );
  NOR2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n555), .A2(n547), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U606 ( .A1(n547), .A2(n565), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n544) );
  NAND2_X1 U610 ( .A1(n547), .A2(n582), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U614 ( .A1(n547), .A2(n562), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n550), .ZN(G1343GAT) );
  NOR2_X1 U617 ( .A1(n572), .A2(n551), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT119), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n555), .A2(n561), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n558) );
  NAND2_X1 U623 ( .A1(n561), .A2(n565), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n582), .A2(n561), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT120), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n570), .A2(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT57), .Z(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n582), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U638 ( .A(n572), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n575), .A2(n586), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  INV_X1 U645 ( .A(n586), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n583), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .Z(n585) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

