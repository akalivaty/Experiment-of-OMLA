//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  INV_X1    g001(.A(G71gat), .ZN(new_n203));
  INV_X1    g002(.A(G78gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT9), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G71gat), .B(G78gat), .Z(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT21), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G231gat), .A2(G233gat), .ZN(new_n213));
  XOR2_X1   g012(.A(new_n213), .B(KEYINPUT96), .Z(new_n214));
  XNOR2_X1  g013(.A(new_n212), .B(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G127gat), .B(G155gat), .Z(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G183gat), .B(G211gat), .Z(new_n218));
  XOR2_X1   g017(.A(new_n217), .B(new_n218), .Z(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT93), .A2(G1gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT16), .B1(KEYINPUT93), .B2(G1gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT94), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n220), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(G1gat), .B2(new_n221), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n227), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n228), .B(new_n229), .C1(new_n208), .C2(new_n209), .ZN(new_n230));
  XOR2_X1   g029(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n219), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G43gat), .B(G50gat), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n234), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n235));
  OR3_X1    g034(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n235), .B(new_n238), .C1(KEYINPUT15), .C2(new_n234), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT92), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n241), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n236), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G29gat), .ZN(new_n245));
  INV_X1    g044(.A(G36gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT15), .A3(new_n234), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n240), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n240), .A2(KEYINPUT17), .A3(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT7), .ZN(new_n254));
  NAND2_X1  g053(.A1(G99gat), .A2(G106gat), .ZN(new_n255));
  INV_X1    g054(.A(G85gat), .ZN(new_n256));
  INV_X1    g055(.A(G92gat), .ZN(new_n257));
  AOI22_X1  g056(.A1(KEYINPUT8), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G99gat), .B(G106gat), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n254), .B(new_n258), .C1(KEYINPUT99), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(KEYINPUT99), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n251), .A2(new_n252), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  AND2_X1   g063(.A1(G232gat), .A2(G233gat), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n249), .A2(new_n264), .B1(KEYINPUT41), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT100), .ZN(new_n268));
  XOR2_X1   g067(.A(G134gat), .B(G162gat), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n265), .A2(KEYINPUT41), .ZN(new_n271));
  XNOR2_X1  g070(.A(G190gat), .B(G218gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n273), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n233), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n262), .B(new_n208), .Z(new_n278));
  INV_X1    g077(.A(KEYINPUT10), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OR3_X1    g079(.A1(new_n262), .A2(new_n279), .A3(new_n208), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G230gat), .A2(G233gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n278), .B2(new_n283), .ZN(new_n285));
  XNOR2_X1  g084(.A(G120gat), .B(G148gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G176gat), .B(G204gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n289), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n228), .A2(new_n229), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(new_n249), .B2(new_n250), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n296), .A2(new_n252), .B1(new_n295), .B2(new_n249), .ZN(new_n297));
  NAND2_X1  g096(.A1(G229gat), .A2(G233gat), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT18), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n249), .B(new_n295), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n298), .B(KEYINPUT13), .Z(new_n301));
  AOI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(KEYINPUT18), .A3(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G113gat), .B(G141gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G169gat), .B(G197gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n309), .B(KEYINPUT12), .Z(new_n310));
  OR2_X1    g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT95), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n304), .A2(new_n310), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n304), .A2(KEYINPUT95), .A3(new_n310), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n277), .A2(new_n294), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G8gat), .B(G36gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(G64gat), .B(G92gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n319), .B(new_n320), .Z(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT65), .ZN(new_n323));
  INV_X1    g122(.A(G183gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT64), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n328), .A2(new_n329), .B1(KEYINPUT24), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(KEYINPUT24), .B2(new_n332), .ZN(new_n334));
  INV_X1    g133(.A(G169gat), .ZN(new_n335));
  INV_X1    g134(.A(G176gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT23), .B1(new_n335), .B2(new_n336), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n334), .A2(new_n343), .A3(KEYINPUT25), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n343), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT25), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n347), .A3(new_n330), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT67), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n325), .A2(KEYINPUT27), .A3(new_n326), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353));
  AOI21_X1  g152(.A(G190gat), .B1(new_n353), .B2(G183gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(KEYINPUT66), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT66), .B1(new_n352), .B2(new_n354), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n351), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n352), .A2(new_n354), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n362), .A2(KEYINPUT67), .A3(new_n356), .A4(new_n355), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n354), .B(KEYINPUT28), .C1(new_n353), .C2(G183gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n337), .A2(KEYINPUT26), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT68), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n341), .B1(KEYINPUT26), .B2(new_n337), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n368), .A2(new_n369), .B1(G183gat), .B2(G190gat), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n366), .B1(new_n365), .B2(new_n370), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n350), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G226gat), .ZN(new_n374));
  INV_X1    g173(.A(G233gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT29), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT22), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT77), .B(G218gat), .ZN(new_n380));
  INV_X1    g179(.A(G211gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(KEYINPUT76), .A2(G197gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(KEYINPUT76), .A2(G197gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(G204gat), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n384), .ZN(new_n386));
  INV_X1    g185(.A(G204gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G211gat), .B(G218gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(KEYINPUT78), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(KEYINPUT78), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n393), .A2(new_n382), .A3(new_n385), .A4(new_n388), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n365), .A2(new_n370), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n350), .A3(new_n376), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n378), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(KEYINPUT69), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n350), .A3(new_n376), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n397), .A2(new_n350), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n377), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n396), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n322), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n376), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n373), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n395), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n378), .A2(new_n396), .A3(new_n398), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n321), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n410), .A2(new_n414), .A3(new_n411), .A4(new_n321), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(G57gat), .B(G85gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT5), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT81), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G127gat), .B(G134gat), .Z(new_n426));
  XNOR2_X1  g225(.A(G113gat), .B(G120gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(KEYINPUT1), .B2(new_n427), .ZN(new_n428));
  XOR2_X1   g227(.A(G113gat), .B(G120gat), .Z(new_n429));
  INV_X1    g228(.A(KEYINPUT1), .ZN(new_n430));
  XNOR2_X1  g229(.A(G127gat), .B(G134gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G148gat), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT80), .B1(new_n434), .B2(G141gat), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436));
  INV_X1    g235(.A(G141gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(G148gat), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n435), .B(new_n438), .C1(new_n437), .C2(G148gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440));
  OR2_X1    g239(.A1(G155gat), .A2(G162gat), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(KEYINPUT2), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G141gat), .B(G148gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n440), .B(new_n441), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT3), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n433), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n443), .A2(new_n446), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(KEYINPUT3), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n422), .B(new_n425), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n428), .A2(new_n432), .A3(KEYINPUT70), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT70), .B1(new_n428), .B2(new_n432), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n447), .B(new_n454), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT4), .B1(new_n450), .B2(new_n433), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n453), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n453), .A3(new_n458), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n452), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n450), .A2(new_n433), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n446), .A2(new_n443), .B1(new_n428), .B2(new_n432), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n424), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g265(.A(new_n433), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT4), .B1(new_n447), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n456), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n428), .A2(new_n432), .A3(KEYINPUT70), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n450), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n468), .B1(new_n471), .B2(KEYINPUT4), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n467), .B1(KEYINPUT3), .B2(new_n450), .ZN(new_n473));
  INV_X1    g272(.A(new_n451), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n424), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n466), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n421), .B1(new_n462), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT84), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n472), .A2(new_n475), .ZN(new_n480));
  INV_X1    g279(.A(new_n466), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n457), .A2(new_n453), .A3(new_n458), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n422), .B(new_n475), .C1(new_n483), .C2(new_n459), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n420), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT6), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n482), .A2(new_n484), .A3(new_n420), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n477), .A2(new_n489), .A3(new_n478), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n416), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT31), .B(G50gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT86), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(G106gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT29), .B1(new_n447), .B2(new_n448), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(new_n395), .ZN(new_n500));
  NAND2_X1  g299(.A1(G228gat), .A2(G233gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT3), .B1(new_n395), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n447), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT29), .B1(new_n389), .B2(new_n390), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n382), .A2(new_n391), .A3(new_n385), .A4(new_n388), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n447), .B1(new_n509), .B2(new_n448), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n506), .B(new_n501), .C1(new_n510), .C2(new_n500), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT3), .B1(new_n507), .B2(new_n508), .ZN(new_n513));
  OAI22_X1  g312(.A1(new_n513), .A2(new_n447), .B1(new_n499), .B2(new_n395), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n506), .B1(new_n514), .B2(new_n501), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n505), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G22gat), .ZN(new_n517));
  INV_X1    g316(.A(G22gat), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n518), .B(new_n505), .C1(new_n512), .C2(new_n515), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n517), .A2(new_n519), .A3(new_n204), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n204), .B1(new_n517), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n498), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n517), .A2(new_n519), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G78gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n517), .A2(new_n519), .A3(new_n204), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(new_n497), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n494), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n479), .A2(new_n487), .A3(new_n490), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT37), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n410), .A2(new_n530), .A3(new_n411), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n409), .A2(new_n396), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n378), .A2(new_n395), .A3(new_n398), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT37), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n321), .A2(KEYINPUT38), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n529), .A2(new_n536), .A3(new_n412), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT37), .B1(new_n399), .B2(new_n406), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT88), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n539), .A3(new_n322), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n530), .B1(new_n410), .B2(new_n411), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT88), .B1(new_n541), .B2(new_n321), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n542), .A3(new_n531), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n537), .B1(new_n543), .B2(KEYINPUT38), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT40), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n473), .A2(new_n474), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(new_n483), .B2(new_n459), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT39), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n424), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n420), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n463), .A2(new_n464), .A3(new_n424), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n551), .A2(KEYINPUT87), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n548), .B1(new_n551), .B2(KEYINPUT87), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n547), .B2(new_n424), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n545), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n547), .A2(new_n424), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n552), .A3(new_n553), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n558), .A2(KEYINPUT40), .A3(new_n420), .A4(new_n549), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n556), .A2(new_n559), .A3(new_n477), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(new_n413), .A3(new_n415), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(new_n526), .A3(new_n522), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n528), .B1(new_n544), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n565));
  NAND2_X1  g364(.A1(G227gat), .A2(G233gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n567));
  INV_X1    g366(.A(new_n350), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n400), .B2(new_n401), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n455), .A2(new_n456), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n567), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n373), .A2(KEYINPUT72), .A3(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT71), .B1(new_n373), .B2(new_n570), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT71), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n402), .A2(new_n576), .A3(new_n571), .A4(new_n350), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n566), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT73), .B(KEYINPUT33), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n565), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n572), .A2(new_n573), .B1(new_n575), .B2(new_n577), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT32), .B1(new_n583), .B2(new_n566), .ZN(new_n584));
  XNOR2_X1  g383(.A(G15gat), .B(G43gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT75), .ZN(new_n586));
  XOR2_X1   g385(.A(G71gat), .B(G99gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  OAI211_X1 g387(.A(KEYINPUT74), .B(new_n580), .C1(new_n583), .C2(new_n566), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n582), .A2(new_n584), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n583), .A2(new_n591), .A3(new_n566), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n583), .B2(new_n566), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n588), .A2(new_n581), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n584), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n590), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n594), .B1(new_n590), .B2(new_n596), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n590), .A2(new_n596), .ZN(new_n601));
  INV_X1    g400(.A(new_n594), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n590), .A2(new_n594), .A3(new_n596), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT36), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n564), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n597), .A2(new_n598), .A3(new_n527), .ZN(new_n607));
  INV_X1    g406(.A(new_n416), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT89), .B(KEYINPUT35), .Z(new_n609));
  NOR3_X1   g408(.A1(new_n608), .A2(new_n529), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n494), .ZN(new_n612));
  INV_X1    g411(.A(new_n527), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n603), .A2(new_n604), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT35), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n318), .B1(new_n606), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n493), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g419(.A(KEYINPUT16), .B(G8gat), .Z(new_n621));
  AND3_X1   g420(.A1(new_n617), .A2(new_n608), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n220), .B1(new_n617), .B2(new_n608), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT42), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(KEYINPUT42), .B2(new_n622), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT101), .ZN(G1325gat));
  INV_X1    g425(.A(G15gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n597), .A2(new_n598), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n617), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n599), .B1(new_n597), .B2(new_n598), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n603), .A2(KEYINPUT36), .A3(new_n604), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n617), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n629), .B1(new_n634), .B2(new_n627), .ZN(G1326gat));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n527), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT43), .B(G22gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1327gat));
  INV_X1    g437(.A(new_n276), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n639), .B1(new_n616), .B2(new_n606), .ZN(new_n640));
  INV_X1    g439(.A(new_n233), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n641), .A2(new_n293), .A3(new_n316), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n643), .A2(G29gat), .A3(new_n493), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT45), .Z(new_n645));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT102), .B1(new_n632), .B2(new_n564), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648));
  AOI211_X1 g447(.A(new_n648), .B(new_n563), .C1(new_n630), .C2(new_n631), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n616), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n276), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n607), .A2(new_n610), .B1(new_n614), .B2(KEYINPUT35), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n563), .B1(new_n630), .B2(new_n631), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n276), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n650), .A2(new_n653), .B1(new_n656), .B2(KEYINPUT44), .ZN(new_n657));
  INV_X1    g456(.A(new_n642), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n646), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n606), .A2(new_n648), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(KEYINPUT102), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n652), .B1(new_n662), .B2(new_n616), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n640), .A2(new_n651), .ZN(new_n664));
  OAI211_X1 g463(.A(KEYINPUT103), .B(new_n642), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT104), .B1(new_n666), .B2(new_n493), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G29gat), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n666), .A2(KEYINPUT104), .A3(new_n493), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n645), .B1(new_n668), .B2(new_n669), .ZN(G1328gat));
  OAI21_X1  g469(.A(G36gat), .B1(new_n666), .B2(new_n416), .ZN(new_n671));
  AND2_X1   g470(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n672));
  NOR2_X1   g471(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n643), .A2(G36gat), .A3(new_n416), .ZN(new_n675));
  MUX2_X1   g474(.A(new_n674), .B(new_n672), .S(new_n675), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(G1329gat));
  OAI21_X1  g476(.A(new_n642), .B1(new_n663), .B2(new_n664), .ZN(new_n678));
  OAI21_X1  g477(.A(G43gat), .B1(new_n678), .B2(new_n632), .ZN(new_n679));
  INV_X1    g478(.A(new_n628), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n643), .A2(G43gat), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(KEYINPUT47), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n659), .A2(new_n633), .A3(new_n665), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G43gat), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n681), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n685), .A2(KEYINPUT106), .A3(G43gat), .ZN(new_n689));
  AOI211_X1 g488(.A(new_n684), .B(KEYINPUT47), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(new_n689), .A3(new_n682), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT107), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n683), .B1(new_n690), .B2(new_n694), .ZN(G1330gat));
  NOR2_X1   g494(.A1(new_n613), .A2(G50gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n643), .B2(KEYINPUT110), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n697), .B1(KEYINPUT110), .B2(new_n643), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G50gat), .B1(new_n678), .B2(new_n613), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n659), .A2(new_n527), .A3(new_n665), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n703), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT109), .B1(new_n703), .B2(G50gat), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n704), .A2(new_n705), .A3(new_n698), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n702), .B1(new_n706), .B2(new_n707), .ZN(G1331gat));
  AND4_X1   g507(.A1(new_n277), .A2(new_n650), .A3(new_n293), .A4(new_n316), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n618), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT111), .B(G57gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1332gat));
  AOI21_X1  g511(.A(new_n416), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT112), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1333gat));
  AOI21_X1  g516(.A(new_n203), .B1(new_n709), .B2(new_n633), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n680), .A2(G71gat), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n709), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g520(.A1(new_n709), .A2(new_n527), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g522(.A(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n233), .A2(new_n276), .A3(new_n316), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(KEYINPUT51), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n729), .A2(KEYINPUT113), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT113), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n731), .A2(new_n732), .A3(new_n294), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n256), .A3(new_n618), .ZN(new_n734));
  NOR4_X1   g533(.A1(new_n657), .A2(new_n641), .A3(new_n294), .A4(new_n317), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(new_n618), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n256), .B2(new_n736), .ZN(G1336gat));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n608), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G92gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n729), .A2(new_n730), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n294), .A2(G92gat), .A3(new_n416), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT52), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n727), .A2(KEYINPUT114), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n727), .A2(KEYINPUT114), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n728), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n744), .A2(KEYINPUT115), .A3(new_n728), .A4(new_n745), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n730), .A3(new_n749), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n750), .A2(new_n741), .B1(G92gat), .B2(new_n738), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n743), .B1(new_n751), .B2(new_n752), .ZN(G1337gat));
  INV_X1    g552(.A(G99gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n733), .A2(new_n754), .A3(new_n628), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n735), .A2(new_n633), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n754), .B2(new_n756), .ZN(G1338gat));
  NAND2_X1  g556(.A1(new_n735), .A2(new_n527), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G106gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n613), .A2(new_n294), .A3(G106gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n740), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n762));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n750), .A2(new_n760), .B1(G106gat), .B2(new_n758), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(G1339gat));
  OR2_X1    g565(.A1(new_n282), .A2(new_n283), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n767), .A2(KEYINPUT54), .A3(new_n284), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT117), .ZN(new_n769));
  INV_X1    g568(.A(new_n284), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n288), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n290), .B1(new_n773), .B2(KEYINPUT55), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n772), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n297), .A2(new_n298), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n300), .A2(new_n301), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n309), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n311), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n778), .A2(new_n276), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n317), .A2(new_n774), .A3(new_n777), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n293), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n276), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n233), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n277), .A2(new_n294), .A3(new_n316), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(new_n607), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n608), .A2(new_n493), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n317), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n293), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n641), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g598(.A1(new_n639), .A2(new_n608), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n493), .A2(G134gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n790), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT56), .Z(new_n803));
  OAI21_X1  g602(.A(G134gat), .B1(new_n792), .B2(new_n639), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1343gat));
  NOR2_X1   g604(.A1(new_n778), .A2(KEYINPUT120), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n774), .A2(new_n777), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n317), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n785), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n783), .B1(new_n810), .B2(new_n639), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n788), .B1(new_n811), .B2(new_n641), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n613), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n789), .A2(new_n527), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n817), .A3(new_n813), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n613), .B1(new_n787), .B2(new_n788), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT119), .B1(new_n819), .B2(KEYINPUT57), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n632), .A2(new_n791), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n317), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G141gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT121), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n816), .A2(new_n822), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n437), .A3(new_n317), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(new_n829), .A3(KEYINPUT58), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n825), .B(new_n828), .C1(KEYINPUT121), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1344gat));
  NAND3_X1  g632(.A1(new_n827), .A2(new_n434), .A3(new_n293), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n821), .A2(new_n823), .ZN(new_n835));
  AOI211_X1 g634(.A(KEYINPUT59), .B(new_n434), .C1(new_n835), .C2(new_n293), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n812), .A2(KEYINPUT122), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n812), .A2(KEYINPUT122), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n613), .A2(KEYINPUT57), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n816), .A2(KEYINPUT57), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n841), .A2(new_n293), .A3(new_n823), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n837), .B1(new_n843), .B2(G148gat), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n834), .B1(new_n836), .B2(new_n844), .ZN(G1345gat));
  AOI21_X1  g644(.A(G155gat), .B1(new_n827), .B2(new_n641), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n641), .A2(G155gat), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT123), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n835), .B2(new_n848), .ZN(G1346gat));
  NAND2_X1  g648(.A1(new_n835), .A2(new_n276), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G162gat), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n493), .A2(G162gat), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n819), .A2(new_n632), .A3(new_n800), .A4(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT124), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(G1347gat));
  NOR2_X1   g654(.A1(new_n618), .A2(new_n416), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n790), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n316), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(new_n335), .ZN(G1348gat));
  NOR2_X1   g658(.A1(new_n857), .A2(new_n294), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(new_n336), .ZN(G1349gat));
  INV_X1    g660(.A(new_n857), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n324), .A2(KEYINPUT27), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n353), .A2(G183gat), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n862), .B(new_n641), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n328), .B1(new_n857), .B2(new_n233), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT60), .Z(G1350gat));
  NOR2_X1   g667(.A1(new_n857), .A2(new_n639), .ZN(new_n869));
  NAND2_X1  g668(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT61), .B(G190gat), .Z(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n869), .B2(new_n872), .ZN(G1351gat));
  AND2_X1   g672(.A1(new_n841), .A2(new_n842), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n632), .A2(new_n856), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n317), .A3(new_n876), .ZN(new_n877));
  XOR2_X1   g676(.A(KEYINPUT125), .B(G197gat), .Z(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n816), .A2(new_n875), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n317), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1352gat));
  NAND3_X1  g682(.A1(new_n874), .A2(new_n293), .A3(new_n876), .ZN(new_n884));
  XOR2_X1   g683(.A(KEYINPUT126), .B(G204gat), .Z(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n294), .A2(new_n885), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT62), .Z(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(G1353gat));
  NAND3_X1  g689(.A1(new_n881), .A2(new_n381), .A3(new_n641), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n841), .A2(new_n641), .A3(new_n842), .A4(new_n876), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n892), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT63), .B1(new_n892), .B2(G211gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(G1354gat));
  AOI21_X1  g694(.A(G218gat), .B1(new_n881), .B2(new_n276), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT127), .Z(new_n897));
  AND2_X1   g696(.A1(new_n874), .A2(new_n876), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n639), .A2(new_n380), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(G1355gat));
endmodule


