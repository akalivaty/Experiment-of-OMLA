//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n468), .B(KEYINPUT68), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n462), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(KEYINPUT70), .A3(G101), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n464), .B1(new_n462), .B2(KEYINPUT69), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n474), .A2(new_n475), .B1(new_n479), .B2(G137), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n470), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n479), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n484), .B2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n476), .A2(new_n478), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI211_X1 g064(.A(KEYINPUT71), .B(new_n484), .C1(new_n476), .C2(new_n478), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n486), .B1(new_n492), .B2(G124), .ZN(G162));
  NAND2_X1  g068(.A1(new_n471), .A2(G102), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n488), .B2(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n497), .B2(new_n484), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n463), .A2(new_n465), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n484), .A2(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n499), .A2(KEYINPUT4), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n500), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT3), .B1(new_n477), .B2(G2104), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n506), .B2(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n505), .A2(new_n508), .A3(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n498), .B1(new_n507), .B2(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n515), .A2(G62), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n516), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n517), .A2(new_n519), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n513), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n512), .A2(new_n514), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n530), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G168));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n521), .A2(new_n541), .B1(new_n523), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n515), .A2(G64), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n516), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n521), .A2(new_n548), .B1(new_n523), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n537), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n550), .B1(KEYINPUT74), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n554), .A2(KEYINPUT74), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT75), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n556), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n531), .A2(G53), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n569), .A2(new_n570), .B1(new_n538), .B2(G91), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n571), .B1(new_n570), .B2(new_n569), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT76), .B(G65), .Z(new_n573));
  AOI22_X1  g148(.A1(new_n515), .A2(new_n573), .B1(G78), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n516), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  NAND4_X1  g155(.A1(new_n517), .A2(new_n519), .A3(G49), .A4(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT77), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n538), .A2(G87), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n537), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n538), .A2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n531), .A2(G48), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n516), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT78), .ZN(new_n595));
  XOR2_X1   g170(.A(KEYINPUT79), .B(G47), .Z(new_n596));
  AOI22_X1  g171(.A1(new_n538), .A2(G85), .B1(new_n531), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n594), .A2(KEYINPUT78), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n537), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(new_n531), .B2(G54), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT80), .Z(new_n607));
  NAND2_X1  g182(.A1(new_n538), .A2(G92), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT10), .Z(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n602), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n602), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n576), .B2(G868), .ZN(G297));
  XOR2_X1   g190(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n563), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n611), .A2(new_n617), .A3(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(G282));
  INV_X1    g199(.A(new_n622), .ZN(G323));
  NAND2_X1  g200(.A1(new_n479), .A2(G135), .ZN(new_n626));
  NOR2_X1   g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(new_n484), .B2(G111), .ZN(new_n628));
  INV_X1    g203(.A(G123), .ZN(new_n629));
  OAI221_X1 g204(.A(new_n626), .B1(new_n627), .B2(new_n628), .C1(new_n491), .C2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT84), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n466), .A2(new_n471), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT13), .B(G2100), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n632), .A2(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT14), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n644), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(G14), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n658), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n658), .B(KEYINPUT17), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n663), .B(new_n660), .C1(new_n657), .C2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n657), .A3(new_n659), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT86), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT87), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n676), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  AOI211_X1 g255(.A(new_n678), .B(new_n680), .C1(new_n673), .C2(new_n677), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT88), .B(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  INV_X1    g261(.A(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G19), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n563), .B2(new_n690), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(G1341), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(G1341), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(G20), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT23), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n576), .B2(new_n690), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1956), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(G164), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G27), .B2(new_n699), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n698), .B1(new_n443), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n443), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n693), .A2(new_n694), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n699), .A2(G26), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(new_n484), .B2(G116), .ZN(new_n707));
  INV_X1    g282(.A(G104), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n484), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT91), .Z(new_n710));
  INV_X1    g285(.A(G140), .ZN(new_n711));
  INV_X1    g286(.A(new_n479), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G128), .B2(new_n492), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n706), .B1(new_n714), .B2(new_n699), .ZN(new_n715));
  INV_X1    g290(.A(G2067), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G5), .A2(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n719), .B(new_n720), .C1(G301), .C2(new_n690), .ZN(new_n721));
  INV_X1    g296(.A(G1961), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g298(.A1(KEYINPUT24), .A2(G34), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n699), .B1(KEYINPUT24), .B2(G34), .ZN(new_n725));
  OAI22_X1  g300(.A1(G160), .A2(new_n699), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT93), .B(G2084), .Z(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(new_n484), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n732), .B(new_n734), .C1(G139), .C2(new_n479), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n699), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n699), .B2(G33), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(new_n442), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n717), .A2(new_n723), .A3(new_n729), .A4(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G168), .A2(new_n690), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n690), .B2(G21), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n726), .A2(new_n728), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n745), .B1(new_n722), .B2(new_n721), .C1(new_n442), .C2(new_n737), .ZN(new_n746));
  INV_X1    g321(.A(G28), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n747), .B2(KEYINPUT30), .ZN(new_n749));
  OR2_X1    g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  NAND2_X1  g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n752), .B1(new_n699), .B2(new_n630), .C1(new_n741), .C2(new_n742), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n739), .A2(new_n746), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n699), .A2(G35), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT96), .Z(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G162), .B2(new_n699), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G2090), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n690), .A2(G4), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n611), .B2(new_n690), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1348), .ZN(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  INV_X1    g339(.A(new_n758), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n699), .A2(G32), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT26), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n770), .A2(new_n771), .B1(G105), .B2(new_n471), .ZN(new_n772));
  INV_X1    g347(.A(G141), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n712), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n492), .B2(G129), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n767), .B1(new_n776), .B2(new_n699), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT27), .B(G1996), .Z(new_n778));
  XOR2_X1   g353(.A(new_n777), .B(new_n778), .Z(new_n779));
  NAND4_X1  g354(.A1(new_n754), .A2(new_n760), .A3(new_n766), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n690), .B1(G290), .B2(KEYINPUT90), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(KEYINPUT90), .B2(G290), .ZN(new_n782));
  INV_X1    g357(.A(G24), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(G16), .B2(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(G1986), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(G1986), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(new_n484), .B2(G107), .ZN(new_n787));
  INV_X1    g362(.A(G95), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n484), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G131), .B2(new_n479), .ZN(new_n790));
  INV_X1    g365(.A(G119), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n491), .B2(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G25), .B(new_n792), .S(G29), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT89), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT35), .B(G1991), .Z(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n785), .A2(new_n786), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n690), .A2(G6), .ZN(new_n799));
  INV_X1    g374(.A(G305), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n690), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(G1981), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(G1981), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n690), .A2(G23), .ZN(new_n805));
  INV_X1    g380(.A(G288), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n690), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT33), .B(G1976), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n690), .A2(G22), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G166), .B2(new_n690), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G1971), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n808), .A2(new_n809), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n809), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n807), .A2(new_n815), .B1(new_n811), .B2(G1971), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n803), .A2(new_n804), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT34), .ZN(new_n818));
  OR3_X1    g393(.A1(new_n798), .A2(new_n818), .A3(KEYINPUT36), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT36), .B1(new_n798), .B2(new_n818), .ZN(new_n820));
  AOI211_X1 g395(.A(new_n704), .B(new_n780), .C1(new_n819), .C2(new_n820), .ZN(G311));
  XNOR2_X1  g396(.A(G311), .B(KEYINPUT98), .ZN(G150));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n537), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G651), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n538), .A2(G93), .B1(new_n531), .B2(G55), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n826), .A2(new_n827), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n562), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n559), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n611), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT100), .Z(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n833), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  NOR2_X1   g423(.A1(new_n735), .A2(new_n775), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n776), .B2(new_n735), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n635), .Z(new_n851));
  AOI21_X1  g426(.A(new_n500), .B1(new_n476), .B2(new_n478), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT4), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT72), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n466), .A2(new_n853), .A3(new_n502), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n509), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n494), .ZN(new_n857));
  OAI21_X1  g432(.A(G126), .B1(new_n503), .B2(new_n504), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n495), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n857), .B1(new_n859), .B2(G2105), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n714), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n479), .A2(G142), .ZN(new_n863));
  NOR2_X1   g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(new_n484), .B2(G118), .ZN(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  OAI221_X1 g441(.A(new_n863), .B1(new_n864), .B2(new_n865), .C1(new_n491), .C2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n792), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n862), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n851), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(G162), .B(G160), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n630), .ZN(new_n872));
  AOI21_X1  g447(.A(G37), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(new_n870), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g450(.A1(new_n833), .A2(new_n619), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n611), .A2(new_n617), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n837), .B(new_n877), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n610), .A2(new_n576), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n610), .A2(new_n576), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n610), .A2(KEYINPUT101), .A3(new_n576), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n882), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n879), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n878), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n883), .A2(new_n879), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n891), .B1(new_n893), .B2(new_n878), .ZN(new_n894));
  XOR2_X1   g469(.A(G166), .B(KEYINPUT102), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n600), .ZN(new_n896));
  XNOR2_X1  g471(.A(G288), .B(G305), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT42), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n894), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n876), .B1(new_n900), .B2(new_n619), .ZN(G295));
  OAI21_X1  g476(.A(new_n876), .B1(new_n900), .B2(new_n619), .ZN(G331));
  XOR2_X1   g477(.A(G171), .B(G168), .Z(new_n903));
  NAND3_X1  g478(.A1(new_n834), .A2(new_n836), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  INV_X1    g480(.A(new_n903), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n832), .B1(new_n558), .B2(new_n561), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(new_n835), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n837), .A2(KEYINPUT103), .A3(new_n906), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n893), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n904), .A2(new_n908), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n890), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n911), .B2(new_n912), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n898), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n898), .B1(new_n914), .B2(new_n917), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT43), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n911), .A2(new_n912), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n923), .A2(new_n919), .A3(new_n913), .A4(new_n916), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n909), .A2(new_n910), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n881), .A2(new_n884), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n927), .A2(new_n888), .B1(new_n886), .B2(new_n892), .ZN(new_n928));
  OAI22_X1  g503(.A1(new_n926), .A2(new_n928), .B1(new_n893), .B2(new_n915), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n898), .ZN(new_n930));
  AND4_X1   g505(.A1(KEYINPUT43), .A2(new_n924), .A3(new_n925), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n922), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n920), .B2(new_n921), .ZN(new_n934));
  AND4_X1   g509(.A1(new_n933), .A2(new_n924), .A3(new_n925), .A4(new_n930), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n936), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g512(.A(G1384), .B1(new_n856), .B2(new_n860), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(KEYINPUT45), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n470), .A2(new_n480), .A3(G40), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n714), .B(G2067), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n775), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n941), .A2(G1996), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT46), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n947), .A2(KEYINPUT46), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT47), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n945), .A2(G1996), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n942), .B1(new_n944), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n947), .A2(new_n776), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(KEYINPUT105), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n954), .A2(KEYINPUT105), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n957), .B(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n792), .A2(new_n796), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n792), .A2(new_n796), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n942), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(G290), .A2(new_n941), .A3(G1986), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT48), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n951), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n961), .B(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n959), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n714), .A2(new_n716), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n941), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n972));
  NAND3_X1  g547(.A1(G303), .A2(G8), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(G166), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n979), .B(new_n980), .C1(G164), .C2(G1384), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT107), .B1(new_n938), .B2(KEYINPUT45), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n981), .B(new_n940), .C1(new_n982), .C2(new_n939), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n940), .B1(new_n938), .B2(new_n984), .ZN(new_n985));
  AOI211_X1 g560(.A(KEYINPUT50), .B(G1384), .C1(new_n856), .C2(new_n860), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n983), .A2(new_n813), .B1(new_n987), .B2(new_n764), .ZN(new_n988));
  OAI21_X1  g563(.A(G8), .B1(new_n988), .B2(KEYINPUT114), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(new_n813), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n764), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n990), .A2(KEYINPUT114), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n978), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n975), .B1(new_n940), .B2(new_n938), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n806), .A2(G1976), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT52), .ZN(new_n997));
  NAND2_X1  g572(.A1(G305), .A2(G1981), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n589), .A2(new_n590), .A3(new_n1000), .A4(new_n591), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G305), .A2(KEYINPUT111), .A3(G1981), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT49), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n994), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n940), .A2(new_n938), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(G288), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1009), .A2(G8), .A3(new_n995), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n997), .B(new_n1008), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n861), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n986), .ZN(new_n1021));
  INV_X1    g596(.A(new_n940), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n938), .A2(new_n984), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(KEYINPUT108), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(new_n1024), .A3(new_n764), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n975), .B1(new_n990), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1016), .B1(new_n1026), .B2(new_n977), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n939), .A2(new_n1022), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n980), .B(G1384), .C1(new_n856), .C2(new_n860), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT115), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1018), .B2(new_n980), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n742), .ZN(new_n1034));
  INV_X1    g609(.A(G2084), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1021), .A2(new_n1024), .A3(new_n1035), .ZN(new_n1036));
  AOI211_X1 g611(.A(new_n975), .B(G286), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n993), .A2(new_n1027), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT63), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(KEYINPUT116), .A3(new_n1039), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1026), .A2(new_n977), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1027), .A2(new_n1044), .A3(KEYINPUT63), .A4(new_n1037), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(new_n975), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G168), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1034), .A2(G286), .A3(new_n1036), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1034), .A2(G168), .A3(new_n1036), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT51), .B1(new_n1054), .B2(G8), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT62), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1052), .ZN(new_n1057));
  AOI21_X1  g632(.A(G286), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1048), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1047), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT62), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1056), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n983), .B2(G2078), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT108), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1020), .B1(new_n938), .B2(new_n984), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1067), .B(new_n940), .C1(new_n1068), .C2(new_n1023), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n722), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1065), .A2(G2078), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .A4(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(KEYINPUT124), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT124), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1066), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AND4_X1   g651(.A1(G171), .A2(new_n993), .A3(new_n1076), .A4(new_n1027), .ZN(new_n1077));
  NOR2_X1   g652(.A1(G288), .A2(G1976), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1008), .A2(new_n1078), .B1(new_n1000), .B2(new_n800), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1079), .A2(KEYINPUT112), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n994), .B1(new_n1079), .B2(KEYINPUT112), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1026), .A2(new_n977), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1080), .A2(new_n1081), .B1(new_n1082), .B2(new_n1016), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT113), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n1085));
  OAI221_X1 g660(.A(new_n1085), .B1(new_n1082), .B2(new_n1016), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1064), .A2(new_n1077), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n576), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n1092), .B(KEYINPUT118), .Z(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT119), .B1(new_n983), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1018), .A2(new_n980), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(KEYINPUT107), .B2(new_n1029), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1022), .B1(new_n939), .B2(new_n979), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1093), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n987), .A2(G1956), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1091), .A2(new_n1094), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1348), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1009), .A2(G2067), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n611), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1094), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1091), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1103), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1109), .A2(KEYINPUT122), .A3(KEYINPUT61), .A4(new_n1102), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G1348), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1069), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1105), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT123), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1117), .A2(new_n1123), .A3(KEYINPUT60), .A4(new_n1118), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1120), .A2(new_n611), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(G1341), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1009), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n983), .B2(G1996), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n562), .A2(KEYINPUT121), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1125), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT61), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1120), .A2(new_n1124), .B1(new_n611), .B2(new_n1122), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1110), .B1(new_n1115), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1066), .A2(G301), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1075), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1073), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1029), .A2(new_n1065), .A3(G2078), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1069), .A2(new_n722), .B1(new_n1145), .B2(new_n1028), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1066), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(G171), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT54), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1141), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1142), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(KEYINPUT125), .A3(KEYINPUT54), .A4(new_n1148), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1143), .A2(new_n1073), .ZN(new_n1156));
  AOI21_X1  g731(.A(G301), .B1(new_n1156), .B2(new_n1066), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1151), .A2(new_n1146), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1155), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AND4_X1   g734(.A1(new_n1027), .A2(new_n1059), .A3(new_n1061), .A4(new_n993), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1154), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1046), .B(new_n1087), .C1(new_n1140), .C2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n600), .B(new_n687), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n963), .B1(new_n942), .B2(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1162), .A2(KEYINPUT126), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT126), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n971), .B1(new_n1165), .B2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g742(.A1(new_n654), .A2(G319), .ZN(new_n1169));
  NOR3_X1   g743(.A1(G227), .A2(G229), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n874), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g745(.A1(new_n936), .A2(new_n1171), .ZN(G308));
  OR2_X1    g746(.A1(new_n936), .A2(new_n1171), .ZN(G225));
endmodule


