//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n225), .B1(new_n202), .B2(new_n226), .C1(new_n203), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT64), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G45), .ZN(new_n249));
  AOI21_X1  g0049(.A(G1), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n252), .A3(G274), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n253), .B1(new_n221), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n226), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n227), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G107), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(new_n257), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n252), .B1(new_n263), .B2(KEYINPUT66), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n256), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G169), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G179), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT67), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n274), .A2(new_n207), .A3(G13), .A4(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n216), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n207), .A2(G20), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n276), .A2(G77), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  XOR2_X1   g0081(.A(KEYINPUT15), .B(G87), .Z(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G20), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n282), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n281), .B1(G77), .B2(new_n276), .C1(new_n290), .C2(new_n279), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n269), .A2(new_n271), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(G190), .B2(new_n266), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n267), .A2(G200), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n252), .ZN(new_n297));
  INV_X1    g0097(.A(G222), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n257), .B1(new_n298), .B2(G1698), .ZN(new_n299));
  OR2_X1    g0099(.A1(KEYINPUT65), .A2(G223), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT65), .A2(G223), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n259), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n297), .B1(G77), .B2(new_n257), .C1(new_n299), .C2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n255), .ZN(new_n304));
  INV_X1    g0104(.A(G274), .ZN(new_n305));
  AND2_X1   g0105(.A1(G1), .A2(G13), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n251), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n304), .A2(G226), .B1(new_n250), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G179), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n287), .A2(new_n284), .B1(G150), .B2(new_n288), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n204), .A2(G20), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n279), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n272), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n278), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G50), .A3(new_n280), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(G50), .B2(new_n272), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n309), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n311), .B(new_n319), .C1(G169), .C2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n296), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT74), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n288), .A2(G50), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n288), .A2(KEYINPUT72), .A3(G50), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n208), .A2(G33), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n329), .A2(new_n220), .B1(new_n208), .B2(G68), .ZN(new_n330));
  OAI211_X1 g0130(.A(KEYINPUT11), .B(new_n278), .C1(new_n328), .C2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT11), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n326), .B2(new_n327), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n279), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n273), .A2(KEYINPUT12), .A3(new_n203), .A4(new_n275), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT12), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n272), .B2(G68), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n331), .A2(new_n334), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n276), .A2(G68), .A3(new_n279), .A4(new_n280), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT73), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n339), .B(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n323), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n339), .B(KEYINPUT73), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n335), .A2(new_n337), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n333), .A2(new_n279), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(KEYINPUT11), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n343), .A2(new_n346), .A3(KEYINPUT74), .A4(new_n334), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT71), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n252), .A2(G238), .A3(new_n254), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n253), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n253), .A2(new_n352), .A3(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G97), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(KEYINPUT70), .A2(G33), .A3(G97), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n226), .A2(G1698), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G226), .B2(G1698), .ZN(new_n363));
  AND2_X1   g0163(.A1(KEYINPUT3), .A2(G33), .ZN(new_n364));
  NOR2_X1   g0164(.A1(KEYINPUT3), .A2(G33), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n361), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n297), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n350), .B1(new_n356), .B2(new_n368), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n253), .A2(new_n352), .A3(new_n351), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n350), .B(new_n368), .C1(new_n370), .C2(new_n353), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n349), .B(G169), .C1(new_n369), .C2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n368), .B1(new_n370), .B2(new_n353), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT13), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(G179), .A3(new_n371), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n371), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n349), .B1(new_n378), .B2(G169), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n348), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n342), .A2(new_n347), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(G200), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n381), .B(new_n382), .C1(new_n383), .C2(new_n378), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n320), .A2(G190), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n319), .A2(KEYINPUT9), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n314), .A2(new_n318), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT9), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT69), .B(new_n386), .C1(new_n387), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT10), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n386), .B1(new_n387), .B2(new_n390), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n309), .A2(G200), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT68), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n391), .B(new_n392), .C1(new_n394), .C2(new_n396), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n322), .A2(new_n385), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n316), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n287), .A2(new_n280), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(KEYINPUT76), .B2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n402), .A2(KEYINPUT76), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n403), .A2(new_n404), .B1(new_n315), .B2(new_n286), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  OR2_X1    g0207(.A1(KEYINPUT3), .A2(G33), .ZN(new_n408));
  NAND2_X1  g0208(.A1(KEYINPUT3), .A2(G33), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n208), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n408), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n409), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n203), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT75), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n202), .A2(new_n203), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G58), .A2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(G20), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n288), .A2(G159), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(new_n414), .C2(KEYINPUT75), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n407), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n420), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n279), .B1(new_n424), .B2(KEYINPUT16), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n406), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  MUX2_X1   g0226(.A(G223), .B(G226), .S(G1698), .Z(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n257), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT77), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n297), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n427), .A2(new_n257), .B1(G33), .B2(G87), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT77), .B1(new_n433), .B2(new_n252), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n253), .B1(new_n226), .B2(new_n255), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(G179), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n433), .A2(new_n252), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n268), .B1(new_n438), .B2(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT18), .B1(new_n426), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n424), .A2(KEYINPUT16), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n278), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT7), .B1(new_n366), .B2(new_n208), .ZN(new_n444));
  INV_X1    g0244(.A(new_n413), .ZN(new_n445));
  OAI21_X1  g0245(.A(G68), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT75), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n423), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT16), .B1(new_n448), .B2(new_n415), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n405), .B1(new_n443), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n440), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n441), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n435), .A2(G190), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n432), .A2(new_n434), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n438), .A2(new_n435), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(G200), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n405), .C1(new_n443), .C2(new_n449), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT17), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n400), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n207), .B(G45), .C1(new_n248), .C2(KEYINPUT5), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n248), .A2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n307), .A3(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G257), .B(new_n252), .C1(new_n464), .C2(new_n466), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n221), .A2(G1698), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n364), .B2(new_n365), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  OAI211_X1 g0275(.A(G250), .B(G1698), .C1(new_n364), .C2(new_n365), .ZN(new_n476));
  INV_X1    g0276(.A(new_n473), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n477), .B(new_n471), .C1(new_n365), .C2(new_n364), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n474), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  AOI211_X1 g0279(.A(KEYINPUT80), .B(new_n470), .C1(new_n297), .C2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT80), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n297), .ZN(new_n482));
  INV_X1    g0282(.A(new_n470), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n480), .A2(new_n484), .A3(new_n383), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n483), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G200), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  AND2_X1   g0288(.A1(G97), .A2(G107), .ZN(new_n489));
  NOR2_X1   g0289(.A1(G97), .A2(G107), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n262), .A2(KEYINPUT6), .A3(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n493), .A2(G20), .B1(G77), .B2(new_n288), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n262), .B1(new_n412), .B2(new_n413), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(KEYINPUT78), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT78), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n497), .B(new_n262), .C1(new_n412), .C2(new_n413), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n278), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n272), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n207), .A2(G33), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n316), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n500), .B1(new_n503), .B2(G97), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n487), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n463), .B1(new_n485), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n486), .A2(KEYINPUT80), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n482), .A2(new_n481), .A3(new_n483), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(G190), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n504), .ZN(new_n510));
  OAI21_X1  g0310(.A(G107), .B1(new_n444), .B2(new_n445), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n497), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n495), .A2(KEYINPUT78), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(new_n494), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n510), .B1(new_n514), .B2(new_n278), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n509), .A2(new_n515), .A3(KEYINPUT81), .A4(new_n487), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n486), .A2(G179), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n507), .A2(new_n508), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(new_n268), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n499), .A2(new_n504), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n506), .A2(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n262), .A2(KEYINPUT23), .A3(G20), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT23), .B1(new_n262), .B2(G20), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n522), .A2(new_n523), .B1(G20), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n208), .B(G87), .C1(new_n364), .C2(new_n365), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT22), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n257), .A2(new_n528), .A3(new_n208), .A4(G87), .ZN(new_n529));
  AOI211_X1 g0329(.A(KEYINPUT24), .B(new_n525), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n529), .ZN(new_n532));
  INV_X1    g0332(.A(new_n525), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n278), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n315), .A2(new_n262), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n536), .A2(KEYINPUT25), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(KEYINPUT25), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(new_n262), .C2(new_n502), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G250), .B(new_n259), .C1(new_n364), .C2(new_n365), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  AND2_X1   g0342(.A1(G257), .A2(G1698), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n364), .B2(new_n365), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n297), .ZN(new_n546));
  OAI211_X1 g0346(.A(G264), .B(new_n252), .C1(new_n464), .C2(new_n466), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(new_n468), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n546), .A2(new_n547), .A3(G190), .A4(new_n468), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n535), .A2(new_n540), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(new_n531), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n539), .B1(new_n553), .B2(new_n278), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n548), .A2(new_n268), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n546), .A2(new_n547), .A3(new_n270), .A4(new_n468), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n551), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n223), .B1(new_n249), .B2(G1), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n207), .A2(new_n305), .A3(G45), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n252), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n524), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G238), .A2(G1698), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n221), .B2(G1698), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n562), .B1(new_n564), .B2(new_n257), .ZN(new_n565));
  OAI211_X1 g0365(.A(G190), .B(new_n561), .C1(new_n565), .C2(new_n252), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n227), .A2(new_n259), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n221), .A2(G1698), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(new_n364), .C2(new_n365), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n524), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n297), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n573), .A2(KEYINPUT84), .A3(G190), .A4(new_n561), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n276), .A2(new_n282), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n359), .A2(KEYINPUT19), .A3(new_n360), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n208), .ZN(new_n578));
  INV_X1    g0378(.A(G97), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n222), .A2(new_n579), .A3(new_n262), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT82), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT82), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n582), .A2(new_n222), .A3(new_n579), .A4(new_n262), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n257), .A2(new_n586), .A3(new_n208), .A4(G68), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n284), .A2(G97), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n208), .B(G68), .C1(new_n364), .C2(new_n365), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT83), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n585), .A2(new_n587), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n576), .B1(new_n593), .B2(new_n278), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n503), .A2(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n573), .A2(new_n561), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G200), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n575), .A2(new_n594), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n592), .A2(new_n587), .A3(new_n590), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n208), .A2(new_n577), .B1(new_n581), .B2(new_n583), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n278), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n576), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n503), .A2(new_n282), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(G169), .B1(new_n573), .B2(new_n561), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n252), .B1(new_n571), .B2(new_n524), .ZN(new_n606));
  INV_X1    g0406(.A(new_n561), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n606), .A2(new_n607), .A3(G179), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n598), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n276), .A2(G116), .A3(new_n279), .A4(new_n501), .ZN(new_n612));
  INV_X1    g0412(.A(G116), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n273), .A2(new_n613), .A3(new_n275), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n277), .A2(new_n216), .B1(G20), .B2(new_n613), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n475), .B(new_n208), .C1(G33), .C2(new_n579), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT20), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n615), .A2(KEYINPUT20), .A3(new_n616), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n612), .B(new_n614), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n259), .A2(G257), .ZN(new_n620));
  NAND2_X1  g0420(.A1(G264), .A2(G1698), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n257), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G303), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n366), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n624), .A3(new_n297), .ZN(new_n625));
  OAI211_X1 g0425(.A(G270), .B(new_n252), .C1(new_n464), .C2(new_n466), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n468), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n619), .A2(G169), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT85), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n619), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n627), .A2(G200), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n625), .A2(G190), .A3(new_n468), .A4(new_n626), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n630), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n619), .A2(G169), .A3(new_n636), .A4(new_n627), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n625), .A2(G179), .A3(new_n468), .A4(new_n626), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n619), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n631), .A2(new_n635), .A3(new_n637), .A4(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n558), .A2(new_n611), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n462), .A2(new_n521), .A3(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n321), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n398), .A2(KEYINPUT89), .A3(new_n399), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT89), .B1(new_n398), .B2(new_n399), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n380), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n269), .A2(new_n271), .A3(new_n291), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n384), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT17), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n459), .B(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n454), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n644), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n462), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n506), .A2(new_n516), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n535), .A2(new_n540), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n555), .A2(new_n556), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n628), .A2(new_n630), .B1(new_n619), .B2(new_n639), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n637), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n268), .B1(new_n480), .B2(new_n484), .ZN(new_n662));
  INV_X1    g0462(.A(new_n517), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n520), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT86), .B1(new_n605), .B2(new_n608), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT86), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n606), .A2(new_n607), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(G169), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n604), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n551), .A2(new_n598), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n656), .A2(new_n661), .A3(new_n664), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n669), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n664), .A2(new_n611), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n598), .A2(new_n669), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT87), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n664), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n662), .A2(new_n663), .A3(KEYINPUT87), .A4(new_n520), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT26), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n674), .B1(new_n679), .B2(KEYINPUT88), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n664), .A2(new_n676), .ZN(new_n681));
  INV_X1    g0481(.A(new_n675), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n673), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT88), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n672), .B1(new_n680), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n654), .B1(new_n655), .B2(new_n687), .ZN(G369));
  AOI21_X1  g0488(.A(new_n557), .B1(new_n535), .B2(new_n540), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n551), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n657), .B2(new_n695), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n699), .B2(new_n689), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n631), .A2(new_n637), .A3(new_n640), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n632), .A2(new_n696), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n641), .B2(new_n702), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n701), .A2(new_n696), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n700), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(new_n697), .A3(new_n709), .ZN(G399));
  NAND3_X1  g0510(.A1(new_n581), .A2(new_n613), .A3(new_n583), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT90), .Z(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n211), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n214), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n568), .A2(new_n574), .B1(G200), .B2(new_n596), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n601), .A2(new_n602), .A3(new_n595), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n720), .A2(new_n721), .B1(new_n604), .B2(new_n609), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n519), .A2(new_n722), .A3(new_n673), .A4(new_n520), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n669), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(KEYINPUT26), .B2(new_n683), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT92), .B1(new_n689), .B2(new_n701), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n659), .A2(new_n727), .A3(new_n637), .A4(new_n660), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n521), .A2(new_n729), .A3(new_n670), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n695), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n680), .A2(new_n686), .ZN(new_n733));
  INV_X1    g0533(.A(new_n672), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n695), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n732), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n642), .A2(new_n664), .A3(new_n656), .A4(new_n696), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n546), .A2(new_n547), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n638), .A2(new_n740), .A3(new_n596), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n507), .A2(new_n741), .A3(new_n508), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n507), .A2(new_n741), .A3(KEYINPUT30), .A4(new_n508), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n667), .A2(G179), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n486), .A2(new_n627), .A3(new_n746), .A4(new_n548), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n695), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n739), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n738), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n719), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR2_X1   g0557(.A1(new_n383), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n270), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G97), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n208), .A2(new_n270), .A3(KEYINPUT96), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT96), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G20), .B2(G179), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT100), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n769), .A2(KEYINPUT100), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n761), .B1(new_n773), .B2(new_n203), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT101), .Z(new_n775));
  NOR2_X1   g0575(.A1(new_n208), .A2(G179), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n768), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT99), .Z(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G107), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n766), .A2(new_n758), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n766), .A2(new_n781), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n779), .B1(new_n202), .B2(new_n780), .C1(new_n220), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n776), .A2(new_n781), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT98), .B(KEYINPUT32), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n788), .A2(G159), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n383), .A2(new_n767), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n776), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n222), .ZN(new_n793));
  INV_X1    g0593(.A(new_n791), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n765), .A2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n366), .B(new_n793), .C1(new_n795), .C2(G50), .ZN(new_n796));
  INV_X1    g0596(.A(new_n789), .ZN(new_n797));
  INV_X1    g0597(.A(G159), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n787), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n790), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n775), .A2(new_n783), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT33), .B(G317), .Z(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n773), .A2(new_n802), .B1(new_n803), .B2(new_n780), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT102), .ZN(new_n805));
  INV_X1    g0605(.A(new_n792), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n257), .B1(new_n806), .B2(G303), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  INV_X1    g0608(.A(new_n760), .ZN(new_n809));
  INV_X1    g0609(.A(new_n795), .ZN(new_n810));
  INV_X1    g0610(.A(G326), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n807), .B1(new_n808), .B2(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G329), .A2(new_n788), .B1(new_n778), .B2(G283), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n782), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n805), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n801), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(KEYINPUT103), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(KEYINPUT103), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n216), .B1(G20), .B2(new_n268), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n208), .A2(G13), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n207), .B1(new_n822), .B2(G45), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n715), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT94), .Z(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n714), .A2(new_n366), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(G355), .B1(new_n613), .B2(new_n714), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n714), .A2(new_n257), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(G45), .B2(new_n214), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT95), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n243), .A2(new_n249), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(G13), .A2(G33), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(G20), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n820), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n827), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n837), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n821), .B(new_n839), .C1(new_n704), .C2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n705), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n704), .A2(G330), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n842), .A2(new_n825), .A3(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT93), .Z(new_n845));
  NAND2_X1  g0645(.A1(new_n841), .A2(new_n845), .ZN(G396));
  NAND4_X1  g0646(.A1(new_n269), .A2(new_n271), .A3(new_n291), .A4(new_n696), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n293), .A2(new_n294), .B1(new_n291), .B2(new_n695), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n649), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n296), .A2(new_n696), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n735), .A2(new_n850), .B1(new_n687), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n825), .B1(new_n852), .B2(new_n754), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n754), .B2(new_n852), .ZN(new_n854));
  INV_X1    g0654(.A(new_n780), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n855), .A2(G143), .B1(G137), .B2(new_n795), .ZN(new_n856));
  INV_X1    g0656(.A(G150), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n798), .B2(new_n782), .C1(new_n773), .C2(new_n857), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT34), .Z(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n787), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n778), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n203), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n257), .B1(new_n792), .B2(new_n201), .C1(new_n809), .C2(new_n202), .ZN(new_n864));
  NOR4_X1   g0664(.A1(new_n859), .A2(new_n861), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n257), .B1(new_n806), .B2(G107), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n761), .B(new_n866), .C1(new_n780), .C2(new_n808), .ZN(new_n867));
  INV_X1    g0667(.A(new_n782), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n868), .A2(G116), .B1(G303), .B2(new_n795), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n778), .A2(G87), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n869), .B(new_n870), .C1(new_n814), .C2(new_n787), .ZN(new_n871));
  INV_X1    g0671(.A(new_n773), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n867), .B(new_n871), .C1(G283), .C2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n820), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n820), .A2(new_n835), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n827), .B1(new_n220), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n876), .C1(new_n850), .C2(new_n836), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n854), .A2(new_n877), .ZN(G384));
  INV_X1    g0678(.A(new_n693), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n454), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n425), .B1(KEYINPUT16), .B2(new_n424), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n693), .B1(new_n881), .B2(new_n405), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n441), .A2(new_n453), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n652), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n450), .A2(new_n451), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n450), .A2(new_n879), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n459), .ZN(new_n888));
  INV_X1    g0688(.A(new_n459), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n881), .A2(new_n405), .B1(new_n440), .B2(new_n693), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n884), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT39), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n897));
  INV_X1    g0697(.A(new_n886), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n885), .A2(new_n886), .A3(new_n459), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n461), .A2(new_n898), .B1(new_n888), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n896), .B(new_n897), .C1(new_n901), .C2(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n648), .A2(new_n696), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n880), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT106), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n847), .B1(new_n687), .B2(new_n851), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT105), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n342), .A2(new_n347), .A3(new_n909), .A4(new_n695), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT105), .B1(new_n381), .B2(new_n696), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n380), .A2(new_n384), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n348), .B(new_n695), .C1(new_n377), .C2(new_n379), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n908), .B(new_n914), .C1(new_n893), .C2(new_n894), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n906), .A2(new_n907), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n907), .B1(new_n906), .B2(new_n915), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n462), .B(new_n732), .C1(new_n735), .C2(new_n737), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n654), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n893), .A2(new_n894), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n849), .B1(new_n912), .B2(new_n913), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT108), .B1(new_n753), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n753), .A2(new_n924), .A3(KEYINPUT108), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n897), .B1(new_n901), .B2(KEYINPUT38), .ZN(new_n929));
  AND4_X1   g0729(.A1(KEYINPUT40), .A2(new_n929), .A3(new_n753), .A4(new_n924), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n462), .A3(new_n753), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n462), .A2(new_n753), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n928), .B2(new_n930), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(G330), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n921), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n936), .A2(KEYINPUT109), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(KEYINPUT109), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n921), .A2(new_n935), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n822), .A2(new_n207), .ZN(new_n940));
  NOR4_X1   g0740(.A1(new_n937), .A2(new_n938), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n493), .B(KEYINPUT104), .Z(new_n942));
  INV_X1    g0742(.A(KEYINPUT35), .ZN(new_n943));
  OAI211_X1 g0743(.A(G116), .B(new_n217), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT36), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n215), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n201), .A2(G68), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n207), .B(G13), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n941), .A2(new_n946), .A3(new_n949), .ZN(G367));
  OAI211_X1 g0750(.A(new_n656), .B(new_n664), .C1(new_n515), .C2(new_n696), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT110), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n519), .A2(new_n520), .A3(new_n695), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n709), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n664), .B1(new_n952), .B2(new_n659), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n956), .A2(KEYINPUT42), .B1(new_n957), .B2(new_n696), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(KEYINPUT42), .B2(new_n956), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n721), .A2(new_n696), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n682), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n669), .B2(new_n960), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n959), .A2(KEYINPUT43), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n707), .B1(new_n952), .B2(new_n953), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n959), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n963), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n964), .B1(new_n963), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n715), .B(KEYINPUT41), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n709), .A2(new_n697), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n952), .B2(new_n953), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n952), .A2(new_n973), .A3(new_n953), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT44), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n706), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n700), .B(new_n708), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(KEYINPUT111), .B2(new_n705), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n705), .B(KEYINPUT111), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n755), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n974), .B(KEYINPUT45), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n977), .B(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n989), .A3(new_n707), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n979), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n972), .B1(new_n991), .B2(new_n756), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n992), .A2(KEYINPUT112), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n823), .B1(new_n992), .B2(KEYINPUT112), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n971), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n830), .A2(new_n238), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n837), .B(new_n820), .C1(new_n714), .C2(new_n282), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n827), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n792), .A2(new_n613), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n366), .B1(new_n579), .B2(new_n777), .C1(new_n999), .C2(KEYINPUT46), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n788), .A2(G317), .B1(G311), .B2(new_n795), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n623), .B2(new_n780), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(KEYINPUT46), .C2(new_n999), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n808), .B2(new_n773), .ZN(new_n1004));
  INV_X1    g0804(.A(G283), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n782), .A2(new_n1005), .B1(new_n262), .B2(new_n809), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT113), .Z(new_n1007));
  OAI22_X1  g0807(.A1(new_n773), .A2(new_n798), .B1(new_n201), .B2(new_n782), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(KEYINPUT114), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n257), .B1(new_n777), .B2(new_n220), .C1(new_n202), .C2(new_n792), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G68), .B2(new_n760), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n788), .A2(G137), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n855), .A2(G150), .B1(G143), .B2(new_n795), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1008), .A2(KEYINPUT114), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1004), .A2(new_n1007), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT47), .Z(new_n1017));
  INV_X1    g0817(.A(new_n820), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n998), .B1(new_n840), .B2(new_n962), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n995), .A2(new_n1019), .ZN(G387));
  AOI22_X1  g0820(.A1(new_n712), .A2(new_n828), .B1(new_n262), .B2(new_n714), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n235), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n830), .B1(new_n1022), .B2(new_n249), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n713), .A2(KEYINPUT115), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n713), .A2(KEYINPUT115), .ZN(new_n1025));
  AND3_X1   g0825(.A1(new_n287), .A2(KEYINPUT50), .A3(new_n201), .ZN(new_n1026));
  AOI21_X1  g0826(.A(KEYINPUT50), .B1(new_n287), .B2(new_n201), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n249), .B1(new_n203), .B2(new_n220), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1021), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1030), .A2(new_n838), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n855), .A2(G50), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n760), .A2(new_n282), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n806), .A2(G77), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1032), .A2(new_n257), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n778), .A2(G97), .B1(G159), .B2(new_n795), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n203), .B2(new_n782), .C1(new_n857), .C2(new_n787), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1035), .B(new_n1037), .C1(new_n287), .C2(new_n872), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT116), .Z(new_n1039));
  INV_X1    g0839(.A(new_n777), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n257), .B1(new_n1040), .B2(G116), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n809), .A2(new_n1005), .B1(new_n792), .B2(new_n808), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n868), .A2(G303), .B1(G322), .B2(new_n795), .ZN(new_n1043));
  INV_X1    g0843(.A(G317), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n780), .C1(new_n773), .C2(new_n814), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT49), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1041), .B1(new_n811), .B2(new_n787), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1039), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n827), .B(new_n1031), .C1(new_n1052), .C2(new_n820), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n700), .A2(new_n837), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1053), .A2(new_n1054), .B1(new_n984), .B2(new_n824), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n756), .A2(new_n984), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n715), .B1(new_n755), .B2(new_n985), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(G393));
  AND2_X1   g0858(.A1(new_n979), .A2(new_n990), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n824), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n830), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n838), .B1(new_n579), .B2(new_n211), .C1(new_n1061), .C2(new_n246), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n810), .A2(new_n857), .B1(new_n780), .B2(new_n798), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT51), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n809), .A2(new_n220), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n366), .B(new_n1065), .C1(G68), .C2(new_n806), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n287), .A2(new_n868), .B1(new_n788), .B2(G143), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n870), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G50), .B2(new_n872), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n808), .A2(new_n782), .B1(new_n787), .B2(new_n803), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n257), .B1(new_n806), .B2(G283), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n779), .B(new_n1071), .C1(new_n613), .C2(new_n809), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(new_n872), .C2(G303), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n810), .A2(new_n1044), .B1(new_n780), .B2(new_n814), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1064), .A2(new_n1069), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n826), .B(new_n1062), .C1(new_n1076), .C2(new_n1018), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT117), .Z(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n954), .B2(new_n840), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1060), .A2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1059), .A2(new_n986), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n991), .A2(new_n715), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(KEYINPUT118), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n753), .A2(new_n850), .A3(G330), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n914), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n683), .A2(KEYINPUT26), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n724), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n730), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n848), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n292), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n696), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n753), .A2(new_n924), .A3(G330), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n847), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1088), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1086), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1095), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1097), .A2(new_n1098), .B1(new_n908), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n462), .A2(G330), .A3(new_n753), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n919), .A2(new_n654), .A3(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n731), .A2(new_n1093), .B1(new_n649), .B2(new_n696), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n904), .B(new_n929), .C1(new_n1105), .C2(new_n1087), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n905), .B1(new_n908), .B2(new_n914), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n903), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1095), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1106), .B(new_n1095), .C1(new_n1107), .C2(new_n903), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1104), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1112), .A2(new_n715), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT119), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n919), .A2(new_n654), .A3(new_n1102), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1099), .A2(KEYINPUT118), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1116), .A2(new_n1105), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1100), .A2(new_n908), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1115), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1114), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1123), .A2(KEYINPUT120), .A3(new_n1114), .A4(new_n1121), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1113), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1110), .A2(new_n824), .A3(new_n1111), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n875), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n826), .B1(new_n287), .B2(new_n1129), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n863), .A2(new_n257), .A3(new_n793), .A4(new_n1065), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n868), .A2(G97), .B1(G283), .B2(new_n795), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G116), .A2(new_n855), .B1(new_n788), .B2(G294), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n773), .A2(new_n262), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n257), .B1(new_n777), .B2(new_n201), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n788), .B2(G125), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT121), .Z(new_n1138));
  INV_X1    g0938(.A(G128), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n810), .A2(new_n1139), .B1(new_n782), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G132), .B2(new_n855), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n792), .A2(new_n857), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT53), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n809), .A2(new_n798), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1144), .B2(new_n1143), .ZN(new_n1146));
  INV_X1    g0946(.A(G137), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1142), .B(new_n1146), .C1(new_n1147), .C2(new_n773), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1134), .A2(new_n1135), .B1(new_n1138), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1130), .B1(new_n1149), .B2(new_n820), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n903), .B2(new_n836), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1128), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1127), .A2(new_n1153), .ZN(G378));
  OAI21_X1  g0954(.A(new_n321), .B1(new_n645), .B2(new_n646), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n388), .A2(new_n693), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n835), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n825), .B1(G50), .B2(new_n1129), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G50), .B1(new_n409), .B2(new_n248), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n282), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n810), .A2(new_n613), .B1(new_n782), .B2(new_n1163), .ZN(new_n1164));
  AOI211_X1 g0964(.A(G41), .B(new_n257), .C1(new_n806), .C2(G77), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n202), .B2(new_n777), .C1(new_n203), .C2(new_n809), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G283), .C2(new_n788), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n780), .A2(new_n262), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT122), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(new_n579), .C2(new_n773), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1162), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G128), .A2(new_n855), .B1(new_n868), .B2(G137), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n795), .A2(G125), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1140), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n760), .A2(G150), .B1(new_n806), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G132), .B2(new_n872), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n283), .B(new_n248), .C1(new_n777), .C2(new_n798), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n788), .B2(G124), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT59), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1182), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1172), .B1(new_n1171), .B2(new_n1170), .C1(new_n1180), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1161), .B1(new_n1185), .B2(new_n820), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1160), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n931), .A2(G330), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n916), .A2(new_n917), .A3(new_n1159), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1158), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1157), .B(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n906), .A2(new_n915), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT106), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n906), .A2(new_n907), .A3(new_n915), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1191), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1188), .B1(new_n1189), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1159), .B1(new_n916), .B2(new_n917), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(new_n1194), .A3(new_n1191), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1188), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1187), .B1(new_n1201), .B2(new_n823), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT123), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1112), .A2(new_n1203), .A3(new_n1115), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1200), .B(new_n1196), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n716), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1199), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(KEYINPUT57), .C1(new_n1205), .C2(new_n1204), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1202), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(G375));
  AOI21_X1  g1014(.A(new_n366), .B1(new_n1040), .B2(G58), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n798), .B2(new_n792), .C1(new_n201), .C2(new_n809), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n868), .A2(G150), .B1(G132), .B2(new_n795), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n1139), .B2(new_n787), .C1(new_n1147), .C2(new_n780), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(new_n872), .C2(new_n1175), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n257), .B1(new_n806), .B2(G97), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1033), .B(new_n1220), .C1(new_n782), .C2(new_n262), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n788), .A2(G303), .B1(G294), .B2(new_n795), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n220), .B2(new_n862), .C1(new_n1005), .C2(new_n780), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(G116), .C2(new_n872), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n820), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n826), .C1(G68), .C2(new_n1129), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n835), .B2(new_n1087), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1119), .B2(new_n824), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n972), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1122), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT124), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(KEYINPUT124), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1228), .B1(new_n1230), .B2(new_n1235), .ZN(G381));
  NAND3_X1  g1036(.A1(new_n995), .A2(new_n1019), .A3(new_n1083), .ZN(new_n1237));
  OR4_X1    g1037(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G378), .A2(G375), .A3(new_n1237), .A4(new_n1238), .ZN(G407));
  NAND3_X1  g1039(.A1(new_n1123), .A2(new_n1114), .A3(new_n1121), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT120), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1125), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1152), .B1(new_n1243), .B2(new_n1113), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n694), .A2(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1213), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(G407), .A2(G213), .A3(new_n1247), .ZN(G409));
  AOI21_X1  g1048(.A(new_n716), .B1(new_n1231), .B2(KEYINPUT60), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT60), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1104), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1235), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1228), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n854), .A3(new_n877), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(G384), .A3(new_n1228), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1244), .B(new_n1202), .C1(new_n1208), .C2(new_n1212), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1211), .B(new_n1229), .C1(new_n1205), .C2(new_n1204), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1211), .A2(new_n824), .B1(new_n1160), .B2(new_n1186), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G378), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1245), .B(new_n1256), .C1(new_n1257), .C2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1208), .A2(new_n1212), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(G378), .A3(new_n1259), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1260), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1245), .A4(new_n1256), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1246), .A2(G2897), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT126), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1245), .B1(new_n1272), .B2(G2897), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1272), .B2(G2897), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1254), .A2(new_n1255), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1254), .A2(KEYINPUT127), .A3(new_n1255), .A4(new_n1274), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1271), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1260), .B1(new_n1213), .B2(G378), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1246), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1262), .A2(new_n1263), .A3(new_n1269), .A4(new_n1281), .ZN(new_n1282));
  XOR2_X1   g1082(.A(G393), .B(G396), .Z(new_n1283));
  AND3_X1   g1083(.A1(new_n995), .A2(new_n1019), .A3(new_n1083), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1083), .B1(new_n995), .B2(new_n1019), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1283), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G387), .A2(G390), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1283), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1237), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1282), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1286), .A2(new_n1289), .A3(new_n1263), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n1261), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT125), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1280), .B2(new_n1246), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1267), .A2(KEYINPUT125), .A3(new_n1245), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1279), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1261), .A2(new_n1293), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1294), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1291), .A2(new_n1300), .ZN(G405));
  NAND2_X1  g1101(.A1(G375), .A2(new_n1244), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1265), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1290), .A2(new_n1265), .A3(new_n1302), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1256), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1304), .A2(new_n1256), .A3(new_n1305), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(G402));
endmodule


