//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G355));
  NOR2_X1   g0005(.A1(G58), .A2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT66), .B(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G58), .A2(G232), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n214), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n213), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT68), .ZN(new_n246));
  AND2_X1   g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n246), .B1(new_n247), .B2(new_n210), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND4_X1  g0049(.A1(new_n249), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n248), .A2(new_n250), .A3(G232), .A4(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(new_n248), .A3(new_n250), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT80), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT80), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(new_n261), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(G223), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(G226), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G87), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n264), .A2(new_n267), .B1(new_n258), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n247), .A2(new_n210), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n257), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G179), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G169), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n257), .B2(new_n271), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT16), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n206), .B1(new_n218), .B2(G58), .ZN(new_n279));
  INV_X1    g0079(.A(G159), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI22_X1  g0082(.A1(new_n279), .A2(new_n211), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT7), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n261), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n263), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n219), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n278), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT70), .B1(new_n214), .B2(new_n258), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT70), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n293), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n210), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT81), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n264), .A2(new_n284), .A3(new_n211), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G68), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n284), .B1(new_n264), .B2(new_n211), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI221_X1 g0101(.A(KEYINPUT16), .B1(new_n280), .B2(new_n282), .C1(new_n279), .C2(new_n211), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT7), .B1(new_n304), .B2(G20), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(G68), .A3(new_n298), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT66), .A2(G68), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT66), .A2(G68), .ZN(new_n308));
  OAI21_X1  g0108(.A(G58), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n211), .B1(new_n309), .B2(new_n207), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n282), .A2(new_n280), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n310), .A2(new_n278), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n306), .A2(KEYINPUT81), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n296), .B1(new_n303), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n251), .A2(G20), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n292), .A2(new_n210), .A3(new_n294), .A4(new_n319), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n318), .A2(new_n320), .B1(new_n319), .B2(new_n316), .ZN(new_n321));
  OAI211_X1 g0121(.A(KEYINPUT18), .B(new_n277), .C1(new_n314), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT82), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n292), .A2(new_n210), .A3(new_n294), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n286), .A2(new_n289), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n218), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n310), .A2(new_n311), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n329), .B2(new_n278), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n306), .A2(KEYINPUT81), .A3(new_n312), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT81), .B1(new_n306), .B2(new_n312), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n321), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n335), .A2(KEYINPUT82), .A3(KEYINPUT18), .A4(new_n277), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT18), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n303), .A2(new_n313), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n321), .B1(new_n338), .B2(new_n330), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n274), .A2(new_n276), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n324), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n272), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n257), .B2(new_n271), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT17), .B1(new_n339), .B2(new_n347), .ZN(new_n348));
  AND4_X1   g0148(.A1(KEYINPUT17), .A2(new_n333), .A3(new_n334), .A4(new_n347), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n270), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n288), .A2(G1698), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G222), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n285), .A2(G223), .A3(G1698), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n288), .A2(G77), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT69), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n352), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n358), .B2(new_n357), .ZN(new_n360));
  INV_X1    g0160(.A(new_n256), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n248), .A2(new_n250), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n363), .A2(new_n252), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n361), .B1(new_n364), .B2(G226), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g0166(.A(KEYINPUT72), .B(G200), .Z(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n360), .A2(G190), .A3(new_n365), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n281), .A2(G150), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n211), .A2(G33), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n371), .B1(new_n201), .B2(new_n211), .C1(new_n315), .C2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G50), .ZN(new_n374));
  INV_X1    g0174(.A(new_n319), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n373), .A2(new_n295), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n320), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(G50), .A3(new_n317), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(KEYINPUT9), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n378), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT9), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n380), .A2(new_n381), .B1(KEYINPUT73), .B2(KEYINPUT10), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n369), .A2(new_n370), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n383), .B(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n361), .B1(new_n364), .B2(G244), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n353), .A2(G232), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT71), .ZN(new_n388));
  INV_X1    g0188(.A(G107), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(KEYINPUT71), .A2(G107), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n387), .B1(new_n285), .B2(new_n393), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n288), .A2(new_n220), .A3(new_n266), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n270), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n386), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(G169), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n316), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT15), .B(G87), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n372), .B2(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n295), .B1(new_n202), .B2(new_n375), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n377), .A2(G77), .A3(new_n317), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(G179), .B2(new_n397), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n398), .B2(G190), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n398), .B2(new_n367), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n366), .A2(new_n275), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n380), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n366), .A2(G179), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n351), .A2(new_n385), .A3(new_n411), .A4(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n218), .A2(new_n211), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n282), .A2(new_n374), .B1(new_n372), .B2(new_n202), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n295), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT11), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  INV_X1    g0222(.A(G68), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT12), .B1(new_n375), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G13), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G1), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n426), .A2(KEYINPUT12), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n417), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n377), .A2(G68), .A3(new_n317), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n421), .A2(new_n422), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  AND4_X1   g0230(.A1(G238), .A2(new_n248), .A3(new_n252), .A4(new_n250), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT75), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n256), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n255), .A2(new_n248), .A3(KEYINPUT75), .A4(new_n250), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n263), .A2(new_n287), .A3(G232), .A4(G1698), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT74), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT74), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n285), .A2(new_n438), .A3(G232), .A4(G1698), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G97), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n285), .A2(G226), .A3(new_n266), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n437), .A2(new_n439), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n270), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT13), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n435), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n435), .B2(new_n443), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n430), .B1(new_n448), .B2(G190), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n435), .A2(new_n443), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT13), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n445), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(G200), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(G169), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT14), .ZN(new_n459));
  XOR2_X1   g0259(.A(KEYINPUT77), .B(KEYINPUT14), .Z(new_n460));
  NAND4_X1  g0260(.A1(new_n453), .A2(G169), .A3(new_n454), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n451), .A2(G179), .A3(new_n445), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT78), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n451), .A2(KEYINPUT78), .A3(G179), .A4(new_n445), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n459), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n457), .B1(new_n467), .B2(new_n430), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT79), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n468), .A2(KEYINPUT79), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n416), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n258), .A2(G1), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n377), .A2(G116), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT87), .B(G116), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n375), .ZN(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(new_n258), .B2(G97), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n476), .A2(G20), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n480), .A2(KEYINPUT20), .A3(new_n295), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT20), .B1(new_n480), .B2(new_n295), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n475), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G257), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n266), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G264), .B2(new_n266), .ZN(new_n487));
  INV_X1    g0287(.A(G303), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n264), .A2(new_n487), .B1(new_n488), .B2(new_n285), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT89), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI221_X1 g0291(.A(KEYINPUT89), .B1(new_n488), .B2(new_n285), .C1(new_n264), .C2(new_n487), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n270), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n251), .A2(G45), .A3(G274), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n248), .A2(new_n496), .A3(new_n250), .A4(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT85), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n497), .B1(new_n494), .B2(new_n495), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(KEYINPUT85), .A3(new_n248), .A4(new_n250), .ZN(new_n503));
  INV_X1    g0303(.A(G45), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(G1), .ZN(new_n505));
  INV_X1    g0305(.A(new_n495), .ZN(new_n506));
  NOR2_X1   g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n508), .A2(new_n248), .A3(new_n250), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n501), .A2(new_n503), .B1(new_n509), .B2(G270), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n493), .A2(new_n510), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n484), .A2(new_n511), .A3(new_n273), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n511), .A2(KEYINPUT21), .A3(G169), .A4(new_n483), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT90), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n275), .B1(new_n493), .B2(new_n510), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT90), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT21), .A4(new_n483), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n512), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n345), .B1(new_n493), .B2(new_n510), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT92), .ZN(new_n520));
  OR3_X1    g0320(.A1(new_n519), .A2(new_n520), .A3(new_n483), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n519), .B2(new_n483), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n493), .A2(new_n510), .A3(G190), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n515), .A2(new_n483), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT91), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT91), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n515), .A2(new_n528), .A3(new_n483), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n518), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  INV_X1    g0332(.A(G97), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n390), .A2(new_n268), .A3(new_n533), .A4(new_n391), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n440), .A2(new_n211), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n372), .A2(KEYINPUT19), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n211), .A2(G68), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n536), .A2(new_n537), .B1(new_n264), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n295), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n401), .A2(new_n375), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n325), .A2(KEYINPUT83), .A3(new_n319), .A4(new_n474), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT83), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n320), .B2(new_n473), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(G87), .A3(new_n544), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n220), .A2(G1698), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n304), .A2(KEYINPUT86), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT86), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n266), .A2(G238), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n264), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g0352(.A(KEYINPUT87), .B(G116), .Z(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G33), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n259), .A2(new_n262), .A3(G244), .A4(new_n263), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(new_n266), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n270), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G250), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n497), .B1(new_n505), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n363), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(G190), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n304), .A2(G244), .A3(G1698), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n562), .A2(new_n548), .A3(new_n554), .A4(new_n551), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(new_n270), .B1(new_n363), .B2(new_n559), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n546), .B(new_n561), .C1(new_n367), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n557), .A2(new_n273), .A3(new_n560), .ZN(new_n566));
  INV_X1    g0366(.A(new_n401), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n542), .A2(new_n567), .A3(new_n544), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n540), .A2(new_n541), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n566), .B(new_n569), .C1(G169), .C2(new_n564), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT88), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT88), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n565), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n501), .A2(new_n503), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AND4_X1   g0377(.A1(G264), .A2(new_n508), .A3(new_n248), .A4(new_n250), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G294), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n485), .A2(G1698), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(G250), .B2(G1698), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n264), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n270), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n577), .A2(new_n585), .A3(G190), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT93), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n583), .A2(new_n270), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n578), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n579), .A2(new_n584), .A3(KEYINPUT93), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n576), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n586), .B1(new_n591), .B2(new_n345), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT22), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n211), .A2(G87), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n288), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT23), .B1(new_n392), .B2(new_n211), .ZN(new_n597));
  OR3_X1    g0397(.A1(new_n211), .A2(KEYINPUT23), .A3(G107), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n594), .A2(new_n268), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n259), .A2(new_n601), .A3(new_n262), .A4(new_n263), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n554), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n211), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n593), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(G20), .B1(new_n554), .B2(new_n602), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n606), .A2(new_n599), .A3(KEYINPUT24), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n295), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n542), .A2(G107), .A3(new_n544), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n319), .A2(G107), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT25), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n592), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n263), .A2(new_n287), .A3(G250), .A4(G1698), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n479), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  AND2_X1   g0417(.A1(KEYINPUT4), .A2(G244), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n285), .A2(new_n617), .A3(new_n266), .A4(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n263), .A2(new_n287), .A3(new_n618), .A4(new_n266), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT84), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n616), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT4), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n555), .B2(G1698), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n352), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n509), .A2(G257), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n576), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(G190), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT6), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n630), .A2(new_n533), .A3(G107), .ZN(new_n631));
  XNOR2_X1  g0431(.A(G97), .B(G107), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n633), .A2(new_n211), .B1(new_n202), .B2(new_n282), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n393), .B1(new_n286), .B2(new_n289), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n295), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n542), .A2(G97), .A3(new_n544), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n375), .A2(new_n533), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n576), .A2(new_n627), .ZN(new_n641));
  OAI21_X1  g0441(.A(G200), .B1(new_n625), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n629), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n626), .A2(new_n273), .A3(new_n628), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n275), .B1(new_n625), .B2(new_n641), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n639), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(G169), .B1(new_n577), .B2(new_n585), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n589), .A2(G179), .A3(new_n576), .A4(new_n590), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n648), .A2(new_n649), .B1(new_n608), .B2(new_n612), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n614), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n472), .A2(new_n531), .A3(new_n575), .A4(new_n651), .ZN(G372));
  XOR2_X1   g0452(.A(new_n383), .B(new_n384), .Z(new_n653));
  INV_X1    g0453(.A(new_n350), .ZN(new_n654));
  AOI211_X1 g0454(.A(new_n406), .B(new_n399), .C1(new_n273), .C2(new_n398), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n456), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n467), .A2(new_n430), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n340), .B1(new_n333), .B2(new_n334), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(KEYINPUT18), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n339), .A2(new_n337), .A3(new_n340), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n653), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n415), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n644), .A2(new_n645), .A3(new_n639), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n570), .A4(new_n565), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(new_n570), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n646), .B1(new_n572), .B2(new_n574), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n667), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n649), .A2(new_n648), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n613), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT94), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n518), .A2(new_n674), .A3(new_n530), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n518), .B2(new_n530), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n614), .A2(new_n647), .A3(new_n571), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n671), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n665), .B1(new_n471), .B2(new_n679), .ZN(G369));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n518), .A2(new_n530), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT94), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n518), .A2(new_n530), .A3(new_n674), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n426), .A2(new_n211), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(KEYINPUT95), .B(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n484), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n683), .A2(new_n684), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n692), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n531), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n681), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n613), .A2(new_n690), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n673), .B(new_n697), .C1(new_n613), .C2(new_n592), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT96), .B1(new_n650), .B2(new_n690), .ZN(new_n699));
  AND4_X1   g0499(.A1(KEYINPUT96), .A2(new_n672), .A3(new_n613), .A4(new_n690), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n690), .B1(new_n518), .B2(new_n530), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n701), .A2(new_n703), .B1(new_n650), .B2(new_n691), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n215), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n534), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n208), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n518), .A2(new_n530), .A3(new_n673), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n678), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n570), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n565), .A2(new_n570), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n666), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n716), .B1(new_n718), .B2(KEYINPUT26), .ZN(new_n719));
  INV_X1    g0519(.A(new_n574), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n573), .B1(new_n565), .B2(new_n570), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n667), .B(new_n666), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n715), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n713), .B1(new_n723), .B2(new_n691), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n677), .A2(new_n678), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n668), .A2(new_n570), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n575), .A2(new_n666), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(KEYINPUT26), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n690), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n724), .B1(new_n729), .B2(new_n713), .ZN(new_n730));
  AND4_X1   g0530(.A1(new_n531), .A2(new_n651), .A3(new_n575), .A4(new_n691), .ZN(new_n731));
  INV_X1    g0531(.A(new_n564), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n626), .A2(new_n628), .ZN(new_n733));
  AOI21_X1  g0533(.A(G179), .B1(new_n493), .B2(new_n510), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n732), .A2(new_n733), .A3(new_n591), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n511), .A2(new_n273), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n579), .A2(new_n584), .A3(KEYINPUT93), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT93), .B1(new_n579), .B2(new_n584), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n625), .A2(new_n641), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n736), .A2(new_n739), .A3(new_n564), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(KEYINPUT98), .A2(KEYINPUT30), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n735), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n742), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n589), .A2(new_n557), .A3(new_n560), .A4(new_n590), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n733), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n744), .B1(new_n746), .B2(new_n736), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n690), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT97), .B(KEYINPUT31), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n690), .B(new_n752), .C1(new_n743), .C2(new_n747), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(G330), .B1(new_n731), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n730), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n712), .B1(new_n757), .B2(G1), .ZN(G364));
  NAND2_X1  g0558(.A1(new_n693), .A2(new_n695), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT99), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n425), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n251), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n707), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n696), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n765), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n211), .A2(G179), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n368), .A2(G190), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT102), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n771), .A2(G303), .B1(new_n774), .B2(G329), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n211), .A2(new_n273), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(G190), .A3(new_n345), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n288), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n776), .A2(new_n772), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n779), .B1(G311), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n368), .A2(new_n343), .A3(new_n769), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n775), .B(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n776), .A2(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(G317), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT33), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n788), .A2(KEYINPUT33), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n786), .A2(new_n343), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G326), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n343), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n211), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n791), .B(new_n793), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n784), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G107), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n771), .A2(G87), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n285), .B1(new_n780), .B2(new_n202), .ZN(new_n801));
  INV_X1    g0601(.A(new_n777), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G58), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n773), .A2(new_n280), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT32), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G68), .A2(new_n787), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n799), .A2(new_n800), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n796), .A2(new_n533), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n792), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n805), .B2(new_n804), .C1(new_n374), .C2(new_n810), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n785), .A2(new_n797), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n210), .B1(G20), .B2(new_n275), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n768), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n304), .A2(new_n706), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n504), .B2(new_n209), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n244), .B2(new_n504), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n706), .A2(new_n288), .ZN(new_n819));
  INV_X1    g0619(.A(G116), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G355), .A2(new_n819), .B1(new_n820), .B2(new_n706), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT100), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT101), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n818), .A2(new_n822), .A3(KEYINPUT101), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G13), .A2(G33), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(G20), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n813), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n827), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n814), .B1(new_n823), .B2(new_n829), .C1(new_n759), .C2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n767), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  NAND2_X1  g0633(.A1(new_n405), .A2(new_n690), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n410), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(new_n408), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n408), .A2(new_n690), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n411), .A2(new_n690), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n729), .A2(new_n838), .B1(new_n679), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n765), .B1(new_n841), .B2(new_n755), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n755), .B2(new_n841), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n813), .A2(new_n825), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n765), .B1(G77), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT103), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n784), .A2(new_n423), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G50), .B2(new_n771), .ZN(new_n849));
  INV_X1    g0649(.A(new_n796), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n264), .B1(new_n850), .B2(G58), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  INV_X1    g0652(.A(new_n774), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n849), .B(new_n851), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT104), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n802), .A2(G143), .B1(new_n781), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(new_n787), .ZN(new_n857));
  INV_X1    g0657(.A(G150), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n856), .B1(new_n857), .B2(new_n858), .C1(new_n859), .C2(new_n810), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT34), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n854), .A2(KEYINPUT104), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n809), .B1(new_n857), .B2(new_n783), .C1(new_n488), .C2(new_n810), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n288), .B1(new_n780), .B2(new_n476), .C1(new_n794), .C2(new_n777), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(G87), .B2(new_n798), .ZN(new_n866));
  INV_X1    g0666(.A(G311), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n866), .B1(new_n389), .B2(new_n770), .C1(new_n867), .C2(new_n853), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n862), .A2(new_n863), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n847), .B1(new_n869), .B2(new_n813), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n838), .B2(new_n826), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n843), .A2(new_n871), .ZN(G384));
  NOR2_X1   g0672(.A1(new_n762), .A2(new_n251), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n748), .A2(new_n751), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT31), .B(new_n690), .C1(new_n743), .C2(new_n747), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n838), .B1(new_n731), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n430), .A2(new_n690), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n657), .A2(new_n456), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT105), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n468), .A2(KEYINPUT105), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n467), .A2(new_n457), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(new_n878), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n877), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n328), .B1(new_n299), .B2(new_n300), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n325), .B1(new_n888), .B2(new_n278), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n331), .B2(new_n332), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n334), .ZN(new_n891));
  INV_X1    g0691(.A(new_n688), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n351), .A2(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n333), .A2(new_n334), .B1(new_n340), .B2(new_n688), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n333), .A2(new_n334), .A3(new_n347), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT37), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT106), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n321), .B1(new_n338), .B2(new_n889), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n898), .B(new_n900), .C1(new_n340), .C2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT37), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n891), .B2(new_n892), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n891), .A2(new_n277), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n900), .B1(new_n906), .B2(new_n898), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n899), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n895), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n893), .B1(new_n342), .B2(new_n350), .ZN(new_n912));
  INV_X1    g0712(.A(new_n898), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n903), .B1(new_n913), .B2(new_n896), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n902), .A2(new_n904), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n907), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n911), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT40), .B1(new_n887), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT17), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n898), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n339), .A2(KEYINPUT17), .A3(new_n347), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(new_n660), .C2(new_n661), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n339), .A2(new_n688), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n897), .A2(new_n898), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT107), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT37), .B1(new_n896), .B2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n927), .A2(new_n929), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n911), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n920), .B1(new_n933), .B2(new_n910), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n919), .B1(new_n887), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n531), .A2(new_n651), .A3(new_n575), .A4(new_n691), .ZN(new_n936));
  INV_X1    g0736(.A(new_n876), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n471), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n681), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n935), .B2(new_n938), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n924), .A2(new_n925), .B1(new_n927), .B2(new_n929), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n942), .B2(new_n930), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n912), .A2(new_n916), .A3(new_n911), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n657), .A2(new_n690), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n910), .A2(new_n917), .A3(KEYINPUT39), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n655), .A2(new_n691), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n679), .B2(new_n840), .ZN(new_n950));
  AND4_X1   g0750(.A1(KEYINPUT105), .A2(new_n657), .A3(new_n456), .A4(new_n878), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT105), .B1(new_n468), .B2(new_n878), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n886), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n950), .A2(new_n918), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n662), .A2(new_n688), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n948), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n665), .B1(new_n730), .B2(new_n471), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n873), .B1(new_n940), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n958), .B2(new_n940), .ZN(new_n960));
  INV_X1    g0760(.A(new_n633), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT35), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(KEYINPUT35), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n962), .A2(G116), .A3(new_n212), .A4(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT36), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n309), .A2(G50), .A3(G77), .A4(new_n207), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(G50), .B2(new_n423), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(G1), .A3(new_n425), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n960), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT108), .Z(G367));
  NAND2_X1  g0770(.A1(new_n701), .A2(new_n703), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n650), .A2(new_n691), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n643), .B(new_n646), .C1(new_n640), .C2(new_n691), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n666), .A2(new_n690), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT44), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n704), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n704), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT45), .B1(new_n704), .B2(new_n976), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n978), .A2(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n702), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n973), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n979), .B1(new_n704), .B2(new_n976), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n988), .B(new_n702), .C1(new_n981), .C2(new_n982), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n701), .B(new_n703), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(new_n696), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(new_n730), .A3(new_n755), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT109), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n992), .A2(new_n730), .A3(new_n755), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT109), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n995), .A2(new_n996), .A3(new_n989), .A4(new_n985), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n756), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n707), .B(KEYINPUT41), .Z(new_n999));
  OAI21_X1  g0799(.A(new_n763), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n701), .A2(new_n703), .A3(new_n976), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT42), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n646), .B1(new_n974), .B2(new_n673), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1001), .A2(KEYINPUT42), .B1(new_n691), .B2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n546), .A2(new_n691), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n717), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n570), .B2(new_n1005), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1002), .A2(new_n1004), .B1(KEYINPUT43), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n984), .A2(new_n976), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1000), .A2(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n794), .A2(new_n857), .B1(new_n810), .B2(new_n867), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n304), .B(new_n1014), .C1(new_n392), .C2(new_n850), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n773), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n802), .A2(G303), .B1(new_n1016), .B2(G317), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n783), .B2(new_n780), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G97), .B2(new_n798), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT46), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n771), .B2(G116), .ZN(new_n1021));
  NOR3_X1   g0821(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n476), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1015), .B(new_n1019), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT110), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n796), .A2(new_n423), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G150), .B2(new_n802), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT111), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n285), .B1(new_n773), .B2(new_n859), .C1(new_n374), .C2(new_n780), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n857), .A2(new_n280), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G143), .C2(new_n792), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n771), .A2(G58), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n798), .A2(G77), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1024), .B1(new_n1027), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT47), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n813), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n236), .A2(new_n815), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n813), .B(new_n827), .C1(new_n706), .C2(new_n567), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n768), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1036), .B(new_n1039), .C1(new_n830), .C2(new_n1007), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1013), .A2(new_n1040), .ZN(G387));
  AOI21_X1  g0841(.A(new_n304), .B1(G326), .B2(new_n1016), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n802), .A2(G317), .B1(new_n781), .B2(G303), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n857), .B2(new_n867), .C1(new_n778), .C2(new_n810), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n771), .A2(G294), .B1(G283), .B2(new_n850), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT113), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT49), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1042), .B1(new_n476), .B2(new_n784), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G68), .A2(new_n781), .B1(new_n1016), .B2(G150), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n374), .B2(new_n777), .C1(new_n533), .C2(new_n784), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n304), .B1(new_n857), .B2(new_n315), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n850), .A2(new_n567), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n810), .B2(new_n280), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n770), .A2(new_n202), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n813), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n819), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1062), .A2(new_n709), .B1(G107), .B2(new_n215), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n233), .A2(new_n504), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n709), .ZN(new_n1065));
  AOI211_X1 g0865(.A(G45), .B(new_n1065), .C1(G68), .C2(G77), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n315), .A2(G50), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT50), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n816), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1063), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT112), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n828), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1061), .B(new_n765), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n701), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1075), .B1(new_n1076), .B2(new_n827), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n764), .B2(new_n992), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n995), .A2(new_n708), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n757), .B2(new_n992), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(G393));
  NOR2_X1   g0881(.A1(new_n241), .A2(new_n816), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n828), .B1(new_n533), .B2(new_n215), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n765), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n288), .B1(new_n780), .B2(new_n794), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n857), .A2(new_n488), .B1(new_n476), .B2(new_n796), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G322), .C2(new_n1016), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n810), .A2(new_n788), .B1(new_n867), .B2(new_n777), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n771), .A2(G283), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1087), .A2(new_n799), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT116), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n264), .B1(new_n1016), .B2(G143), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n784), .B2(new_n268), .C1(new_n219), .C2(new_n770), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT115), .Z(new_n1095));
  OAI22_X1  g0895(.A1(new_n810), .A2(new_n858), .B1(new_n280), .B2(new_n777), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n787), .A2(G50), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n850), .A2(G77), .B1(new_n781), .B2(new_n316), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1092), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1084), .B1(new_n1101), .B2(new_n813), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n977), .A2(new_n827), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT114), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n985), .A2(new_n1105), .A3(new_n989), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n983), .A2(KEYINPUT114), .A3(new_n984), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(KEYINPUT117), .B(new_n1104), .C1(new_n1108), .C2(new_n763), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT117), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n763), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1104), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1106), .A2(new_n993), .A3(new_n1107), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT118), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT118), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1106), .A2(new_n1117), .A3(new_n993), .A4(new_n1107), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n708), .B1(new_n994), .B2(new_n997), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1114), .A2(new_n1121), .ZN(G390));
  AOI21_X1  g0922(.A(new_n885), .B1(new_n881), .B2(new_n882), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n838), .B(G330), .C1(new_n731), .C2(new_n876), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n946), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n943), .B2(new_n944), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n953), .A2(KEYINPUT119), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT119), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n883), .A2(new_n1129), .A3(new_n886), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n723), .A2(new_n691), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n949), .B1(new_n1132), .B2(new_n836), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1127), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n950), .A2(new_n953), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1135), .A2(new_n1126), .B1(new_n945), .B2(new_n947), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1125), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n725), .A2(new_n728), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n837), .B1(new_n1138), .B2(new_n839), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1126), .B1(new_n1139), .B2(new_n1123), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n945), .A2(new_n947), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n838), .B(G330), .C1(new_n731), .C2(new_n754), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n953), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1133), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1142), .B(new_n1145), .C1(new_n1147), .C2(new_n1127), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1137), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n681), .B1(new_n937), .B2(new_n936), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1150), .A2(new_n469), .A3(new_n470), .A4(new_n416), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n665), .C1(new_n730), .C2(new_n471), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1128), .A2(new_n1130), .A3(new_n1124), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1133), .B1(new_n1144), .B2(new_n953), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1144), .A2(new_n953), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n950), .B1(new_n1156), .B2(new_n1125), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1152), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1149), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1137), .A2(new_n1148), .A3(new_n1158), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n707), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1137), .A2(new_n1148), .A3(new_n764), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n288), .B1(new_n781), .B2(new_n1165), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n852), .B2(new_n777), .C1(new_n784), .C2(new_n374), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G125), .B2(new_n774), .ZN(new_n1168));
  OR3_X1    g0968(.A1(new_n770), .A2(KEYINPUT53), .A3(new_n858), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT53), .B1(new_n770), .B2(new_n858), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1171), .A2(new_n810), .B1(new_n857), .B2(new_n859), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G159), .B2(new_n850), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n810), .A2(new_n783), .B1(new_n780), .B2(new_n533), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n392), .B2(new_n787), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT120), .Z(new_n1177));
  OAI22_X1  g0977(.A1(new_n796), .A2(new_n202), .B1(new_n777), .B2(new_n820), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1178), .B(new_n848), .C1(G294), .C2(new_n774), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n800), .A2(new_n288), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT121), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1174), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT122), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n813), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n765), .B1(new_n316), .B2(new_n845), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT123), .Z(new_n1189));
  INV_X1    g0989(.A(new_n1141), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n826), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1163), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1162), .A2(new_n1193), .ZN(G378));
  INV_X1    g0994(.A(new_n1152), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1161), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n681), .B1(new_n887), .B2(new_n934), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n835), .A2(new_n408), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n949), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n937), .B2(new_n936), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n953), .A2(new_n918), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n920), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n380), .A2(new_n892), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n653), .A2(new_n664), .A3(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n380), .B(new_n892), .C1(new_n385), .C2(new_n415), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1206), .B(new_n1208), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1197), .A2(new_n1202), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n956), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n956), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1209), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n953), .A2(new_n1200), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT40), .B1(new_n943), .B2(new_n944), .ZN(new_n1216));
  OAI21_X1  g1016(.A(G330), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n919), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1197), .A2(new_n1202), .A3(new_n1209), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1213), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n707), .B1(new_n1196), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1161), .A2(new_n1195), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n956), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1218), .A2(new_n1213), .A3(new_n1219), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1222), .A2(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n787), .A2(G97), .B1(new_n781), .B2(new_n567), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT124), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n777), .A2(new_n389), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1231), .B(new_n1025), .C1(G116), .C2(new_n792), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1059), .B1(G283), .B2(new_n774), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n304), .A2(G41), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n798), .B2(G58), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1230), .A2(new_n1232), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT58), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n777), .A2(new_n1171), .B1(new_n780), .B2(new_n859), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G132), .B2(new_n787), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G150), .A2(new_n850), .B1(new_n792), .B2(G125), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n770), .C2(new_n1164), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n798), .A2(G159), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G33), .B(G41), .C1(new_n1016), .C2(G124), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1234), .B(new_n374), .C1(G33), .C2(G41), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1238), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n813), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n765), .C1(G50), .C2(new_n845), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1214), .B2(new_n825), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1226), .B2(new_n764), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1228), .A2(new_n1254), .ZN(G375));
  NAND2_X1  g1055(.A1(new_n1123), .A2(new_n1143), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1257), .A2(new_n950), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1152), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n999), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1159), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1131), .A2(new_n826), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n285), .B1(new_n781), .B2(new_n392), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1032), .B(new_n1263), .C1(new_n783), .C2(new_n777), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n853), .A2(new_n488), .B1(new_n533), .B2(new_n770), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1057), .B1(new_n857), .B2(new_n476), .C1(new_n794), .C2(new_n810), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n798), .A2(G58), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n781), .A2(G150), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n802), .A2(G137), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1268), .A2(new_n304), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G50), .A2(new_n850), .B1(new_n792), .B2(G132), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n857), .B2(new_n1164), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n853), .A2(new_n1171), .B1(new_n280), .B2(new_n770), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1271), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n813), .B1(new_n1267), .B2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1276), .B(new_n765), .C1(G68), .C2(new_n845), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1258), .A2(new_n763), .B1(new_n1262), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1261), .A2(new_n1279), .ZN(G381));
  INV_X1    g1080(.A(G375), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1040), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1000), .B2(new_n1012), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1078), .A2(new_n1284), .A3(new_n1080), .A4(new_n832), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(G378), .A2(G390), .A3(G381), .A4(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1281), .A2(new_n1283), .A3(new_n1286), .ZN(G407));
  AOI21_X1  g1087(.A(new_n708), .B1(new_n1149), .B2(new_n1159), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1192), .B1(new_n1288), .B2(new_n1161), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n689), .A2(G213), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1281), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(new_n1292), .A3(G213), .ZN(G409));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(G393), .B(new_n832), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(G390), .A2(new_n1013), .A3(new_n1040), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1283), .A2(G390), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G390), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G387), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1283), .A2(G390), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1295), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G378), .B(new_n1254), .C1(new_n1222), .C2(new_n1227), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1223), .A2(new_n1260), .A3(new_n1226), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1254), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1289), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1291), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT60), .B1(new_n1258), .B2(new_n1152), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1311), .A2(new_n1259), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1155), .A2(new_n1157), .A3(new_n1152), .A4(KEYINPUT60), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n707), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G384), .B(new_n1279), .C1(new_n1312), .C2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1259), .B2(new_n1311), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1284), .B1(new_n1316), .B2(new_n1278), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1315), .A2(new_n1317), .ZN(new_n1318));
  XOR2_X1   g1118(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1319));
  AND3_X1   g1119(.A1(new_n1310), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1291), .A2(G2897), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1315), .A2(new_n1317), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1321), .B1(new_n1310), .B2(new_n1325), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1320), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(new_n1290), .A3(new_n1318), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1305), .B1(new_n1327), .B2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1299), .A2(new_n1321), .A3(new_n1303), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1310), .A2(KEYINPUT63), .A3(new_n1318), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT125), .B1(new_n1328), .B2(new_n1290), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT125), .ZN(new_n1338));
  AOI211_X1 g1138(.A(new_n1338), .B(new_n1291), .C1(new_n1306), .C2(new_n1309), .ZN(new_n1339));
  NOR3_X1   g1139(.A1(new_n1337), .A2(new_n1339), .A3(new_n1325), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1336), .A2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1294), .B1(new_n1331), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1319), .ZN(new_n1343));
  OAI221_X1 g1143(.A(new_n1321), .B1(new_n1310), .B2(new_n1325), .C1(new_n1329), .C2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1330), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1304), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1325), .B1(new_n1310), .B2(KEYINPUT125), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1347), .B1(KEYINPUT125), .B2(new_n1310), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1348), .A2(new_n1335), .A3(new_n1333), .A4(new_n1334), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1346), .A2(KEYINPUT127), .A3(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1342), .A2(new_n1350), .ZN(G405));
  NOR2_X1   g1151(.A1(new_n1281), .A2(G378), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1306), .ZN(new_n1353));
  OR3_X1    g1153(.A1(new_n1352), .A2(new_n1353), .A3(new_n1318), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1318), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1304), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1354), .A2(new_n1305), .A3(new_n1355), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(G402));
endmodule


