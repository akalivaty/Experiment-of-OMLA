//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT82), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(KEYINPUT22), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(KEYINPUT22), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(G204gat), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(G204gat), .B1(new_n210), .B2(new_n211), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G211gat), .B(G218gat), .Z(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT75), .B(G197gat), .ZN(new_n218));
  INV_X1    g017(.A(G204gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n212), .ZN(new_n221));
  INV_X1    g020(.A(new_n216), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(new_n209), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G226gat), .A2(G233gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT24), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NOR3_X1   g038(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n228), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245));
  INV_X1    g044(.A(G169gat), .ZN(new_n246));
  INV_X1    g045(.A(G176gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n238), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n249), .A2(new_n233), .A3(new_n237), .A4(new_n235), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT65), .A3(new_n228), .ZN(new_n251));
  NOR2_X1   g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(new_n234), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n232), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT24), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n248), .A2(new_n238), .B1(G169gat), .B2(G176gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n251), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT67), .B1(new_n229), .B2(KEYINPUT27), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n230), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n263), .A2(KEYINPUT28), .A3(new_n230), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OR3_X1    g068(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n237), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n232), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n227), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n226), .B1(new_n261), .B2(new_n273), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n225), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  INV_X1    g078(.A(G64gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G92gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n274), .A2(new_n227), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT29), .B1(new_n261), .B2(new_n273), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n285), .B(new_n224), .C1(new_n227), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n278), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n288), .A2(KEYINPUT77), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT77), .B1(new_n288), .B2(new_n289), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n284), .B1(new_n278), .B2(new_n287), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n278), .A2(new_n284), .A3(new_n287), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(KEYINPUT30), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n203), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n288), .A2(new_n289), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n288), .A2(KEYINPUT77), .A3(new_n289), .ZN(new_n300));
  AND4_X1   g099(.A1(new_n203), .A2(new_n295), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n202), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G127gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G134gat), .ZN(new_n304));
  INV_X1    g103(.A(G134gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G127gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT68), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(new_n303), .B2(G134gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT69), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G134gat), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n311), .B(new_n312), .C1(new_n313), .C2(KEYINPUT68), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G113gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G120gat), .ZN(new_n317));
  INV_X1    g116(.A(G120gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G113gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT71), .B1(new_n318), .B2(G113gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(new_n316), .A3(G120gat), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n319), .A2(KEYINPUT70), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT70), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n318), .A3(G113gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT1), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT72), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n313), .B(new_n332), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n315), .A2(new_n322), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n250), .A2(KEYINPUT65), .A3(new_n228), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT65), .B1(new_n250), .B2(new_n228), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n259), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n232), .ZN(new_n340));
  INV_X1    g139(.A(new_n272), .ZN(new_n341));
  AOI211_X1 g140(.A(new_n340), .B(new_n341), .C1(new_n267), .C2(new_n268), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n335), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n344), .B(KEYINPUT64), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n261), .A2(new_n273), .A3(new_n334), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n348), .B(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G15gat), .B(G43gat), .Z(new_n352));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n346), .B1(new_n343), .B2(new_n347), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(KEYINPUT33), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT32), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n347), .ZN(new_n360));
  AOI221_X4 g159(.A(new_n357), .B1(KEYINPUT33), .B2(new_n354), .C1(new_n360), .C2(new_n345), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n351), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n261), .A2(new_n334), .A3(new_n273), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n334), .B1(new_n261), .B2(new_n273), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n345), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT32), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n354), .C1(KEYINPUT33), .C2(new_n355), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n356), .A2(new_n358), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n348), .B(new_n349), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n362), .A2(KEYINPUT74), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n367), .A2(new_n368), .A3(new_n369), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G57gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(G85gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT5), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382));
  OR2_X1    g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(KEYINPUT2), .ZN(new_n384));
  INV_X1    g183(.A(G148gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G141gat), .ZN(new_n386));
  INV_X1    g185(.A(G141gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G148gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n386), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n384), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n386), .A2(new_n388), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n382), .B(new_n383), .C1(new_n393), .C2(KEYINPUT2), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n335), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n315), .A2(new_n322), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n392), .A2(new_n394), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n331), .A2(new_n333), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n381), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n381), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(KEYINPUT3), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n392), .A2(new_n394), .A3(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n310), .A2(new_n314), .B1(new_n321), .B2(new_n320), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n328), .B1(G113gat), .B2(new_n318), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n316), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n323), .B(new_n325), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n321), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n313), .B(KEYINPUT72), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n403), .B(new_n405), .C1(new_n406), .C2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n402), .B1(new_n415), .B2(new_n400), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n412), .A2(new_n406), .A3(new_n395), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT4), .ZN(new_n418));
  AOI211_X1 g217(.A(new_n380), .B(new_n401), .C1(new_n416), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT80), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n400), .A2(new_n414), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n400), .A2(new_n423), .A3(KEYINPUT4), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(new_n380), .A3(new_n381), .A4(new_n413), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n379), .B1(new_n419), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n416), .A2(new_n418), .ZN(new_n430));
  INV_X1    g229(.A(new_n401), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(KEYINPUT5), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(new_n426), .A3(new_n378), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n428), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT6), .B(new_n379), .C1(new_n419), .C2(new_n427), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT31), .B(G50gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(G228gat), .A2(G233gat), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT29), .B1(new_n217), .B2(new_n223), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n404), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI211_X1 g240(.A(KEYINPUT81), .B(KEYINPUT29), .C1(new_n217), .C2(new_n223), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n395), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n405), .A2(new_n275), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n225), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n438), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n439), .A2(new_n395), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n445), .A2(new_n447), .A3(new_n403), .A4(new_n438), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n437), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G78gat), .B(G106gat), .Z(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(G22gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n437), .ZN(new_n453));
  INV_X1    g252(.A(new_n445), .ZN(new_n454));
  INV_X1    g253(.A(new_n223), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n222), .B1(new_n221), .B2(new_n209), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n275), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT81), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n440), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n404), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n454), .B1(new_n460), .B2(new_n395), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n453), .B(new_n448), .C1(new_n461), .C2(new_n438), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n450), .A2(new_n452), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n452), .B1(new_n450), .B2(new_n462), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n374), .A2(new_n436), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT85), .B1(new_n302), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n295), .A2(new_n299), .A3(new_n300), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT82), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n292), .A2(new_n203), .A3(new_n295), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT35), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n463), .A2(new_n464), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n373), .B2(new_n371), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n471), .A2(new_n472), .A3(new_n474), .A4(new_n436), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n468), .B1(new_n435), .B2(new_n434), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n370), .B(new_n362), .C1(new_n463), .C2(new_n464), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n202), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n362), .A2(KEYINPUT36), .A3(new_n370), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n374), .B2(KEYINPUT36), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n378), .B1(new_n432), .B2(new_n426), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n425), .A2(new_n413), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n402), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT40), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n378), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n396), .A2(new_n381), .A3(new_n400), .ZN(new_n492));
  AOI211_X1 g291(.A(new_n487), .B(new_n492), .C1(new_n486), .C2(new_n402), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n485), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n491), .A2(new_n493), .B1(KEYINPUT83), .B2(new_n489), .ZN(new_n497));
  AND4_X1   g296(.A1(new_n469), .A2(new_n496), .A3(new_n470), .A4(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n278), .B2(new_n287), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n278), .A2(new_n499), .A3(new_n287), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n283), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT38), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n500), .A2(new_n501), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n502), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT38), .B1(new_n504), .B2(new_n500), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n288), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n465), .B1(new_n510), .B2(new_n436), .ZN(new_n511));
  OAI221_X1 g310(.A(new_n484), .B1(new_n477), .B2(new_n465), .C1(new_n498), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n482), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  NOR2_X1   g313(.A1(G29gat), .A2(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT86), .B1(G29gat), .B2(G36gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n517), .B(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G43gat), .B(G50gat), .Z(new_n521));
  INV_X1    g320(.A(KEYINPUT15), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G29gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT87), .B(G36gat), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n520), .B(new_n523), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n521), .A2(new_n522), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n528), .A2(KEYINPUT17), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT88), .ZN(new_n531));
  INV_X1    g330(.A(G1gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n532), .A2(KEYINPUT16), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(new_n531), .ZN(new_n535));
  INV_X1    g334(.A(G8gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n528), .A2(KEYINPUT17), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n529), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n537), .A2(new_n528), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n537), .A2(new_n528), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(new_n540), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n542), .B(KEYINPUT13), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n539), .A2(KEYINPUT18), .A3(new_n541), .A4(new_n542), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT11), .B(G169gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G197gat), .ZN(new_n553));
  XOR2_X1   g352(.A(G113gat), .B(G141gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT12), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n545), .A2(new_n549), .A3(new_n556), .A4(new_n550), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G64gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n280), .A2(G57gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(KEYINPUT9), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G71gat), .ZN(new_n570));
  INV_X1    g369(.A(G78gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT89), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n567), .B(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT90), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n569), .A2(KEYINPUT90), .A3(new_n572), .A4(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n572), .A2(new_n567), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n566), .B(new_n580), .C1(KEYINPUT9), .C2(new_n568), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT91), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT93), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(G99gat), .A3(G106gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n588), .A3(KEYINPUT8), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT94), .B(G85gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(G92gat), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT95), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n589), .B(new_n593), .C1(G92gat), .C2(new_n590), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G99gat), .B(G106gat), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT96), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT7), .B1(new_n598), .B2(KEYINPUT92), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(KEYINPUT92), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(KEYINPUT92), .A3(KEYINPUT7), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n595), .A2(new_n597), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n596), .A2(KEYINPUT96), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n592), .A2(new_n594), .B1(new_n601), .B2(new_n602), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(new_n597), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n584), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n579), .A2(new_n583), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n604), .A2(new_n605), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n608), .A2(new_n607), .A3(new_n597), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT10), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n613), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n562), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n562), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n610), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT98), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n318), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n619), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n619), .A2(new_n629), .A3(new_n621), .A4(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n619), .A2(new_n621), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n625), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n561), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n606), .A2(new_n609), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n528), .ZN(new_n637));
  AND3_X1   g436(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n529), .A2(new_n636), .A3(new_n538), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  XNOR2_X1  g443(.A(G190gat), .B(G218gat), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OR3_X1    g447(.A1(new_n643), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n643), .B2(new_n644), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G127gat), .B(G155gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n207), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n537), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(G183gat), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(G183gat), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(G231gat), .A3(G233gat), .A4(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  INV_X1    g461(.A(G231gat), .ZN(new_n663));
  INV_X1    g462(.A(G233gat), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n662), .A2(new_n658), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n655), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n661), .A2(new_n665), .A3(new_n655), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n670), .ZN(new_n673));
  INV_X1    g472(.A(new_n671), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(new_n666), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n652), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT97), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n652), .A2(new_n676), .A3(KEYINPUT97), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n513), .A2(new_n635), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n436), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n532), .ZN(G1324gat));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n296), .A2(new_n301), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n682), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n685), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G8gat), .B1(new_n682), .B2(new_n687), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n689), .A2(KEYINPUT100), .A3(KEYINPUT42), .A4(new_n690), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT101), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n693), .A2(new_n700), .A3(new_n696), .A4(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(G1325gat));
  INV_X1    g501(.A(G15gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n484), .B(KEYINPUT102), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n682), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n374), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n682), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(new_n703), .B2(new_n708), .ZN(G1326gat));
  NOR2_X1   g508(.A1(new_n682), .A2(new_n465), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT43), .B(G22gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  AOI21_X1  g511(.A(new_n652), .B1(new_n482), .B2(new_n512), .ZN(new_n713));
  INV_X1    g512(.A(new_n676), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n635), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(G29gat), .A3(new_n436), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n484), .B1(new_n498), .B2(new_n511), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n477), .B2(new_n465), .ZN(new_n724));
  INV_X1    g523(.A(new_n468), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n436), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(KEYINPUT104), .A3(new_n473), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n480), .B1(new_n467), .B2(new_n475), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n721), .B(new_n651), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n713), .B2(new_n721), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n716), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n436), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT105), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n720), .B1(new_n735), .B2(new_n524), .ZN(G1328gat));
  INV_X1    g535(.A(new_n717), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(new_n525), .A3(new_n686), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT46), .Z(new_n739));
  NOR2_X1   g538(.A1(new_n733), .A2(new_n687), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n525), .B2(new_n740), .ZN(G1329gat));
  OAI21_X1  g540(.A(G43gat), .B1(new_n733), .B2(new_n484), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n717), .A2(G43gat), .A3(new_n707), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(KEYINPUT47), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G43gat), .B1(new_n733), .B2(new_n705), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(new_n743), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n746), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  INV_X1    g547(.A(G50gat), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n477), .A2(new_n465), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n722), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n730), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT44), .B1(new_n752), .B2(new_n652), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n715), .B1(new_n753), .B2(new_n731), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n749), .B1(new_n754), .B2(new_n473), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n473), .A2(new_n749), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n717), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n755), .A2(KEYINPUT106), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n759));
  OAI21_X1  g558(.A(G50gat), .B1(new_n733), .B2(new_n465), .ZN(new_n760));
  INV_X1    g559(.A(new_n757), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n748), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT106), .B1(new_n755), .B2(new_n757), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n759), .A3(new_n761), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(KEYINPUT48), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(G1331gat));
  AND2_X1   g566(.A1(new_n681), .A2(new_n561), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n469), .A2(new_n496), .A3(new_n470), .A4(new_n497), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n769), .B(new_n465), .C1(new_n436), .C2(new_n510), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(new_n484), .A3(new_n724), .A4(new_n727), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n482), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n768), .A2(new_n634), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n436), .B(KEYINPUT107), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n563), .ZN(G1332gat));
  NOR2_X1   g576(.A1(new_n773), .A2(new_n687), .ZN(new_n778));
  NOR2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  AND2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n778), .B2(new_n779), .ZN(G1333gat));
  AND2_X1   g581(.A1(new_n768), .A2(new_n772), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n783), .A2(G71gat), .A3(new_n634), .A4(new_n704), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n570), .B1(new_n773), .B2(new_n707), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n784), .A2(new_n786), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT108), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT50), .B1(new_n793), .B2(new_n787), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n791), .A2(new_n794), .ZN(G1334gat));
  NOR2_X1   g594(.A1(new_n773), .A2(new_n465), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT109), .B(G78gat), .Z(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1335gat));
  NOR2_X1   g597(.A1(new_n676), .A2(new_n560), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n732), .A2(new_n634), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g599(.A(KEYINPUT94), .B(G85gat), .Z(new_n801));
  NOR3_X1   g600(.A1(new_n800), .A2(new_n436), .A3(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n651), .B(new_n799), .C1(new_n729), .C2(new_n730), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n651), .A4(new_n799), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n634), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n436), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n802), .B1(new_n811), .B2(new_n801), .ZN(G1336gat));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n652), .B1(new_n482), .B2(new_n771), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT51), .B1(new_n814), .B2(new_n799), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n803), .A2(new_n804), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n813), .B1(new_n803), .B2(new_n804), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n687), .A2(G92gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n634), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G92gat), .B1(new_n800), .B2(new_n687), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT52), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n809), .A2(KEYINPUT111), .A3(new_n821), .ZN(new_n826));
  XNOR2_X1  g625(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n828));
  INV_X1    g627(.A(new_n821), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n808), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n826), .A2(new_n823), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n825), .A2(new_n831), .ZN(G1337gat));
  OAI21_X1  g631(.A(G99gat), .B1(new_n800), .B2(new_n705), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n808), .A2(G99gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n707), .ZN(G1338gat));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n732), .A2(new_n634), .A3(new_n473), .A4(new_n799), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(G106gat), .ZN(new_n838));
  INV_X1    g637(.A(new_n634), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n839), .A2(G106gat), .A3(new_n465), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT53), .B1(new_n807), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n820), .A2(new_n840), .B1(G106gat), .B2(new_n837), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n836), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT110), .B1(new_n805), .B2(new_n806), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n846), .B2(new_n818), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n838), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n838), .A2(new_n841), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT113), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n845), .A2(new_n850), .ZN(G1339gat));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT10), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n606), .A2(new_n609), .A3(new_n584), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n611), .B1(new_n613), .B2(new_n612), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n617), .A3(new_n620), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n857), .A2(new_n619), .A3(KEYINPUT54), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n625), .B1(new_n619), .B2(KEYINPUT54), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n852), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n620), .B1(new_n856), .B2(new_n617), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n626), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n857), .A2(new_n619), .A3(KEYINPUT54), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(KEYINPUT55), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n631), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT114), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n860), .A2(new_n631), .A3(new_n868), .A4(new_n865), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n560), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n547), .A2(new_n548), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n542), .B1(new_n539), .B2(new_n541), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n555), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n634), .A2(new_n559), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n651), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n559), .A2(new_n873), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n649), .B2(new_n650), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n867), .A2(new_n877), .A3(new_n869), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n714), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n679), .A2(new_n839), .A3(new_n561), .A4(new_n680), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n686), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(new_n479), .A3(new_n774), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n316), .A3(new_n560), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n810), .A3(new_n474), .ZN(new_n885));
  OAI21_X1  g684(.A(G113gat), .B1(new_n885), .B2(new_n561), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT115), .Z(G1340gat));
  NAND3_X1  g687(.A1(new_n883), .A2(new_n318), .A3(new_n634), .ZN(new_n889));
  OAI21_X1  g688(.A(G120gat), .B1(new_n885), .B2(new_n839), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1341gat));
  NOR3_X1   g690(.A1(new_n885), .A2(new_n303), .A3(new_n714), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n883), .A2(new_n676), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT116), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n894), .B2(new_n303), .ZN(G1342gat));
  NAND4_X1  g694(.A1(new_n883), .A2(KEYINPUT56), .A3(new_n305), .A4(new_n651), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n305), .A3(new_n479), .A4(new_n774), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n652), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n882), .A2(new_n810), .A3(new_n651), .A4(new_n474), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(G134gat), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n901), .B2(G134gat), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT118), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n896), .A2(new_n899), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n907), .B(new_n908), .C1(new_n904), .C2(new_n903), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n909), .ZN(G1343gat));
  AND2_X1   g709(.A1(new_n866), .A2(KEYINPUT119), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n560), .B1(new_n866), .B2(KEYINPUT119), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n874), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n652), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n676), .B1(new_n914), .B2(new_n878), .ZN(new_n915));
  INV_X1    g714(.A(new_n881), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n473), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT57), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n880), .A2(new_n881), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n473), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n687), .A2(new_n810), .A3(new_n484), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G141gat), .B1(new_n923), .B2(new_n561), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n882), .A2(new_n774), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n704), .A2(new_n465), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n925), .A2(new_n387), .A3(new_n560), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT58), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT58), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n924), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1344gat));
  AND2_X1   g731(.A1(new_n925), .A2(new_n926), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n385), .A3(new_n634), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n935));
  AOI211_X1 g734(.A(KEYINPUT59), .B(new_n385), .C1(new_n935), .C2(new_n634), .ZN(new_n936));
  XOR2_X1   g735(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n937));
  AND2_X1   g736(.A1(new_n880), .A2(new_n881), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT57), .B1(new_n938), .B2(new_n465), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n877), .A2(new_n631), .A3(new_n860), .A4(new_n865), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n676), .B1(new_n914), .B2(new_n940), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n920), .B(new_n473), .C1(new_n941), .C2(new_n916), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n939), .A2(new_n634), .A3(new_n922), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n937), .B1(new_n943), .B2(G148gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n934), .B1(new_n936), .B2(new_n944), .ZN(G1345gat));
  AOI21_X1  g744(.A(G155gat), .B1(new_n933), .B2(new_n676), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n676), .A2(G155gat), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT121), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n935), .B2(new_n948), .ZN(G1346gat));
  OAI21_X1  g748(.A(G162gat), .B1(new_n923), .B2(new_n652), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n951));
  INV_X1    g750(.A(G162gat), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n925), .A2(new_n952), .A3(new_n651), .A4(new_n926), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n950), .B2(new_n953), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(new_n955), .ZN(G1347gat));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n810), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n686), .A2(new_n479), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT123), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n960), .A2(G169gat), .A3(new_n561), .ZN(new_n961));
  INV_X1    g760(.A(new_n474), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n880), .B2(new_n881), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n774), .A2(new_n687), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n246), .B1(new_n965), .B2(new_n560), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n961), .A2(new_n966), .ZN(G1348gat));
  OAI21_X1  g766(.A(new_n247), .B1(new_n960), .B2(new_n839), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n965), .A2(G176gat), .A3(new_n634), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n968), .A2(new_n969), .ZN(G1349gat));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(KEYINPUT60), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n971), .A2(KEYINPUT60), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n963), .A2(new_n676), .A3(new_n964), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n963), .A2(new_n976), .A3(new_n676), .A4(new_n964), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n975), .A2(G183gat), .A3(new_n977), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n957), .A2(new_n676), .A3(new_n263), .A4(new_n959), .ZN(new_n979));
  AOI211_X1 g778(.A(new_n972), .B(new_n973), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  AND4_X1   g779(.A1(new_n971), .A2(new_n978), .A3(KEYINPUT60), .A4(new_n979), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n980), .A2(new_n981), .ZN(G1350gat));
  AOI21_X1  g781(.A(new_n230), .B1(new_n965), .B2(new_n651), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT61), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n960), .A2(G190gat), .A3(new_n652), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(new_n985), .ZN(G1351gat));
  NAND2_X1  g785(.A1(new_n939), .A2(new_n942), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n939), .A2(KEYINPUT126), .A3(new_n942), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n705), .A2(new_n964), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(G197gat), .B1(new_n993), .B2(new_n561), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n957), .A2(new_n686), .A3(new_n926), .ZN(new_n995));
  INV_X1    g794(.A(G197gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n995), .A2(new_n996), .A3(new_n560), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n994), .A2(new_n997), .ZN(G1352gat));
  OAI21_X1  g797(.A(G204gat), .B1(new_n993), .B2(new_n839), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n995), .A2(new_n1000), .A3(new_n219), .A4(new_n634), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n957), .A2(new_n219), .A3(new_n686), .A4(new_n926), .ZN(new_n1002));
  OAI21_X1  g801(.A(KEYINPUT62), .B1(new_n1002), .B2(new_n839), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n999), .A2(new_n1004), .ZN(G1353gat));
  NAND4_X1  g804(.A1(new_n939), .A2(new_n676), .A3(new_n942), .A4(new_n992), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G211gat), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT63), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(KEYINPUT63), .ZN(new_n1010));
  OR2_X1    g809(.A1(new_n1008), .A2(KEYINPUT63), .ZN(new_n1011));
  NAND4_X1  g810(.A1(new_n1006), .A2(G211gat), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n995), .A2(new_n207), .A3(new_n676), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .ZN(G1354gat));
  OAI21_X1  g813(.A(G218gat), .B1(new_n993), .B2(new_n652), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n995), .A2(new_n208), .A3(new_n651), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(G1355gat));
endmodule


