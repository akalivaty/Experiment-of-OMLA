

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  XOR2_X1 U325 ( .A(n447), .B(KEYINPUT79), .Z(n293) );
  INV_X1 U326 ( .A(KEYINPUT95), .ZN(n350) );
  XNOR2_X1 U327 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U328 ( .A(n370), .B(n352), .ZN(n356) );
  XNOR2_X1 U329 ( .A(KEYINPUT106), .B(KEYINPUT37), .ZN(n420) );
  XNOR2_X1 U330 ( .A(n421), .B(n420), .ZN(n526) );
  XOR2_X1 U331 ( .A(KEYINPUT36), .B(n562), .Z(n590) );
  INV_X1 U332 ( .A(KEYINPUT58), .ZN(n481) );
  XOR2_X1 U333 ( .A(n309), .B(n308), .Z(n562) );
  XNOR2_X1 U334 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U335 ( .A(n456), .B(KEYINPUT110), .ZN(n457) );
  XNOR2_X1 U336 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n458), .B(n457), .ZN(G1331GAT) );
  XOR2_X1 U338 ( .A(G162GAT), .B(G50GAT), .Z(n334) );
  XOR2_X1 U339 ( .A(G43GAT), .B(KEYINPUT7), .Z(n295) );
  XNOR2_X1 U340 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n427) );
  XNOR2_X1 U342 ( .A(n334), .B(n427), .ZN(n296) );
  XOR2_X1 U343 ( .A(G190GAT), .B(G36GAT), .Z(n347) );
  XNOR2_X1 U344 ( .A(n296), .B(n347), .ZN(n301) );
  XOR2_X1 U345 ( .A(G92GAT), .B(G99GAT), .Z(n298) );
  XNOR2_X1 U346 ( .A(G85GAT), .B(KEYINPUT75), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n447) );
  NAND2_X1 U348 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n293), .B(n299), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n309) );
  XOR2_X1 U351 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n303) );
  XNOR2_X1 U352 ( .A(G134GAT), .B(G218GAT), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U354 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n305) );
  XNOR2_X1 U355 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U357 ( .A(n307), .B(n306), .Z(n308) );
  XOR2_X1 U358 ( .A(G22GAT), .B(G211GAT), .Z(n311) );
  XNOR2_X1 U359 ( .A(G71GAT), .B(G183GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U361 ( .A(n312), .B(G78GAT), .Z(n314) );
  XOR2_X1 U362 ( .A(G127GAT), .B(G15GAT), .Z(n365) );
  XNOR2_X1 U363 ( .A(G155GAT), .B(n365), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n314), .B(n313), .ZN(n319) );
  XNOR2_X1 U365 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n315), .B(KEYINPUT13), .ZN(n446) );
  XOR2_X1 U367 ( .A(n446), .B(KEYINPUT12), .Z(n317) );
  NAND2_X1 U368 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U370 ( .A(n319), .B(n318), .Z(n327) );
  XOR2_X1 U371 ( .A(KEYINPUT14), .B(G8GAT), .Z(n321) );
  XNOR2_X1 U372 ( .A(G1GAT), .B(G64GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U374 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n323) );
  XNOR2_X1 U375 ( .A(KEYINPUT82), .B(KEYINPUT81), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U378 ( .A(n327), .B(n326), .Z(n485) );
  INV_X1 U379 ( .A(n485), .ZN(n584) );
  XNOR2_X1 U380 ( .A(G78GAT), .B(KEYINPUT73), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n328), .B(KEYINPUT74), .ZN(n329) );
  XOR2_X1 U382 ( .A(n329), .B(G204GAT), .Z(n331) );
  XNOR2_X1 U383 ( .A(G148GAT), .B(G106GAT), .ZN(n330) );
  XOR2_X1 U384 ( .A(n331), .B(n330), .Z(n452) );
  XOR2_X1 U385 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n333) );
  XNOR2_X1 U386 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U388 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n336) );
  XOR2_X1 U389 ( .A(G141GAT), .B(G22GAT), .Z(n424) );
  XNOR2_X1 U390 ( .A(n334), .B(n424), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n340) );
  AND2_X1 U393 ( .A1(G228GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n345) );
  XNOR2_X1 U395 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n341), .B(KEYINPUT2), .ZN(n406) );
  XOR2_X1 U397 ( .A(G197GAT), .B(KEYINPUT21), .Z(n343) );
  XNOR2_X1 U398 ( .A(G218GAT), .B(G211GAT), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n358) );
  XNOR2_X1 U400 ( .A(n406), .B(n358), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U402 ( .A(n452), .B(n346), .Z(n476) );
  XOR2_X1 U403 ( .A(G8GAT), .B(G169GAT), .Z(n426) );
  XNOR2_X1 U404 ( .A(n347), .B(n426), .ZN(n362) );
  XOR2_X1 U405 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n349) );
  XNOR2_X1 U406 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n370) );
  NAND2_X1 U408 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XOR2_X1 U409 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n354) );
  XNOR2_X1 U410 ( .A(G92GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U412 ( .A(n356), .B(n355), .Z(n360) );
  XNOR2_X1 U413 ( .A(G64GAT), .B(G176GAT), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n357), .B(KEYINPUT76), .ZN(n439) );
  XNOR2_X1 U415 ( .A(n358), .B(n439), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U417 ( .A(n362), .B(n361), .Z(n471) );
  INV_X1 U418 ( .A(n471), .ZN(n507) );
  XOR2_X1 U419 ( .A(G176GAT), .B(KEYINPUT84), .Z(n364) );
  XNOR2_X1 U420 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n380) );
  XOR2_X1 U422 ( .A(G120GAT), .B(G71GAT), .Z(n440) );
  XOR2_X1 U423 ( .A(n440), .B(n365), .Z(n367) );
  XNOR2_X1 U424 ( .A(G99GAT), .B(G43GAT), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n376) );
  XOR2_X1 U426 ( .A(G113GAT), .B(KEYINPUT0), .Z(n369) );
  XNOR2_X1 U427 ( .A(G134GAT), .B(KEYINPUT83), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n407) );
  XNOR2_X1 U429 ( .A(n407), .B(n370), .ZN(n374) );
  XOR2_X1 U430 ( .A(G169GAT), .B(KEYINPUT66), .Z(n372) );
  XNOR2_X1 U431 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U434 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U435 ( .A1(G227GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U437 ( .A(n380), .B(n379), .Z(n383) );
  INV_X1 U438 ( .A(n383), .ZN(n511) );
  NOR2_X1 U439 ( .A1(n507), .A2(n511), .ZN(n381) );
  NOR2_X1 U440 ( .A1(n476), .A2(n381), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n382), .B(KEYINPUT25), .ZN(n389) );
  INV_X1 U442 ( .A(n476), .ZN(n384) );
  OR2_X1 U443 ( .A1(n384), .A2(n383), .ZN(n386) );
  INV_X1 U444 ( .A(KEYINPUT26), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n551) );
  XNOR2_X1 U446 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n387) );
  XOR2_X1 U447 ( .A(n387), .B(n507), .Z(n412) );
  NAND2_X1 U448 ( .A1(n551), .A2(n412), .ZN(n388) );
  NAND2_X1 U449 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n390), .B(KEYINPUT98), .ZN(n410) );
  XOR2_X1 U451 ( .A(G127GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U452 ( .A(G29GAT), .B(G85GAT), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U454 ( .A(KEYINPUT4), .B(G141GAT), .Z(n394) );
  XNOR2_X1 U455 ( .A(G120GAT), .B(G148GAT), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U457 ( .A(n396), .B(n395), .Z(n401) );
  XOR2_X1 U458 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n398) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U461 ( .A(KEYINPUT5), .B(n399), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U463 ( .A(KEYINPUT92), .B(KEYINPUT1), .Z(n403) );
  XNOR2_X1 U464 ( .A(KEYINPUT91), .B(G57GAT), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U466 ( .A(n405), .B(n404), .Z(n409) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n491) );
  XOR2_X1 U469 ( .A(G1GAT), .B(n491), .Z(n527) );
  INV_X1 U470 ( .A(n527), .ZN(n504) );
  NAND2_X1 U471 ( .A1(n410), .A2(n504), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n411), .B(KEYINPUT99), .ZN(n416) );
  NAND2_X1 U473 ( .A1(n412), .A2(n527), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n413), .B(KEYINPUT97), .ZN(n538) );
  XOR2_X1 U475 ( .A(n476), .B(KEYINPUT28), .Z(n539) );
  NAND2_X1 U476 ( .A1(n538), .A2(n539), .ZN(n414) );
  INV_X1 U477 ( .A(n511), .ZN(n540) );
  NOR2_X1 U478 ( .A1(n414), .A2(n540), .ZN(n415) );
  NOR2_X1 U479 ( .A1(n416), .A2(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n417), .B(KEYINPUT100), .ZN(n488) );
  NOR2_X1 U481 ( .A1(n584), .A2(n488), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n418), .B(KEYINPUT105), .ZN(n419) );
  NOR2_X1 U483 ( .A1(n590), .A2(n419), .ZN(n421) );
  XOR2_X1 U484 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n423) );
  XNOR2_X1 U485 ( .A(G1GAT), .B(G197GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U487 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U490 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n431) );
  NAND2_X1 U491 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U493 ( .A(n433), .B(n432), .Z(n438) );
  XOR2_X1 U494 ( .A(G15GAT), .B(G36GAT), .Z(n435) );
  XNOR2_X1 U495 ( .A(G113GAT), .B(G50GAT), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n436), .B(KEYINPUT30), .ZN(n437) );
  XOR2_X1 U498 ( .A(n438), .B(n437), .Z(n515) );
  INV_X1 U499 ( .A(n515), .ZN(n575) );
  XOR2_X1 U500 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n442) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n451) );
  XOR2_X1 U503 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n444) );
  NAND2_X1 U504 ( .A1(G230GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U505 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U506 ( .A(n445), .B(KEYINPUT77), .Z(n449) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n581) );
  NAND2_X1 U511 ( .A1(n575), .A2(n581), .ZN(n489) );
  NOR2_X1 U512 ( .A1(n526), .A2(n489), .ZN(n455) );
  XNOR2_X1 U513 ( .A(KEYINPUT38), .B(KEYINPUT107), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n455), .B(n454), .ZN(n512) );
  NOR2_X1 U515 ( .A1(n512), .A2(n539), .ZN(n458) );
  INV_X1 U516 ( .A(G50GAT), .ZN(n456) );
  XOR2_X1 U517 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n480) );
  XNOR2_X1 U518 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n473) );
  INV_X1 U519 ( .A(n562), .ZN(n462) );
  XNOR2_X1 U520 ( .A(KEYINPUT41), .B(n581), .ZN(n555) );
  NAND2_X1 U521 ( .A1(n575), .A2(n555), .ZN(n459) );
  XOR2_X1 U522 ( .A(KEYINPUT46), .B(n459), .Z(n460) );
  NOR2_X1 U523 ( .A1(n584), .A2(n460), .ZN(n461) );
  NAND2_X1 U524 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n463), .B(KEYINPUT47), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n590), .A2(n485), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n464), .B(KEYINPUT45), .ZN(n465) );
  NAND2_X1 U528 ( .A1(n465), .A2(n581), .ZN(n466) );
  NOR2_X1 U529 ( .A1(n466), .A2(n575), .ZN(n467) );
  NOR2_X1 U530 ( .A1(n468), .A2(n467), .ZN(n470) );
  XOR2_X1 U531 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n469) );
  XNOR2_X1 U532 ( .A(n470), .B(n469), .ZN(n537) );
  NAND2_X1 U533 ( .A1(n537), .A2(n471), .ZN(n472) );
  XOR2_X1 U534 ( .A(n473), .B(n472), .Z(n474) );
  NOR2_X1 U535 ( .A1(n527), .A2(n474), .ZN(n475) );
  XNOR2_X1 U536 ( .A(KEYINPUT65), .B(n475), .ZN(n573) );
  NOR2_X1 U537 ( .A1(n476), .A2(n573), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n477), .B(KEYINPUT55), .ZN(n478) );
  NOR2_X2 U539 ( .A1(n511), .A2(n478), .ZN(n570) );
  NAND2_X1 U540 ( .A1(n570), .A2(n562), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(n484) );
  XNOR2_X1 U542 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n482) );
  NOR2_X1 U543 ( .A1(n562), .A2(n485), .ZN(n486) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(n486), .Z(n487) );
  OR2_X1 U545 ( .A1(n488), .A2(n487), .ZN(n516) );
  NOR2_X1 U546 ( .A1(n489), .A2(n516), .ZN(n500) );
  INV_X1 U547 ( .A(n500), .ZN(n490) );
  NOR2_X1 U548 ( .A1(n491), .A2(n490), .ZN(n493) );
  NOR2_X1 U549 ( .A1(G1GAT), .A2(n500), .ZN(n492) );
  NOR2_X1 U550 ( .A1(n493), .A2(n492), .ZN(n495) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n494) );
  XNOR2_X1 U552 ( .A(n495), .B(n494), .ZN(G1324GAT) );
  NAND2_X1 U553 ( .A1(n471), .A2(n500), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n496), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n498) );
  NAND2_X1 U556 ( .A1(n500), .A2(n540), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n502) );
  INV_X1 U560 ( .A(n539), .ZN(n532) );
  NAND2_X1 U561 ( .A1(n500), .A2(n532), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G22GAT), .B(n503), .ZN(G1327GAT) );
  NOR2_X1 U564 ( .A1(n512), .A2(n504), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n507), .A2(n512), .ZN(n508) );
  XOR2_X1 U568 ( .A(G36GAT), .B(n508), .Z(G1329GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n510) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n512), .A2(n511), .ZN(n513) );
  XOR2_X1 U573 ( .A(n514), .B(n513), .Z(G1330GAT) );
  XOR2_X1 U574 ( .A(n555), .B(KEYINPUT111), .Z(n566) );
  NAND2_X1 U575 ( .A1(n566), .A2(n515), .ZN(n525) );
  NOR2_X1 U576 ( .A1(n525), .A2(n516), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n527), .A2(n522), .ZN(n517) );
  XNOR2_X1 U578 ( .A(KEYINPUT42), .B(n517), .ZN(n518) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U580 ( .A1(n471), .A2(n522), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n522), .A2(n540), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n520), .B(KEYINPUT112), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G71GAT), .B(n521), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U586 ( .A1(n522), .A2(n532), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  XOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT113), .Z(n529) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n471), .A2(n533), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n533), .A2(n540), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n535) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U599 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  NAND2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n552) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U602 ( .A1(n552), .A2(n541), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n575), .A2(n548), .ZN(n542) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U606 ( .A1(n548), .A2(n566), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n545), .Z(G1341GAT) );
  NAND2_X1 U609 ( .A1(n548), .A2(n584), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U613 ( .A1(n548), .A2(n562), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n554) );
  INV_X1 U616 ( .A(n551), .ZN(n574) );
  NOR2_X1 U617 ( .A1(n574), .A2(n552), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n575), .A2(n561), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U621 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT117), .Z(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n584), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(KEYINPUT118), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n575), .A2(n570), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n570), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n584), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT120), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G183GAT), .B(n572), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n577) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n585), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(n578), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U647 ( .A(n585), .ZN(n589) );
  OR2_X1 U648 ( .A1(n589), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n588) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(n592), .B(n591), .Z(G1355GAT) );
endmodule

