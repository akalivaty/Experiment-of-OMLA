//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G125), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT68), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n466), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n467), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n478), .A2(new_n479), .A3(new_n465), .A4(new_n470), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n469), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(G137), .B1(G101), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(G112), .B2(new_n465), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n481), .A2(G136), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n478), .A2(new_n479), .A3(G2105), .A4(new_n470), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n478), .A2(new_n479), .A3(new_n496), .A4(new_n470), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n463), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(G114), .B2(new_n465), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n492), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n499), .A2(new_n504), .ZN(G164));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OAI211_X1 g082(.A(G50), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT71), .A2(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT71), .A2(G88), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n509), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n508), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n510), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n510), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n522), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n515), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n524), .A2(new_n523), .B1(new_n506), .B2(new_n507), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n520), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n515), .ZN(new_n538));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT72), .B(G81), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n520), .A2(new_n539), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NOR2_X1   g122(.A1(new_n506), .A2(new_n507), .ZN(new_n548));
  INV_X1    g123(.A(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(KEYINPUT73), .A3(G53), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n520), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n554), .A3(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n552), .B(new_n556), .C1(new_n520), .C2(new_n553), .ZN(new_n557));
  INV_X1    g132(.A(new_n533), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n525), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n555), .A2(new_n557), .A3(new_n559), .A4(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  OAI21_X1  g141(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n567));
  INV_X1    g142(.A(G87), .ZN(new_n568));
  INV_X1    g143(.A(G49), .ZN(new_n569));
  OAI221_X1 g144(.A(new_n567), .B1(new_n533), .B2(new_n568), .C1(new_n569), .C2(new_n520), .ZN(G288));
  NAND3_X1  g145(.A1(new_n510), .A2(G48), .A3(G543), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n533), .ZN(new_n573));
  OAI21_X1  g148(.A(G61), .B1(new_n523), .B2(new_n524), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n515), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(KEYINPUT74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(KEYINPUT74), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n558), .A2(G85), .B1(new_n550), .B2(G47), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n515), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n509), .A2(new_n510), .A3(G92), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n525), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n550), .B2(G54), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n584), .B1(new_n591), .B2(G868), .ZN(G321));
  XOR2_X1   g167(.A(G321), .B(KEYINPUT75), .Z(G284));
  NAND2_X1  g168(.A1(G286), .A2(G868), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n551), .A2(new_n554), .A3(KEYINPUT9), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n557), .A2(new_n563), .A3(new_n559), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n594), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n594), .B1(new_n597), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G860), .ZN(G148));
  INV_X1    g176(.A(new_n542), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n591), .A2(KEYINPUT76), .A3(new_n600), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n586), .A2(new_n590), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G559), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  MUX2_X1   g182(.A(new_n602), .B(new_n607), .S(G868), .Z(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n463), .A2(new_n482), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2100), .ZN(new_n613));
  INV_X1    g188(.A(new_n492), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G123), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT77), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G111), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G2105), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n481), .B2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(G2096), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(G2096), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n613), .A2(new_n622), .A3(new_n623), .ZN(G156));
  INV_X1    g199(.A(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n627), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n630), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT78), .Z(G401));
  INV_X1    g215(.A(KEYINPUT18), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n644), .B2(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT79), .ZN(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n661), .A2(new_n654), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(new_n661), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT80), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n665), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n671), .B1(new_n670), .B2(new_n672), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n675), .ZN(new_n678));
  INV_X1    g253(.A(new_n671), .ZN(new_n679));
  INV_X1    g254(.A(new_n672), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n669), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n678), .B1(new_n681), .B2(new_n673), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n682), .ZN(G229));
  NAND2_X1  g258(.A1(G303), .A2(G16), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G22), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(KEYINPUT83), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(KEYINPUT83), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(G1971), .A3(new_n689), .ZN(new_n693));
  NOR2_X1   g268(.A1(G6), .A2(G16), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n579), .B2(G16), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n692), .A2(new_n693), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n685), .A2(G23), .ZN(new_n701));
  INV_X1    g276(.A(G288), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n685), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n704), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n701), .B(new_n706), .C1(new_n702), .C2(new_n685), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n705), .A2(new_n707), .B1(new_n695), .B2(new_n697), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT84), .B1(new_n700), .B2(new_n709), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n690), .A2(new_n691), .B1(new_n696), .B2(new_n698), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n711), .A2(new_n712), .A3(new_n708), .A4(new_n693), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n710), .A2(new_n713), .A3(KEYINPUT34), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n481), .A2(G131), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT81), .ZN(new_n719));
  OR2_X1    g294(.A1(G95), .A2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n720), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT82), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G119), .B2(new_n614), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G25), .B2(G29), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  AND2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  MUX2_X1   g305(.A(G24), .B(G290), .S(G16), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n716), .A2(new_n717), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(KEYINPUT36), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n716), .A2(new_n736), .A3(new_n717), .A4(new_n733), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n463), .A2(G127), .ZN(new_n739));
  NAND2_X1  g314(.A1(G115), .A2(G2104), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n465), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G139), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n480), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT88), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n747));
  NAND3_X1  g322(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n745), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n746), .B1(new_n745), .B2(new_n749), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n742), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G33), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT90), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(KEYINPUT90), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G2072), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n754), .A2(G35), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n493), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n754), .A2(G26), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT28), .ZN(new_n766));
  INV_X1    g341(.A(G140), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n480), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT86), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  INV_X1    g346(.A(G116), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n614), .B2(G128), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n766), .B1(new_n776), .B2(new_n754), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g354(.A(G2067), .B(new_n766), .C1(new_n776), .C2(new_n754), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n763), .A2(new_n764), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G164), .A2(new_n754), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G27), .B2(new_n754), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT93), .B(G2078), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT24), .A2(G34), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT24), .ZN(new_n787));
  INV_X1    g362(.A(G34), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n484), .A2(G29), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n783), .A2(new_n784), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n785), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n795), .A2(G28), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n754), .B1(new_n795), .B2(G28), .ZN(new_n797));
  AND2_X1   g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  NOR2_X1   g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  OAI22_X1  g374(.A1(new_n796), .A2(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n685), .A2(G5), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G301), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1961), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n685), .A2(G19), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT85), .Z(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n542), .B2(new_n685), .ZN(new_n807));
  INV_X1    g382(.A(G1341), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n685), .A2(G21), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G168), .B2(new_n685), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(G1966), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(G1966), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n814), .B(new_n815), .C1(new_n803), .C2(new_n802), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n685), .A2(G20), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT23), .Z(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G299), .B2(G16), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT95), .B(G1956), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n820), .B(new_n821), .Z(new_n822));
  NAND4_X1  g397(.A1(new_n781), .A2(new_n794), .A3(new_n817), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n685), .A2(G4), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n591), .B2(new_n685), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(G1348), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(G1348), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n621), .A2(new_n754), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n790), .A2(new_n791), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT91), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(KEYINPUT91), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n754), .A2(G32), .ZN(new_n833));
  NAND3_X1  g408(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT26), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n836), .A2(new_n837), .B1(G105), .B2(new_n482), .ZN(new_n838));
  INV_X1    g413(.A(G129), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n492), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n481), .A2(G141), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n833), .B1(new_n842), .B2(new_n754), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT27), .B(G1996), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT92), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n843), .B(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n829), .A2(new_n831), .A3(new_n832), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n823), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n763), .A2(new_n764), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT94), .Z(new_n850));
  INV_X1    g425(.A(G2072), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n757), .A2(new_n851), .A3(new_n758), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n760), .A2(new_n848), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT96), .B1(new_n738), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n856));
  AOI211_X1 g431(.A(new_n856), .B(new_n853), .C1(new_n735), .C2(new_n737), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(G311));
  NAND2_X1  g433(.A1(new_n738), .A2(new_n854), .ZN(G150));
  NAND2_X1  g434(.A1(new_n591), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n515), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT97), .B(G55), .Z(new_n864));
  XOR2_X1   g439(.A(KEYINPUT98), .B(G93), .Z(new_n865));
  OAI22_X1  g440(.A1(new_n520), .A2(new_n864), .B1(new_n533), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n542), .A2(new_n867), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n541), .A2(new_n538), .B1(new_n863), .B2(new_n866), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n861), .B(new_n870), .Z(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n872));
  INV_X1    g447(.A(G860), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n867), .A2(new_n873), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(G145));
  XNOR2_X1  g453(.A(new_n621), .B(new_n493), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n484), .B(KEYINPUT99), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n842), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n752), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n742), .B(new_n842), .C1(new_n750), .C2(new_n751), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n724), .B(new_n611), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n775), .B(G164), .ZN(new_n888));
  OR2_X1    g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n890));
  INV_X1    g465(.A(G130), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n890), .B1(new_n492), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n481), .B2(G142), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n888), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n886), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n883), .A3(new_n884), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n887), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n894), .B1(new_n887), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n881), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n887), .A2(new_n896), .ZN(new_n900));
  INV_X1    g475(.A(new_n894), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n881), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n887), .A2(new_n894), .A3(new_n896), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n899), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g483(.A(KEYINPUT102), .B1(new_n867), .B2(G868), .ZN(new_n909));
  INV_X1    g484(.A(G868), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n607), .B(new_n870), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n591), .A2(new_n597), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n605), .A2(G299), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n912), .A2(KEYINPUT41), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT41), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n912), .A2(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(G288), .B(KEYINPUT100), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(G305), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G290), .B(G303), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n921), .A2(G305), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n924), .B1(new_n928), .B2(new_n922), .ZN(new_n929));
  OAI22_X1  g504(.A1(new_n927), .A2(new_n929), .B1(KEYINPUT101), .B2(KEYINPUT42), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n920), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n917), .A2(new_n930), .A3(new_n919), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n910), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n932), .A2(KEYINPUT101), .A3(KEYINPUT42), .A4(new_n933), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n909), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n917), .A2(new_n930), .A3(new_n919), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n930), .B1(new_n917), .B2(new_n919), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n935), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND4_X1   g517(.A1(new_n939), .A2(new_n937), .A3(G868), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n938), .A2(new_n943), .ZN(G295));
  NOR2_X1   g519(.A1(new_n938), .A2(new_n943), .ZN(G331));
  OR2_X1    g520(.A1(new_n927), .A2(new_n929), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n531), .B2(new_n535), .ZN(new_n948));
  NAND2_X1  g523(.A1(G171), .A2(KEYINPUT103), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n870), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n948), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n869), .A3(new_n868), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n952), .A3(G168), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G168), .B1(new_n950), .B2(new_n952), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n916), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n955), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n957), .A2(new_n913), .A3(new_n912), .A4(new_n953), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n946), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n927), .A2(new_n929), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  INV_X1    g536(.A(new_n913), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n605), .A2(G299), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT41), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n953), .B2(new_n957), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n954), .A2(new_n955), .A3(new_n918), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n960), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n959), .A2(new_n969), .A3(new_n906), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n956), .A2(new_n958), .ZN(new_n973));
  AOI21_X1  g548(.A(G37), .B1(new_n973), .B2(new_n960), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n974), .B2(new_n959), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT44), .ZN(G397));
  INV_X1    g552(.A(KEYINPUT57), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n978), .B1(new_n597), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(G299), .A2(KEYINPUT114), .A3(KEYINPUT57), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n499), .B2(new_n504), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n482), .A2(G101), .ZN(new_n986));
  INV_X1    g561(.A(G137), .ZN(new_n987));
  OAI211_X1 g562(.A(G40), .B(new_n986), .C1(new_n480), .C2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n466), .B2(new_n475), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT45), .B(new_n982), .C1(new_n499), .C2(new_n504), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT56), .B(G2072), .Z(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n985), .A2(new_n989), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n980), .A2(new_n981), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n983), .A2(KEYINPUT50), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n996), .B(new_n982), .C1(new_n499), .C2(new_n504), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n989), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1956), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(KEYINPUT113), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT113), .B1(new_n998), .B2(new_n999), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n994), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n993), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1002), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(new_n1000), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n980), .A2(new_n981), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1348), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n998), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n504), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n463), .A2(new_n498), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(new_n989), .A3(new_n778), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1016), .A2(new_n989), .A3(KEYINPUT115), .A4(new_n778), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1011), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(new_n605), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1003), .B1(new_n1009), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT60), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n605), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI211_X1 g605(.A(KEYINPUT118), .B(new_n605), .C1(new_n1021), .C2(new_n1025), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT60), .B1(new_n1033), .B2(new_n1011), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT118), .B1(new_n1034), .B2(new_n605), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1026), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1003), .B(KEYINPUT61), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1016), .A2(new_n989), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT58), .B(G1341), .Z(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1996), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n985), .A2(new_n1044), .A3(new_n989), .A4(new_n990), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n542), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1040), .B1(new_n1047), .B2(KEYINPUT59), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(KEYINPUT116), .A3(KEYINPUT59), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n602), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1048), .A2(new_n1049), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n993), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1005), .A2(new_n1000), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1056), .A2(new_n1007), .B1(new_n1057), .B2(new_n994), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1039), .B(new_n1055), .C1(new_n1058), .C2(KEYINPUT61), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1024), .B1(new_n1038), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n998), .A2(new_n803), .ZN(new_n1062));
  INV_X1    g637(.A(G2078), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n985), .A2(new_n1063), .A3(new_n989), .A4(new_n990), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT119), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n1064), .B2(KEYINPUT119), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT120), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1070), .B(new_n1062), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1064), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G301), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(G301), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1063), .A2(KEYINPUT53), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n1078), .B(new_n988), .C1(G2105), .C2(new_n473), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(new_n985), .A3(new_n990), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1077), .A2(new_n1062), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1061), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n985), .A2(new_n989), .A3(new_n990), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n691), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n995), .A2(new_n764), .A3(new_n989), .A4(new_n997), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G8), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT107), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n511), .A2(new_n512), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n508), .B1(new_n533), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(G62), .B1(new_n523), .B2(new_n524), .ZN(new_n1091));
  NAND2_X1  g666(.A1(G75), .A2(G543), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n515), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT55), .B(G8), .C1(new_n1090), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT105), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT105), .ZN(new_n1096));
  NAND4_X1  g671(.A1(G303), .A2(new_n1096), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT106), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(new_n1097), .A3(KEYINPUT106), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n1088), .A2(new_n1100), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1088), .B1(new_n1105), .B2(new_n1101), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1087), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT107), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1105), .A2(new_n1088), .A3(new_n1101), .ZN(new_n1110));
  INV_X1    g685(.A(G8), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT49), .ZN(new_n1114));
  AOI211_X1 g689(.A(G1981), .B(new_n573), .C1(new_n577), .C2(new_n578), .ZN(new_n1115));
  INV_X1    g690(.A(G1981), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT108), .B(G86), .Z(new_n1117));
  OAI21_X1  g692(.A(new_n571), .B1(new_n533), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n576), .B1(new_n1118), .B2(KEYINPUT109), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT109), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n571), .B(new_n1120), .C1(new_n533), .C2(new_n1117), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1116), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1114), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n573), .ZN(new_n1124));
  INV_X1    g699(.A(new_n578), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n576), .A2(KEYINPUT74), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1116), .B(new_n1124), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1118), .A2(KEYINPUT109), .ZN(new_n1128));
  INV_X1    g703(.A(new_n576), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1121), .ZN(new_n1130));
  OAI211_X1 g705(.A(KEYINPUT49), .B(new_n1127), .C1(new_n1130), .C2(new_n1116), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1111), .B1(new_n1016), .B2(new_n989), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1123), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n702), .A2(G1976), .ZN(new_n1134));
  INV_X1    g709(.A(G1976), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT52), .B1(G288), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT52), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1133), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1107), .A2(new_n1113), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1966), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1083), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n995), .A2(new_n791), .A3(new_n989), .A4(new_n997), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(G168), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(G8), .ZN(new_n1146));
  AOI21_X1  g721(.A(G168), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT51), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT51), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1145), .A2(new_n1150), .A3(G8), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1141), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1074), .A2(new_n1062), .A3(new_n1080), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT54), .B1(new_n1154), .B2(G301), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1060), .A2(new_n1082), .A3(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1064), .A2(KEYINPUT119), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(KEYINPUT53), .A3(new_n1065), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1070), .B1(new_n1160), .B2(new_n1062), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1071), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1074), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1148), .A2(new_n1164), .A3(new_n1151), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1163), .A2(new_n1141), .A3(new_n1165), .A4(G171), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1075), .A2(KEYINPUT121), .A3(new_n1141), .A4(new_n1165), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT62), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1127), .B(KEYINPUT110), .Z(new_n1172));
  NOR2_X1   g747(.A1(G288), .A2(G1976), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n1133), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT111), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1132), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1140), .ZN(new_n1178));
  OAI22_X1  g753(.A1(new_n1176), .A2(new_n1177), .B1(new_n1113), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g754(.A(new_n1111), .B(G286), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1107), .A2(new_n1113), .A3(new_n1140), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT63), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1182), .A2(KEYINPUT112), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1181), .B(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(KEYINPUT112), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1179), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1158), .A2(new_n1171), .A3(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n989), .A2(new_n984), .A3(new_n983), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1044), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT104), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n775), .B(new_n778), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(new_n1044), .B2(new_n842), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1191), .A2(new_n842), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n725), .A2(new_n728), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n725), .A2(new_n728), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1188), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(G290), .B(G1986), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1199), .B1(new_n1188), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1187), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT46), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1190), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT124), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT47), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1192), .A2(new_n842), .ZN(new_n1207));
  AOI22_X1  g782(.A1(new_n1191), .A2(KEYINPUT46), .B1(new_n1188), .B2(new_n1207), .ZN(new_n1208));
  AND3_X1   g783(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1206), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1210));
  NOR2_X1   g785(.A1(G290), .A2(G1986), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1188), .A2(new_n1211), .ZN(new_n1212));
  XOR2_X1   g787(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1213));
  XNOR2_X1  g788(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1214), .B1(new_n1199), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g791(.A(KEYINPUT125), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1217));
  OAI22_X1  g792(.A1(new_n1209), .A2(new_n1210), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT123), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1194), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1195), .B(KEYINPUT122), .Z(new_n1221));
  NOR2_X1   g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n775), .A2(G2067), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1219), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  OAI221_X1 g799(.A(KEYINPUT123), .B1(G2067), .B2(new_n775), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1225));
  AND2_X1   g800(.A1(new_n1225), .A2(new_n1188), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1218), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1202), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g803(.A1(new_n639), .A2(new_n459), .A3(G227), .ZN(new_n1230));
  AND3_X1   g804(.A1(new_n677), .A2(new_n682), .A3(new_n1230), .ZN(new_n1231));
  OAI211_X1 g805(.A(new_n907), .B(new_n1231), .C1(new_n971), .C2(new_n975), .ZN(G225));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n1233));
  NOR2_X1   g807(.A1(G225), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g808(.A1(new_n677), .A2(new_n682), .A3(new_n1230), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n1236));
  NAND3_X1  g810(.A1(new_n974), .A2(new_n972), .A3(new_n959), .ZN(new_n1237));
  AOI21_X1  g811(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g812(.A(KEYINPUT127), .B1(new_n1238), .B2(new_n907), .ZN(new_n1239));
  NOR2_X1   g813(.A1(new_n1234), .A2(new_n1239), .ZN(G308));
endmodule


