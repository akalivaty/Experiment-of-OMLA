//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n615, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n466), .B2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n474), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n475), .A2(new_n469), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g056(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n468), .A2(G2105), .A3(new_n470), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(G136), .B2(new_n472), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n470), .A2(new_n465), .A3(new_n467), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n469), .C1(new_n491), .C2(KEYINPUT69), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(KEYINPUT4), .A2(new_n490), .B1(new_n495), .B2(new_n474), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n470), .A2(new_n465), .A3(new_n467), .A4(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT70), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(new_n494), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n474), .A2(new_n504), .A3(new_n489), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(new_n501), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n502), .A2(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT71), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n514), .A2(new_n515), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n517), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(G62), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  XOR2_X1   g106(.A(new_n531), .B(KEYINPUT72), .Z(new_n532));
  AOI21_X1  g107(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n528), .A2(new_n533), .ZN(G166));
  NAND2_X1  g109(.A1(new_n522), .A2(new_n523), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n514), .B2(new_n515), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(G51), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n537), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  AOI22_X1  g118(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n529), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n516), .A2(G52), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n526), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n529), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n516), .A2(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n526), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  AND3_X1   g135(.A1(new_n522), .A2(G65), .A3(new_n523), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT75), .Z(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n524), .A2(G91), .A3(new_n525), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n515), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n567), .C2(new_n513), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT74), .B1(new_n569), .B2(KEYINPUT73), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(KEYINPUT74), .B2(new_n569), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n566), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  OR2_X1    g151(.A1(G171), .A2(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g152(.A1(G171), .A2(KEYINPUT76), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(G301));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g155(.A1(G166), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n528), .B2(new_n533), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G303));
  AOI22_X1  g158(.A1(new_n536), .A2(G87), .B1(G49), .B2(new_n516), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G288));
  AOI22_X1  g161(.A1(new_n536), .A2(G86), .B1(G48), .B2(new_n516), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n522), .A2(G61), .A3(new_n523), .ZN(new_n588));
  AND2_X1   g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n536), .A2(G85), .B1(G47), .B2(new_n516), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n529), .B2(new_n593), .ZN(G290));
  NAND3_X1  g169(.A1(new_n524), .A2(G92), .A3(new_n525), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n535), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G54), .B2(new_n516), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n597), .A2(new_n601), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT78), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  MUX2_X1   g183(.A(G301), .B(new_n607), .S(new_n608), .Z(G321));
  XOR2_X1   g184(.A(G321), .B(KEYINPUT79), .Z(G284));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n575), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(G868), .B2(new_n575), .ZN(G280));
  INV_X1    g188(.A(new_n607), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  OAI21_X1  g191(.A(G868), .B1(new_n607), .B2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n472), .A2(G135), .ZN(new_n620));
  INV_X1    g195(.A(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n469), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n620), .B1(new_n621), .B2(new_n484), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT80), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n474), .A2(new_n477), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n627), .A2(new_n628), .A3(new_n632), .ZN(G156));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n639), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT81), .Z(new_n651));
  NOR2_X1   g226(.A1(G2072), .A2(G2078), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n442), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(KEYINPUT17), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n649), .B(new_n650), .C1(new_n442), .C2(new_n652), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n655), .A3(new_n649), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2096), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT82), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n667), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT83), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n677), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT84), .B(G1986), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  MUX2_X1   g261(.A(G23), .B(G288), .S(G16), .Z(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT33), .B(G1976), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  NOR2_X1   g264(.A1(G6), .A2(G16), .ZN(new_n690));
  INV_X1    g265(.A(G305), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G16), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1971), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n689), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT34), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G1986), .Z(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G25), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n472), .A2(G131), .ZN(new_n707));
  INV_X1    g282(.A(G119), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n469), .A2(G107), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n710));
  OAI22_X1  g285(.A1(new_n484), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n705), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n701), .A2(new_n702), .A3(new_n704), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT36), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT24), .B(G34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(new_n705), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT90), .Z(new_n720));
  INV_X1    g295(.A(G160), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n705), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT91), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G2084), .ZN(new_n724));
  NOR2_X1   g299(.A1(G29), .A2(G33), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT87), .Z(new_n726));
  NAND3_X1  g301(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT25), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(new_n469), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n728), .B1(new_n730), .B2(KEYINPUT89), .ZN(new_n731));
  INV_X1    g306(.A(G139), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n471), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(KEYINPUT88), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(KEYINPUT88), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n731), .B1(KEYINPUT89), .B2(new_n730), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n726), .B1(new_n736), .B2(new_n705), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2072), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n705), .A2(G32), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT26), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n742), .A2(new_n743), .B1(G105), .B2(new_n477), .ZN(new_n744));
  INV_X1    g319(.A(G129), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n484), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G141), .B2(new_n472), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n705), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT27), .B(G1996), .Z(new_n749));
  OAI211_X1 g324(.A(new_n724), .B(new_n738), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT92), .Z(new_n751));
  NOR2_X1   g326(.A1(G171), .A2(new_n695), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G5), .B2(new_n695), .ZN(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT85), .B(G1341), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT86), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n555), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G16), .B2(G19), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n755), .B(new_n756), .C1(new_n758), .C2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n762), .A2(G28), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n705), .B1(new_n762), .B2(G28), .ZN(new_n764));
  AND2_X1   g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  NOR2_X1   g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  OAI22_X1  g341(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G168), .A2(new_n695), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n695), .B2(G21), .ZN(new_n769));
  INV_X1    g344(.A(G1966), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n625), .A2(G29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n748), .A2(new_n749), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n760), .A2(new_n758), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n695), .A2(G20), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT23), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n575), .B2(new_n695), .ZN(new_n778));
  INV_X1    g353(.A(G1956), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G29), .A2(G35), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G162), .B2(G29), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G2090), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n761), .A2(new_n775), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n695), .A2(G4), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n614), .B2(new_n695), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n769), .A2(new_n770), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT93), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n784), .A2(new_n785), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(KEYINPUT95), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n705), .A2(G26), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT28), .ZN(new_n798));
  INV_X1    g373(.A(G128), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n469), .A2(G116), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n484), .A2(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G140), .B2(new_n472), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n798), .B1(new_n803), .B2(new_n705), .ZN(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n723), .A2(G2084), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n794), .A2(new_n796), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G27), .A2(G29), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G164), .B2(G29), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n795), .B2(KEYINPUT95), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n751), .A2(new_n792), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n717), .A2(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  NOR2_X1   g391(.A1(new_n607), .A2(new_n615), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n529), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n516), .A2(G55), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n526), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n555), .B(new_n825), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n819), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n828));
  AOI21_X1  g403(.A(G860), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  OAI21_X1  g405(.A(G860), .B1(new_n821), .B2(new_n824), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(G145));
  XNOR2_X1  g408(.A(new_n736), .B(new_n747), .ZN(new_n834));
  OR2_X1    g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n836));
  INV_X1    g411(.A(G130), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n484), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G142), .B2(new_n472), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n630), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n834), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n498), .A2(new_n842), .A3(new_n500), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n498), .B2(new_n500), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n507), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n803), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n712), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n841), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n625), .B(G160), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(G162), .Z(new_n850));
  OR2_X1    g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(G37), .B1(new_n848), .B2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n826), .B1(new_n607), .B2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n555), .B(new_n825), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n857), .A2(new_n615), .A3(new_n606), .A4(new_n604), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n602), .A2(G299), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n605), .A2(new_n575), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n860), .A2(KEYINPUT41), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n859), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n860), .A2(KEYINPUT98), .A3(new_n861), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n858), .A3(new_n856), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n867), .A2(new_n871), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n871), .B1(new_n867), .B2(new_n876), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n691), .B(G290), .ZN(new_n879));
  XNOR2_X1  g454(.A(G166), .B(G288), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(KEYINPUT99), .B2(KEYINPUT42), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n877), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n867), .A2(new_n876), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n870), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n867), .A2(new_n871), .A3(new_n876), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(G868), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n825), .A2(G868), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n855), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n882), .B1(new_n877), .B2(new_n878), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n886), .A2(new_n884), .A3(new_n887), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n608), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n895), .A2(KEYINPUT100), .A3(new_n890), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n892), .A2(new_n896), .ZN(G295));
  NAND2_X1  g472(.A1(new_n889), .A2(new_n891), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n900));
  NOR2_X1   g475(.A1(G168), .A2(G171), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n857), .B(new_n902), .C1(G301), .C2(G286), .ZN(new_n903));
  AOI21_X1  g478(.A(G286), .B1(new_n577), .B2(new_n578), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n826), .B1(new_n904), .B2(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n862), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n866), .A2(new_n905), .A3(new_n903), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n881), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n903), .A2(new_n905), .B1(new_n873), .B2(new_n874), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n881), .B1(new_n913), .B2(new_n908), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n900), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n881), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n866), .A2(new_n905), .A3(new_n903), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n912), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n918), .A2(KEYINPUT103), .A3(new_n909), .A4(new_n910), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n899), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n907), .A2(new_n908), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT101), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n907), .A2(new_n923), .A3(new_n908), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n916), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n911), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT43), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n920), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n918), .A2(new_n899), .A3(new_n909), .A4(new_n910), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n929), .A2(KEYINPUT102), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n899), .B1(new_n925), .B2(new_n926), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(KEYINPUT102), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n930), .B(new_n931), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n934), .ZN(G397));
  NAND2_X1  g510(.A1(new_n501), .A2(KEYINPUT97), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n498), .A2(new_n842), .A3(new_n500), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G1384), .B1(new_n938), .B2(new_n507), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n473), .A2(G40), .A3(new_n476), .A4(new_n478), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT45), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n712), .ZN(new_n943));
  INV_X1    g518(.A(new_n714), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n803), .B(new_n805), .ZN(new_n946));
  INV_X1    g521(.A(G1996), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n747), .B(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n949), .B2(new_n942), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n803), .A2(new_n805), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n942), .B1(new_n952), .B2(KEYINPUT126), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(KEYINPUT126), .B2(new_n952), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT127), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n941), .A2(new_n947), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT46), .ZN(new_n959));
  INV_X1    g534(.A(new_n747), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n941), .B1(new_n946), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  INV_X1    g538(.A(new_n945), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n943), .A2(new_n944), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n949), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n968));
  OR3_X1    g543(.A1(new_n942), .A2(G1986), .A3(G290), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n967), .A2(new_n942), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  NOR4_X1   g546(.A1(new_n956), .A2(new_n957), .A3(new_n963), .A4(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G8), .ZN(new_n973));
  INV_X1    g548(.A(new_n940), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n939), .ZN(new_n975));
  INV_X1    g550(.A(G1981), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n590), .B2(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g552(.A1(G305), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n587), .B(new_n590), .C1(KEYINPUT107), .C2(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(KEYINPUT49), .A3(new_n979), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n975), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(G288), .A2(G1976), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(G305), .A2(G1981), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n975), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n581), .A2(G8), .A3(new_n582), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT106), .B(KEYINPUT55), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n581), .A2(G8), .A3(new_n582), .A4(new_n990), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(G1384), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n845), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT104), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT104), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n845), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n502), .A2(new_n510), .A3(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n998), .A2(new_n1000), .B1(new_n995), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1971), .B1(new_n1003), .B2(new_n974), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n940), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT105), .B1(new_n939), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n845), .A2(KEYINPUT105), .A3(new_n1006), .A4(new_n1001), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1005), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G2090), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n994), .B(G8), .C1(new_n1004), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n975), .B1(new_n1013), .B2(G288), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n975), .B(new_n1016), .C1(new_n1013), .C2(G288), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n984), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n988), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT63), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1018), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n502), .A2(new_n510), .A3(new_n1006), .A4(new_n1001), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n974), .B(new_n1022), .C1(new_n1006), .C2(new_n939), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(G2090), .ZN(new_n1024));
  OAI21_X1  g599(.A(G8), .B1(new_n1004), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n994), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1021), .A2(new_n1027), .A3(new_n1012), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n845), .A2(new_n1001), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n940), .B1(new_n1029), .B2(new_n995), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n502), .A2(new_n510), .A3(new_n996), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT108), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n502), .A2(new_n510), .A3(KEYINPUT108), .A4(new_n996), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n770), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n845), .A2(new_n1006), .A3(new_n1001), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT105), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1008), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n1005), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(G8), .A3(G168), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1020), .B1(new_n1028), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1020), .ZN(new_n1046));
  OAI21_X1  g621(.A(G8), .B1(new_n1011), .B2(new_n1004), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1026), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1046), .A2(new_n1012), .A3(new_n1021), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1019), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(KEYINPUT122), .A2(G8), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n1043), .B2(G286), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT51), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(new_n1051), .C1(new_n1043), .C2(G286), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1043), .A2(G8), .A3(G286), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT62), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1053), .A2(new_n1059), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n998), .A2(new_n1000), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1002), .A2(new_n995), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1061), .A2(new_n811), .A3(new_n1062), .A4(new_n974), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1010), .A2(new_n754), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(G2078), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1030), .A2(new_n1033), .A3(new_n1067), .A4(new_n1034), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G301), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1028), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1058), .A2(new_n1060), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1050), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n574), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n572), .B(KEYINPUT110), .C1(new_n568), .C2(new_n573), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1076), .A2(new_n564), .A3(new_n565), .A4(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT109), .B(KEYINPUT57), .Z(new_n1079));
  AND3_X1   g654(.A1(new_n1078), .A2(KEYINPUT111), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT111), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1080), .A2(new_n1081), .B1(new_n1082), .B2(G299), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT112), .B(KEYINPUT56), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(G2072), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1061), .A2(new_n1062), .A3(new_n974), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1023), .A2(new_n779), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI221_X1 g665(.A(KEYINPUT113), .B1(G299), .B2(new_n1082), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1083), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1348), .B1(new_n1040), .B2(new_n1005), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n974), .A2(new_n939), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(G2067), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n605), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1093), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1010), .A2(new_n790), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1097), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n602), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1103), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n605), .A2(KEYINPUT121), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1098), .A2(KEYINPUT121), .A3(KEYINPUT60), .A4(new_n605), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1092), .A2(KEYINPUT61), .A3(new_n1094), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(KEYINPUT120), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1083), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1090), .A2(new_n1115), .A3(KEYINPUT119), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1094), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1083), .B1(new_n1089), .B2(new_n1088), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1114), .B(new_n1116), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1092), .A2(new_n1121), .A3(KEYINPUT61), .A4(new_n1094), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n1124));
  INV_X1    g699(.A(new_n555), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT114), .B(G1996), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n940), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1000), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n999), .B1(new_n845), .B2(new_n996), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1062), .B(new_n1127), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT58), .B(G1341), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n1096), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1125), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT59), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT115), .B(new_n1125), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1138), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1003), .A2(new_n1127), .B1(new_n1096), .B2(new_n1131), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT115), .B1(new_n1143), .B2(new_n1125), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(KEYINPUT116), .A4(KEYINPUT59), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1137), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1113), .B(new_n1123), .C1(new_n1124), .C2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1147), .A2(new_n1124), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1100), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1028), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1061), .A2(new_n1030), .A3(new_n1067), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1065), .A2(G301), .A3(new_n1066), .A4(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1071), .A2(KEYINPUT123), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1153), .B2(KEYINPUT123), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1151), .B(new_n1057), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1065), .A2(new_n1066), .A3(new_n1152), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(G171), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1159), .A2(KEYINPUT124), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(KEYINPUT124), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(new_n1155), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT125), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1160), .A2(new_n1163), .A3(new_n1166), .A4(new_n1161), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1157), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1074), .B1(new_n1150), .B2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(G290), .B(G1986), .Z(new_n1170));
  AOI21_X1  g745(.A(new_n942), .B1(new_n967), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n972), .B1(new_n1169), .B2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g747(.A1(G401), .A2(new_n461), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n685), .A2(new_n663), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g749(.A(new_n1175), .B1(new_n851), .B2(new_n852), .ZN(new_n1176));
  OAI211_X1 g750(.A(new_n1176), .B(new_n930), .C1(new_n932), .C2(new_n933), .ZN(G225));
  INV_X1    g751(.A(G225), .ZN(G308));
endmodule


