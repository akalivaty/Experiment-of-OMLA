//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT27), .B(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT28), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n211), .B1(KEYINPUT26), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(KEYINPUT26), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n215), .A2(new_n216), .B1(G183gat), .B2(G190gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(KEYINPUT23), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G183gat), .B(G190gat), .Z(new_n222));
  AOI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(KEYINPUT24), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT64), .B(G169gat), .Z(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(G176gat), .ZN(new_n226));
  AOI211_X1 g025(.A(KEYINPUT25), .B(new_n211), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n209), .A2(new_n217), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n210), .B1(new_n214), .B2(new_n225), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  INV_X1    g029(.A(new_n223), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT25), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G113gat), .ZN(new_n237));
  INV_X1    g036(.A(G120gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT1), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G113gat), .A2(G120gat), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n234), .A2(new_n235), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n236), .B(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n233), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(new_n242), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(G227gat), .A3(G233gat), .A4(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT33), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n204), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(KEYINPUT32), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT67), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n244), .ZN(new_n251));
  INV_X1    g050(.A(G227gat), .ZN(new_n252));
  INV_X1    g051(.A(G233gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT34), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n254), .B(KEYINPUT34), .Z(new_n257));
  NAND3_X1  g056(.A1(new_n249), .A2(new_n257), .A3(KEYINPUT67), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(KEYINPUT36), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT36), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n249), .A2(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n247), .A2(new_n248), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n247), .A2(new_n248), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n255), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n260), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G211gat), .A2(G218gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(KEYINPUT22), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(G211gat), .A2(G218gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n272), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G155gat), .ZN(new_n276));
  INV_X1    g075(.A(G162gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT2), .ZN(new_n279));
  NOR2_X1   g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(KEYINPUT70), .B(G148gat), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G141gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT69), .B(G141gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G148gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(KEYINPUT2), .ZN(new_n288));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289));
  AOI211_X1 g088(.A(new_n280), .B(new_n278), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n275), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n270), .A2(KEYINPUT75), .A3(new_n272), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n294), .B(new_n296), .C1(new_n275), .C2(KEYINPUT75), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n292), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n286), .A2(new_n290), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(G228gat), .A2(G233gat), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT3), .B1(new_n275), .B2(new_n294), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(new_n291), .ZN(new_n303));
  OAI22_X1  g102(.A1(new_n300), .A2(new_n301), .B1(new_n295), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT31), .B(G50gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G22gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(KEYINPUT76), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n308), .B2(new_n307), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n304), .B(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n242), .B1(new_n299), .B2(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n293), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT5), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n242), .A2(new_n291), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT4), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n242), .A2(new_n291), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G1gat), .B(G29gat), .Z(new_n325));
  XNOR2_X1  g124(.A(G57gat), .B(G85gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT72), .B(KEYINPUT0), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(KEYINPUT4), .B2(new_n319), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n322), .A2(new_n330), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n316), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n242), .B(new_n291), .ZN(new_n335));
  INV_X1    g134(.A(new_n315), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT5), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n324), .B(new_n329), .C1(new_n334), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n331), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n333), .A3(new_n320), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n317), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT5), .A3(new_n337), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(KEYINPUT73), .A3(new_n329), .A4(new_n324), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT6), .ZN(new_n347));
  INV_X1    g146(.A(new_n329), .ZN(new_n348));
  INV_X1    g147(.A(new_n324), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n338), .B1(new_n343), .B2(new_n317), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n341), .A2(new_n346), .A3(new_n347), .A4(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n351), .A2(new_n347), .ZN(new_n353));
  INV_X1    g152(.A(G226gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(new_n253), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n355), .B1(new_n233), .B2(new_n294), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n233), .A2(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n275), .ZN(new_n361));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(KEYINPUT68), .ZN(new_n365));
  INV_X1    g164(.A(new_n358), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(new_n356), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(KEYINPUT68), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n361), .B(new_n364), .C1(new_n369), .C2(new_n275), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n352), .A2(new_n353), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT38), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT37), .ZN(new_n373));
  INV_X1    g172(.A(new_n275), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n373), .B1(new_n360), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n369), .A2(new_n374), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n364), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n275), .B1(new_n367), .B2(new_n368), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n359), .A2(new_n374), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n373), .B2(new_n364), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n379), .A2(KEYINPUT79), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n361), .B1(new_n369), .B2(new_n275), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n386), .A2(KEYINPUT37), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n380), .B1(new_n386), .B2(KEYINPUT37), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT38), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n388), .B2(new_n378), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n385), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n315), .B1(new_n323), .B2(new_n314), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT39), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n348), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT39), .B1(new_n335), .B2(new_n336), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT40), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n351), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n397), .A2(new_n398), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n401), .A2(KEYINPUT78), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(KEYINPUT78), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OR4_X1    g203(.A1(KEYINPUT30), .A2(new_n381), .A3(new_n382), .A4(new_n380), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n370), .A2(new_n383), .A3(KEYINPUT30), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT77), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT77), .B1(new_n405), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n312), .B1(new_n392), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n352), .A2(new_n353), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n405), .A2(new_n406), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT74), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n414), .A2(new_n415), .A3(new_n311), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n266), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n249), .A2(new_n257), .A3(KEYINPUT67), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n257), .B1(new_n249), .B2(KEYINPUT67), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n311), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n414), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT35), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n407), .A2(new_n408), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n261), .A2(new_n264), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n426), .A2(new_n422), .A3(new_n411), .A4(new_n311), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n421), .A2(new_n422), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n417), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n308), .A2(G15gat), .ZN(new_n430));
  INV_X1    g229(.A(G15gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G22gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G1gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT16), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n430), .B(new_n432), .C1(new_n436), .C2(G1gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(KEYINPUT85), .A3(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(G8gat), .C1(KEYINPUT85), .C2(new_n437), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n437), .A2(KEYINPUT86), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(KEYINPUT86), .ZN(new_n441));
  INV_X1    g240(.A(G8gat), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .A4(new_n435), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(G43gat), .A2(G50gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(G43gat), .A2(G50gat), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT15), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT14), .ZN(new_n448));
  INV_X1    g247(.A(G29gat), .ZN(new_n449));
  INV_X1    g248(.A(G36gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n453), .A2(KEYINPUT81), .B1(G29gat), .B2(G36gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n452), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT81), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n447), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G43gat), .ZN(new_n459));
  INV_X1    g258(.A(G50gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G43gat), .A2(G50gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n463), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n451), .A2(KEYINPUT83), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n466), .A2(new_n448), .A3(new_n449), .A4(new_n450), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n467), .A3(new_n452), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n445), .A2(new_n446), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT82), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n461), .A2(KEYINPUT82), .A3(new_n470), .A4(new_n462), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n464), .B(new_n468), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n470), .A3(new_n462), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n472), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n480), .A2(KEYINPUT84), .A3(new_n468), .A4(new_n464), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n458), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n444), .B1(new_n482), .B2(KEYINPUT17), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n454), .A2(new_n457), .ZN(new_n484));
  INV_X1    g283(.A(new_n447), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G29gat), .A2(G36gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n447), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n479), .B2(new_n472), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT84), .B1(new_n489), .B2(new_n468), .ZN(new_n490));
  AND4_X1   g289(.A1(KEYINPUT84), .A2(new_n480), .A3(new_n468), .A4(new_n464), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n486), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n483), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n492), .A2(new_n444), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT18), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n495), .A2(KEYINPUT18), .A3(new_n496), .A4(new_n497), .ZN(new_n501));
  INV_X1    g300(.A(new_n444), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n482), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n496), .B(KEYINPUT13), .Z(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT80), .B(G197gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT11), .B(G169gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT12), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n500), .A2(new_n501), .A3(new_n506), .A4(new_n513), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n429), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G127gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(G71gat), .B2(G78gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(KEYINPUT88), .A2(G71gat), .A3(G78gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT88), .B1(G71gat), .B2(G78gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G71gat), .ZN(new_n526));
  INV_X1    g325(.A(G78gat), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT87), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G71gat), .A2(G78gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT88), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(new_n531), .A3(new_n522), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(G57gat), .B(G64gat), .Z(new_n534));
  INV_X1    g333(.A(new_n529), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(KEYINPUT9), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G64gat), .ZN(new_n538));
  INV_X1    g337(.A(G57gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(KEYINPUT89), .ZN(new_n540));
  OR3_X1    g339(.A1(new_n539), .A2(new_n538), .A3(KEYINPUT89), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT9), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n535), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(G231gat), .B(G233gat), .C1(new_n544), .C2(KEYINPUT21), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n537), .A2(new_n543), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT21), .ZN(new_n547));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n519), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n545), .A2(new_n519), .A3(new_n549), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n551), .B2(new_n554), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n439), .B(new_n443), .C1(new_n546), .C2(new_n547), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n558), .A2(KEYINPUT90), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(KEYINPUT90), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n276), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n557), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n555), .B2(new_n556), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G190gat), .B(G218gat), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574));
  OAI211_X1 g373(.A(KEYINPUT17), .B(new_n486), .C1(new_n490), .C2(new_n491), .ZN(new_n575));
  OR2_X1    g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT96), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(KEYINPUT7), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT93), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n581), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT95), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n581), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n584), .A2(KEYINPUT93), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n582), .A2(KEYINPUT7), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n576), .A2(new_n597), .A3(new_n577), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n586), .A2(new_n592), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n577), .A2(KEYINPUT94), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n577), .A2(KEYINPUT94), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT8), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n580), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n598), .A2(new_n592), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n607), .A2(new_n608), .A3(new_n579), .A4(new_n602), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n575), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n482), .A2(KEYINPUT17), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n574), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n610), .B1(new_n482), .B2(KEYINPUT17), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(new_n494), .A3(KEYINPUT97), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n482), .B2(new_n611), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n573), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  AOI211_X1 g421(.A(new_n620), .B(new_n572), .C1(new_n614), .C2(new_n616), .ZN(new_n623));
  XOR2_X1   g422(.A(G134gat), .B(G162gat), .Z(new_n624));
  NOR2_X1   g423(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n622), .A2(new_n623), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n628), .B(new_n629), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n615), .A2(new_n494), .A3(KEYINPUT97), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT97), .B1(new_n615), .B2(new_n494), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n621), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n572), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n617), .A2(new_n621), .A3(new_n573), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n571), .B1(new_n631), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n632), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n622), .B2(new_n623), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n636), .A2(new_n637), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n630), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(KEYINPUT99), .A3(new_n571), .ZN(new_n646));
  XOR2_X1   g445(.A(G120gat), .B(G148gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT101), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n610), .A2(new_n544), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n546), .A2(new_n604), .A3(new_n609), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n651), .A2(new_n658), .A3(new_n652), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n610), .A2(new_n544), .A3(KEYINPUT10), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n654), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT100), .B1(new_n653), .B2(new_n654), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n657), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n654), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n659), .B2(new_n660), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n650), .B1(new_n655), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n641), .A2(new_n646), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n518), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n411), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n436), .A2(new_n442), .ZN(new_n676));
  AND4_X1   g475(.A1(new_n424), .A2(new_n671), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n442), .B1(new_n671), .B2(new_n424), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT42), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(KEYINPUT42), .B2(new_n677), .ZN(G1325gat));
  NAND3_X1  g479(.A1(new_n671), .A2(new_n431), .A3(new_n426), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n259), .A2(new_n682), .A3(new_n265), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n259), .B2(new_n265), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n518), .A2(new_n670), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n681), .B1(new_n431), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n312), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  INV_X1    g489(.A(new_n645), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n571), .A2(new_n668), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n518), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n449), .A3(new_n672), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n691), .A2(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n429), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n571), .B(KEYINPUT104), .ZN(new_n700));
  INV_X1    g499(.A(new_n517), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n700), .A2(new_n701), .A3(new_n668), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n685), .B1(new_n410), .B2(new_n416), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n645), .B1(new_n703), .B2(new_n428), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n699), .B(new_n702), .C1(new_n704), .C2(KEYINPUT44), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n411), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n697), .A2(new_n706), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n694), .A2(new_n450), .A3(new_n424), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT46), .Z(new_n709));
  OAI21_X1  g508(.A(G36gat), .B1(new_n705), .B2(new_n423), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1329gat));
  OAI21_X1  g510(.A(G43gat), .B1(new_n705), .B2(new_n685), .ZN(new_n712));
  INV_X1    g511(.A(new_n693), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n425), .A2(G43gat), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n429), .A2(new_n517), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(KEYINPUT47), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n715), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n717), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI211_X1 g521(.A(KEYINPUT106), .B(KEYINPUT47), .C1(new_n712), .C2(new_n719), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n716), .B1(new_n722), .B2(new_n723), .ZN(G1330gat));
  OAI21_X1  g523(.A(G50gat), .B1(new_n705), .B2(new_n311), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n694), .A2(new_n460), .A3(new_n312), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g527(.A1(new_n703), .A2(new_n428), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n641), .A2(new_n646), .A3(new_n701), .A4(new_n668), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT107), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n729), .A2(KEYINPUT108), .A3(new_n731), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n672), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g537(.A1(new_n736), .A2(new_n424), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  INV_X1    g542(.A(new_n685), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n734), .A2(new_n744), .A3(new_n735), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G71gat), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n734), .A2(new_n526), .A3(new_n426), .A4(new_n735), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1334gat));
  NAND2_X1  g549(.A1(new_n736), .A2(new_n312), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g551(.A1(new_n517), .A2(new_n571), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n704), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n704), .A2(KEYINPUT51), .A3(new_n753), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n588), .A2(new_n590), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n672), .A2(new_n759), .A3(new_n668), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n517), .A2(new_n571), .A3(new_n669), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n699), .B(new_n763), .C1(new_n704), .C2(KEYINPUT44), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n411), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n765), .B2(new_n759), .ZN(G1336gat));
  NAND4_X1  g565(.A1(new_n758), .A2(new_n591), .A3(new_n424), .A4(new_n668), .ZN(new_n767));
  OAI21_X1  g566(.A(G92gat), .B1(new_n764), .B2(new_n423), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(G1337gat));
  AOI21_X1  g573(.A(new_n669), .B1(new_n756), .B2(new_n757), .ZN(new_n775));
  INV_X1    g574(.A(G99gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n776), .A3(new_n426), .ZN(new_n777));
  OAI21_X1  g576(.A(G99gat), .B1(new_n764), .B2(new_n685), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1338gat));
  NOR2_X1   g578(.A1(new_n311), .A2(G106gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT112), .B1(new_n764), .B2(new_n311), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n764), .A2(KEYINPUT112), .A3(new_n311), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n781), .B(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G106gat), .B1(new_n764), .B2(new_n311), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n788), .B2(new_n782), .ZN(G1339gat));
  AND4_X1   g588(.A1(new_n701), .A2(new_n641), .A3(new_n669), .A4(new_n646), .ZN(new_n790));
  INV_X1    g589(.A(new_n664), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n666), .A2(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n650), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n659), .A2(new_n665), .A3(new_n660), .ZN(new_n795));
  AND4_X1   g594(.A1(KEYINPUT113), .A2(new_n662), .A3(KEYINPUT54), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n792), .B1(new_n661), .B2(new_n654), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT113), .B1(new_n797), .B2(new_n795), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n662), .A2(KEYINPUT54), .A3(new_n795), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n797), .A2(KEYINPUT113), .A3(new_n795), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(KEYINPUT114), .A3(new_n794), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n791), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n496), .B1(new_n495), .B2(new_n497), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n504), .A2(new_n505), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n512), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n512), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n812), .A2(new_n516), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n793), .A2(new_n650), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n806), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n808), .A2(new_n691), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  AND4_X1   g620(.A1(new_n516), .A2(new_n668), .A3(new_n812), .A4(new_n814), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n818), .A2(new_n819), .B1(new_n515), .B2(new_n516), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n808), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n821), .B1(new_n824), .B2(new_n691), .ZN(new_n825));
  INV_X1    g624(.A(new_n700), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n790), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n411), .ZN(new_n828));
  INV_X1    g627(.A(new_n420), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT116), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n424), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(KEYINPUT116), .A3(new_n829), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n831), .A2(KEYINPUT117), .A3(new_n832), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n701), .A2(G113gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n827), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n311), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n423), .A2(new_n672), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n841), .A2(new_n425), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n237), .B1(new_n843), .B2(new_n517), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(KEYINPUT118), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  INV_X1    g646(.A(new_n838), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n848), .B1(new_n835), .B2(new_n836), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n847), .B1(new_n849), .B2(new_n844), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n846), .A2(new_n850), .ZN(G1340gat));
  NAND3_X1  g650(.A1(new_n837), .A2(new_n238), .A3(new_n668), .ZN(new_n852));
  INV_X1    g651(.A(new_n843), .ZN(new_n853));
  OAI21_X1  g652(.A(G120gat), .B1(new_n853), .B2(new_n669), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n853), .B2(new_n826), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n571), .A2(new_n519), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n833), .B2(new_n857), .ZN(G1342gat));
  OR3_X1    g657(.A1(new_n833), .A2(G134gat), .A3(new_n645), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n853), .B2(new_n645), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(G1343gat));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  INV_X1    g664(.A(new_n571), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n790), .B1(new_n825), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n311), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n865), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n868), .B1(new_n827), .B2(new_n311), .ZN(new_n872));
  INV_X1    g671(.A(new_n822), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT114), .B1(new_n806), .B2(new_n794), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n650), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n800), .B(new_n875), .C1(new_n804), .C2(new_n805), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n664), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n816), .B1(new_n804), .B2(new_n805), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n517), .B1(KEYINPUT55), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n873), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n645), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n571), .B1(new_n881), .B2(new_n821), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT119), .B(new_n869), .C1(new_n882), .C2(new_n790), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n871), .A2(new_n872), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n744), .A2(new_n842), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n517), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n284), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR4_X1   g687(.A1(new_n683), .A2(new_n684), .A3(new_n424), .A4(new_n311), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n701), .A2(G141gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n828), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n864), .B1(new_n888), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT121), .B(new_n894), .C1(new_n886), .C2(new_n887), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n828), .A2(new_n889), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n886), .A2(new_n887), .B1(new_n899), .B2(new_n890), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n896), .A2(new_n897), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  OAI221_X1 g702(.A(new_n903), .B1(new_n898), .B2(new_n900), .C1(new_n896), .C2(new_n897), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1344gat));
  NAND3_X1  g704(.A1(new_n899), .A2(new_n282), .A3(new_n668), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n867), .A2(KEYINPUT123), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n311), .B1(new_n867), .B2(KEYINPUT123), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n840), .A2(new_n312), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n868), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n668), .A3(new_n885), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n907), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n884), .A2(new_n885), .ZN(new_n917));
  AOI211_X1 g716(.A(KEYINPUT59), .B(new_n282), .C1(new_n917), .C2(new_n668), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n906), .B1(new_n916), .B2(new_n918), .ZN(G1345gat));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n276), .A3(new_n571), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n917), .A2(new_n700), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n276), .ZN(G1346gat));
  AOI21_X1  g721(.A(G162gat), .B1(new_n899), .B2(new_n691), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n645), .A2(new_n277), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n917), .B2(new_n924), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n423), .A2(new_n672), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n827), .A2(new_n420), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n517), .A3(new_n224), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT124), .Z(new_n930));
  NOR3_X1   g729(.A1(new_n841), .A2(new_n425), .A3(new_n927), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n701), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(new_n933), .ZN(G1348gat));
  OAI21_X1  g733(.A(G176gat), .B1(new_n932), .B2(new_n669), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n928), .A2(new_n213), .A3(new_n668), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1349gat));
  OAI21_X1  g736(.A(G183gat), .B1(new_n932), .B2(new_n826), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n928), .A2(new_n205), .A3(new_n571), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  OAI221_X1 g741(.A(G190gat), .B1(KEYINPUT125), .B2(new_n942), .C1(new_n932), .C2(new_n645), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(KEYINPUT125), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n206), .A3(new_n691), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1351gat));
  NOR2_X1   g746(.A1(new_n744), .A2(new_n927), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n911), .ZN(new_n950));
  AOI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n517), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n913), .A2(new_n949), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n517), .A2(G197gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(G1352gat));
  INV_X1    g753(.A(new_n950), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n955), .A2(G204gat), .A3(new_n669), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT62), .ZN(new_n957));
  INV_X1    g756(.A(new_n952), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n958), .B2(new_n669), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1353gat));
  NOR3_X1   g759(.A1(new_n955), .A2(G211gat), .A3(new_n866), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n571), .B(new_n948), .C1(new_n910), .C2(new_n912), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  INV_X1    g767(.A(G218gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n969), .B1(new_n952), .B2(new_n691), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n950), .A2(new_n969), .A3(new_n691), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n973), .ZN(new_n975));
  OAI21_X1  g774(.A(KEYINPUT127), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(G1355gat));
endmodule


