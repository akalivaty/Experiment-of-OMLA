

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U325 ( .A(KEYINPUT82), .B(n556), .ZN(n540) );
  XNOR2_X1 U326 ( .A(n381), .B(n295), .ZN(n296) );
  XNOR2_X1 U327 ( .A(n424), .B(n296), .ZN(n297) );
  XNOR2_X1 U328 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U329 ( .A(n305), .B(n304), .ZN(n310) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U332 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XNOR2_X1 U333 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n375) );
  XOR2_X1 U334 ( .A(G162GAT), .B(KEYINPUT80), .Z(n294) );
  XNOR2_X1 U335 ( .A(G50GAT), .B(G218GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n424) );
  XOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .Z(n381) );
  AND2_X1 U338 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U339 ( .A(n297), .B(KEYINPUT65), .Z(n305) );
  XOR2_X1 U340 ( .A(G85GAT), .B(G92GAT), .Z(n299) );
  XNOR2_X1 U341 ( .A(G99GAT), .B(G106GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n334) );
  XNOR2_X1 U343 ( .A(n334), .B(KEYINPUT9), .ZN(n303) );
  XOR2_X1 U344 ( .A(KEYINPUT11), .B(KEYINPUT81), .Z(n301) );
  XNOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(KEYINPUT8), .B(KEYINPUT71), .Z(n307) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G29GAT), .ZN(n306) );
  XNOR2_X1 U349 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U350 ( .A(KEYINPUT7), .B(n308), .Z(n322) );
  INV_X1 U351 ( .A(n322), .ZN(n309) );
  XNOR2_X1 U352 ( .A(n310), .B(n309), .ZN(n556) );
  XOR2_X1 U353 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n312) );
  XNOR2_X1 U354 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n311) );
  XNOR2_X1 U355 ( .A(n312), .B(n311), .ZN(n326) );
  XOR2_X1 U356 ( .A(KEYINPUT73), .B(G197GAT), .Z(n314) );
  XNOR2_X1 U357 ( .A(G15GAT), .B(G113GAT), .ZN(n313) );
  XNOR2_X1 U358 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U359 ( .A(n315), .B(G50GAT), .Z(n317) );
  XOR2_X1 U360 ( .A(G169GAT), .B(G8GAT), .Z(n391) );
  XNOR2_X1 U361 ( .A(n391), .B(G36GAT), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U363 ( .A(KEYINPUT72), .B(G1GAT), .Z(n360) );
  XOR2_X1 U364 ( .A(n360), .B(KEYINPUT29), .Z(n319) );
  NAND2_X1 U365 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U367 ( .A(n321), .B(n320), .Z(n324) );
  XOR2_X1 U368 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XNOR2_X1 U369 ( .A(n322), .B(n420), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U371 ( .A(n326), .B(n325), .Z(n559) );
  XOR2_X1 U372 ( .A(KEYINPUT78), .B(KEYINPUT75), .Z(n328) );
  XNOR2_X1 U373 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n327) );
  XOR2_X1 U374 ( .A(n328), .B(n327), .Z(n342) );
  XOR2_X1 U375 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n330) );
  NAND2_X1 U376 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U378 ( .A(n331), .B(KEYINPUT79), .Z(n336) );
  XOR2_X1 U379 ( .A(G78GAT), .B(G148GAT), .Z(n333) );
  XNOR2_X1 U380 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n429) );
  XNOR2_X1 U382 ( .A(n429), .B(n334), .ZN(n335) );
  XNOR2_X1 U383 ( .A(n336), .B(n335), .ZN(n338) );
  XNOR2_X1 U384 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n337) );
  XNOR2_X1 U385 ( .A(n337), .B(KEYINPUT13), .ZN(n358) );
  XOR2_X1 U386 ( .A(n338), .B(n358), .Z(n340) );
  XOR2_X1 U387 ( .A(G120GAT), .B(G71GAT), .Z(n446) );
  XOR2_X1 U388 ( .A(G176GAT), .B(G64GAT), .Z(n380) );
  XNOR2_X1 U389 ( .A(n446), .B(n380), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n342), .B(n341), .ZN(n576) );
  XNOR2_X1 U392 ( .A(n576), .B(KEYINPUT41), .ZN(n561) );
  NOR2_X1 U393 ( .A1(n559), .A2(n561), .ZN(n344) );
  XNOR2_X1 U394 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n365) );
  XOR2_X1 U396 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n346) );
  XNOR2_X1 U397 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n364) );
  XOR2_X1 U399 ( .A(G155GAT), .B(G78GAT), .Z(n348) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(G71GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U402 ( .A(G64GAT), .B(G211GAT), .Z(n350) );
  XNOR2_X1 U403 ( .A(G22GAT), .B(G8GAT), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U405 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U406 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n354) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U409 ( .A(KEYINPUT14), .B(n355), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n359) );
  XOR2_X1 U411 ( .A(n359), .B(n358), .Z(n362) );
  XOR2_X1 U412 ( .A(G15GAT), .B(G127GAT), .Z(n447) );
  XNOR2_X1 U413 ( .A(n360), .B(n447), .ZN(n361) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n567) );
  NAND2_X1 U416 ( .A1(n365), .A2(n567), .ZN(n366) );
  NOR2_X1 U417 ( .A1(n556), .A2(n366), .ZN(n367) );
  XNOR2_X1 U418 ( .A(n367), .B(KEYINPUT47), .ZN(n373) );
  INV_X1 U419 ( .A(n567), .ZN(n579) );
  XNOR2_X1 U420 ( .A(KEYINPUT36), .B(n540), .ZN(n583) );
  NAND2_X1 U421 ( .A1(n579), .A2(n583), .ZN(n369) );
  XOR2_X1 U422 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n371) );
  INV_X1 U424 ( .A(n559), .ZN(n572) );
  NOR2_X1 U425 ( .A1(n572), .A2(n576), .ZN(n370) );
  NAND2_X1 U426 ( .A1(n371), .A2(n370), .ZN(n372) );
  NAND2_X1 U427 ( .A1(n373), .A2(n372), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n527) );
  XNOR2_X1 U429 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n376), .B(G183GAT), .ZN(n377) );
  XOR2_X1 U431 ( .A(n377), .B(KEYINPUT88), .Z(n379) );
  XNOR2_X1 U432 ( .A(KEYINPUT18), .B(KEYINPUT89), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n441) );
  XOR2_X1 U434 ( .A(n381), .B(n380), .Z(n383) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U437 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n385) );
  XNOR2_X1 U438 ( .A(G218GAT), .B(G92GAT), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U440 ( .A(n387), .B(n386), .Z(n393) );
  XOR2_X1 U441 ( .A(KEYINPUT21), .B(G211GAT), .Z(n389) );
  XNOR2_X1 U442 ( .A(KEYINPUT91), .B(G204GAT), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U444 ( .A(G197GAT), .B(n390), .Z(n430) );
  XNOR2_X1 U445 ( .A(n391), .B(n430), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n441), .B(n394), .ZN(n491) );
  NAND2_X1 U448 ( .A1(n527), .A2(n491), .ZN(n396) );
  XOR2_X1 U449 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n416) );
  XOR2_X1 U451 ( .A(KEYINPUT1), .B(G57GAT), .Z(n398) );
  XNOR2_X1 U452 ( .A(G141GAT), .B(G1GAT), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n398), .B(n397), .ZN(n415) );
  XOR2_X1 U454 ( .A(G162GAT), .B(G148GAT), .Z(n400) );
  XNOR2_X1 U455 ( .A(G127GAT), .B(G120GAT), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U457 ( .A(G29GAT), .B(G85GAT), .Z(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n411) );
  XNOR2_X1 U459 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n403), .B(KEYINPUT5), .ZN(n404) );
  XOR2_X1 U461 ( .A(n404), .B(KEYINPUT94), .Z(n409) );
  XNOR2_X1 U462 ( .A(G113GAT), .B(G134GAT), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n405), .B(KEYINPUT0), .ZN(n444) );
  XOR2_X1 U464 ( .A(G155GAT), .B(KEYINPUT3), .Z(n407) );
  XNOR2_X1 U465 ( .A(KEYINPUT92), .B(KEYINPUT2), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n427) );
  XNOR2_X1 U467 ( .A(n444), .B(n427), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n413) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U472 ( .A(n415), .B(n414), .Z(n487) );
  NOR2_X1 U473 ( .A1(n416), .A2(n487), .ZN(n569) );
  XOR2_X1 U474 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n418) );
  XNOR2_X1 U475 ( .A(G106GAT), .B(KEYINPUT90), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U477 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U480 ( .A(n423), .B(KEYINPUT93), .Z(n426) );
  XNOR2_X1 U481 ( .A(n424), .B(KEYINPUT22), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U483 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n466) );
  NAND2_X1 U486 ( .A1(n569), .A2(n466), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n433), .B(KEYINPUT122), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n434), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U489 ( .A(G176GAT), .B(KEYINPUT20), .Z(n436) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U492 ( .A(KEYINPUT87), .B(G99GAT), .Z(n438) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(G190GAT), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n443) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U498 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n529) );
  NAND2_X1 U501 ( .A1(n450), .A2(n529), .ZN(n566) );
  INV_X1 U502 ( .A(n566), .ZN(n451) );
  NAND2_X1 U503 ( .A1(n451), .A2(n540), .ZN(n455) );
  XOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n453) );
  INV_X1 U505 ( .A(n487), .ZN(n511) );
  NOR2_X1 U506 ( .A1(n559), .A2(n576), .ZN(n485) );
  NAND2_X1 U507 ( .A1(n529), .A2(n491), .ZN(n456) );
  NAND2_X1 U508 ( .A1(n466), .A2(n456), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(KEYINPUT25), .ZN(n462) );
  XNOR2_X1 U510 ( .A(KEYINPUT27), .B(KEYINPUT97), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(n491), .ZN(n465) );
  NOR2_X1 U512 ( .A1(n466), .A2(n529), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT26), .ZN(n570) );
  INV_X1 U514 ( .A(n570), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n465), .A2(n460), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U517 ( .A1(n487), .A2(n463), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n464), .B(KEYINPUT98), .ZN(n470) );
  NOR2_X1 U519 ( .A1(n511), .A2(n465), .ZN(n526) );
  XOR2_X1 U520 ( .A(n466), .B(KEYINPUT67), .Z(n467) );
  XNOR2_X1 U521 ( .A(KEYINPUT28), .B(n467), .ZN(n522) );
  NAND2_X1 U522 ( .A1(n526), .A2(n522), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n468), .A2(n529), .ZN(n469) );
  NOR2_X1 U524 ( .A1(n470), .A2(n469), .ZN(n482) );
  NOR2_X1 U525 ( .A1(n540), .A2(n567), .ZN(n471) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(n471), .Z(n472) );
  NOR2_X1 U527 ( .A1(n482), .A2(n472), .ZN(n499) );
  NAND2_X1 U528 ( .A1(n485), .A2(n499), .ZN(n480) );
  NOR2_X1 U529 ( .A1(n511), .A2(n480), .ZN(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT34), .B(n473), .Z(n474) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  INV_X1 U532 ( .A(n491), .ZN(n513) );
  NOR2_X1 U533 ( .A1(n513), .A2(n480), .ZN(n475) );
  XOR2_X1 U534 ( .A(G8GAT), .B(n475), .Z(G1325GAT) );
  INV_X1 U535 ( .A(n529), .ZN(n515) );
  NOR2_X1 U536 ( .A1(n480), .A2(n515), .ZN(n479) );
  XOR2_X1 U537 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n477) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT100), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n522), .A2(n480), .ZN(n481) );
  XOR2_X1 U542 ( .A(G22GAT), .B(n481), .Z(G1327GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n489) );
  NOR2_X1 U544 ( .A1(n579), .A2(n482), .ZN(n483) );
  NAND2_X1 U545 ( .A1(n583), .A2(n483), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(KEYINPUT37), .ZN(n510) );
  NAND2_X1 U547 ( .A1(n510), .A2(n485), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(n486), .Z(n496) );
  NAND2_X1 U549 ( .A1(n487), .A2(n496), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U551 ( .A(G29GAT), .B(n490), .Z(G1328GAT) );
  NAND2_X1 U552 ( .A1(n496), .A2(n491), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n496), .A2(n529), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  XOR2_X1 U558 ( .A(G50GAT), .B(KEYINPUT103), .Z(n498) );
  INV_X1 U559 ( .A(n522), .ZN(n531) );
  NAND2_X1 U560 ( .A1(n531), .A2(n496), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  NOR2_X1 U562 ( .A1(n572), .A2(n561), .ZN(n509) );
  NAND2_X1 U563 ( .A1(n509), .A2(n499), .ZN(n505) );
  NOR2_X1 U564 ( .A1(n511), .A2(n505), .ZN(n500) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n500), .Z(n501) );
  XNOR2_X1 U566 ( .A(KEYINPUT42), .B(n501), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n513), .A2(n505), .ZN(n502) );
  XOR2_X1 U568 ( .A(G64GAT), .B(n502), .Z(G1333GAT) );
  NOR2_X1 U569 ( .A1(n515), .A2(n505), .ZN(n503) );
  XOR2_X1 U570 ( .A(KEYINPUT104), .B(n503), .Z(n504) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U572 ( .A1(n522), .A2(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U575 ( .A(G78GAT), .B(n508), .Z(G1335GAT) );
  NAND2_X1 U576 ( .A1(n510), .A2(n509), .ZN(n521) );
  NOR2_X1 U577 ( .A1(n511), .A2(n521), .ZN(n512) );
  XOR2_X1 U578 ( .A(G85GAT), .B(n512), .Z(G1336GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n521), .ZN(n514) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n521), .ZN(n517) );
  XNOR2_X1 U582 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(n518), .ZN(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(n524) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U589 ( .A(n524), .B(n523), .Z(n525) );
  XNOR2_X1 U590 ( .A(KEYINPUT108), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U591 ( .A(G113GAT), .B(KEYINPUT113), .Z(n533) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT112), .B(n528), .Z(n545) );
  NAND2_X1 U594 ( .A1(n529), .A2(n545), .ZN(n530) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n541), .A2(n572), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  INV_X1 U599 ( .A(n561), .ZN(n548) );
  NAND2_X1 U600 ( .A1(n541), .A2(n548), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n539) );
  XOR2_X1 U603 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n537) );
  NAND2_X1 U604 ( .A1(n541), .A2(n579), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n545), .A2(n570), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT117), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n572), .A2(n555), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n552) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT118), .Z(n550) );
  NAND2_X1 U617 ( .A1(n555), .A2(n548), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  XOR2_X1 U620 ( .A(G155GAT), .B(KEYINPUT119), .Z(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n579), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(KEYINPUT120), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n558), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n566), .ZN(n560) );
  XOR2_X1 U627 ( .A(G169GAT), .B(n560), .Z(G1348GAT) );
  NOR2_X1 U628 ( .A1(n566), .A2(n561), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n563) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  NAND2_X1 U636 ( .A1(n569), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT125), .B(n571), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n582), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U642 ( .A1(n582), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

