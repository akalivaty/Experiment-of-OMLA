//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT75), .A2(G104), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT75), .A2(G104), .ZN(new_n190));
  OAI22_X1  g004(.A1(new_n189), .A2(new_n190), .B1(KEYINPUT3), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(G101), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT3), .A2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G104), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n191), .A2(new_n192), .A3(new_n193), .A4(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n189), .B2(new_n190), .ZN(new_n198));
  NAND2_X1  g012(.A1(G104), .A2(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(G101), .A3(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT68), .B1(new_n202), .B2(G119), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G116), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G119), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n203), .A2(new_n206), .A3(KEYINPUT5), .A4(new_n207), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n202), .A2(KEYINPUT5), .A3(G119), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(G113), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G113), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT2), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G113), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n215), .A2(new_n207), .A3(new_n206), .A4(new_n203), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n210), .A2(KEYINPUT82), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT82), .B1(new_n210), .B2(new_n216), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n201), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT83), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n210), .A2(new_n216), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n197), .A2(new_n200), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n224), .B(new_n201), .C1(new_n217), .C2(new_n218), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n220), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G110), .B(G122), .ZN(new_n227));
  XOR2_X1   g041(.A(new_n227), .B(KEYINPUT80), .Z(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT8), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n226), .A2(KEYINPUT84), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT84), .B1(new_n226), .B2(new_n229), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n201), .A2(new_n216), .A3(new_n210), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n191), .A2(new_n193), .A3(new_n196), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G101), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n236), .A3(G101), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n212), .A2(new_n214), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n241), .A2(KEYINPUT69), .A3(new_n216), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT69), .B1(new_n241), .B2(new_n216), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n232), .B(new_n228), .C1(new_n238), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G143), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT65), .B1(new_n248), .B2(G146), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n246), .A3(G143), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n247), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n248), .A2(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n246), .A2(G143), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT0), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT64), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(KEYINPUT0), .B2(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n252), .A2(new_n253), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n255), .ZN(new_n266));
  OAI211_X1 g080(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n248), .C2(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G128), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT67), .B1(new_n255), .B2(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n249), .A2(new_n251), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G128), .A4(new_n254), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n264), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G224), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT81), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT7), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n265), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n265), .B2(new_n274), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT85), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT85), .ZN(new_n283));
  AOI211_X1 g097(.A(new_n283), .B(new_n279), .C1(new_n265), .C2(new_n274), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n245), .B(new_n280), .C1(new_n282), .C2(new_n284), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n230), .A2(new_n231), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n232), .B1(new_n238), .B2(new_n244), .ZN(new_n287));
  INV_X1    g101(.A(new_n228), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT6), .A3(new_n245), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT6), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(new_n291), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n265), .A2(new_n274), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(new_n277), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n188), .B1(new_n286), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n226), .A2(new_n229), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n226), .A2(KEYINPUT84), .A3(new_n229), .ZN(new_n302));
  INV_X1    g116(.A(new_n285), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n304), .A2(new_n296), .A3(new_n187), .A4(new_n295), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT79), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n275), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT70), .A2(G953), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G237), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(G214), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(G143), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT18), .ZN(new_n318));
  INV_X1    g132(.A(G131), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(G125), .B(G140), .Z(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(G146), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n316), .B(new_n248), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G131), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n320), .B(new_n322), .C1(new_n318), .C2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n321), .B(KEYINPUT19), .Z(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n246), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n317), .A2(new_n319), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n323), .A2(G131), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OR3_X1    g144(.A1(new_n264), .A2(KEYINPUT16), .A3(G140), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT16), .ZN(new_n332));
  OAI211_X1 g146(.A(G146), .B(new_n331), .C1(new_n321), .C2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT73), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n325), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G113), .B(G122), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n336), .B(G104), .Z(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n317), .A2(new_n319), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT17), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n324), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n328), .A2(KEYINPUT17), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n331), .B1(new_n321), .B2(new_n332), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n246), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n342), .A2(new_n343), .A3(new_n333), .A4(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n337), .A3(new_n325), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G475), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(new_n296), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT20), .ZN(new_n351));
  AOI21_X1  g165(.A(G475), .B1(new_n339), .B2(new_n347), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n296), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n347), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n337), .B1(new_n346), .B2(new_n325), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n296), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G475), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n258), .A2(G143), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT13), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT86), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n360), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT87), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n258), .A2(G143), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n362), .A3(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n248), .A2(G128), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n360), .A2(new_n362), .A3(new_n364), .A4(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G134), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G134), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n369), .A2(new_n367), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n202), .A2(G122), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n202), .A2(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G107), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n195), .A3(new_n381), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n373), .A2(KEYINPUT88), .A3(G134), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n376), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n379), .B1(KEYINPUT14), .B2(new_n381), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(KEYINPUT90), .C1(KEYINPUT14), .C2(new_n381), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n389), .B(G107), .C1(KEYINPUT90), .C2(new_n388), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n377), .B1(new_n369), .B2(new_n367), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n378), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n392), .A2(KEYINPUT89), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(KEYINPUT89), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n390), .B(new_n384), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n387), .A2(new_n395), .ZN(new_n396));
  XOR2_X1   g210(.A(KEYINPUT9), .B(G234), .Z(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G217), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n398), .A2(new_n399), .A3(G953), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n387), .A2(new_n395), .A3(new_n400), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n296), .ZN(new_n405));
  INV_X1    g219(.A(G478), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(KEYINPUT15), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n405), .B(new_n407), .Z(new_n408));
  INV_X1    g222(.A(G952), .ZN(new_n409));
  AOI211_X1 g223(.A(G953), .B(new_n409), .C1(G234), .C2(G237), .ZN(new_n410));
  AOI211_X1 g224(.A(new_n296), .B(new_n314), .C1(G234), .C2(G237), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT21), .B(G898), .Z(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n410), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AND4_X1   g229(.A1(new_n355), .A2(new_n359), .A3(new_n408), .A4(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G221), .B1(new_n398), .B2(G902), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G469), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT11), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n377), .B2(G137), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n377), .A2(G137), .ZN(new_n422));
  INV_X1    g236(.A(G137), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT11), .A3(G134), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G131), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n421), .A2(new_n424), .A3(new_n319), .A4(new_n422), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n428), .A2(KEYINPUT77), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n270), .A2(new_n273), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n201), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n258), .B1(new_n255), .B2(KEYINPUT1), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n252), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n222), .B1(new_n273), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n429), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT12), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n314), .A2(G227), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G140), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT10), .ZN(new_n441));
  INV_X1    g255(.A(new_n273), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(new_n433), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n443), .B2(new_n222), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n270), .A2(new_n273), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n197), .A2(KEYINPUT10), .A3(new_n200), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT76), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n235), .A2(new_n263), .A3(new_n237), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT76), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n201), .A2(new_n449), .A3(new_n430), .A4(KEYINPUT10), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n444), .A2(new_n447), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n440), .B1(new_n451), .B2(new_n428), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n437), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n447), .A2(new_n450), .ZN(new_n454));
  INV_X1    g268(.A(new_n428), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n448), .A4(new_n444), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n428), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n440), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n419), .B(new_n296), .C1(new_n453), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n419), .A2(new_n296), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n440), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n451), .A2(new_n428), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n463), .B1(new_n437), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n456), .A2(new_n457), .A3(new_n440), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n465), .A2(KEYINPUT78), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT78), .B1(new_n465), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g282(.A(G469), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n418), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n310), .A2(new_n416), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT32), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n428), .A2(new_n263), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT66), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n423), .A2(G134), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n422), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G131), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n430), .A2(new_n427), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n428), .A2(new_n263), .A3(KEYINPUT66), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n477), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n244), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n270), .A2(new_n273), .B1(G131), .B2(new_n479), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n486), .A2(new_n427), .B1(new_n428), .B2(new_n263), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n244), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT28), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT28), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n487), .B2(new_n244), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n485), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(G101), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n314), .A2(G210), .A3(new_n315), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n483), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n487), .A2(KEYINPUT30), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n484), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT31), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n488), .A4(new_n496), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n488), .A3(new_n496), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT31), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT71), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT71), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT31), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n505), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(G472), .A2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n474), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT31), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n509), .B1(new_n506), .B2(KEYINPUT31), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n498), .B(new_n504), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(KEYINPUT32), .A3(new_n512), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n502), .A2(new_n488), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n496), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT29), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n489), .A2(new_n491), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n487), .A2(new_n244), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n496), .B1(new_n492), .B2(KEYINPUT29), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n522), .B(new_n296), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G472), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n514), .A2(new_n518), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n205), .A2(KEYINPUT23), .A3(G128), .ZN(new_n531));
  XNOR2_X1  g345(.A(G119), .B(G128), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(KEYINPUT23), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT24), .B(G110), .Z(new_n534));
  OAI22_X1  g348(.A1(new_n533), .A2(G110), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(G146), .B2(new_n321), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n334), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n532), .ZN(new_n538));
  XOR2_X1   g352(.A(new_n538), .B(KEYINPUT72), .Z(new_n539));
  NAND2_X1  g353(.A1(new_n345), .A2(new_n333), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n533), .A2(G110), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n314), .A2(G221), .A3(G234), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT22), .Z(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G137), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n544), .B(KEYINPUT22), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n423), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n546), .A2(new_n548), .A3(KEYINPUT74), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n543), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n537), .A2(new_n549), .A3(new_n550), .A4(new_n542), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n530), .B1(new_n555), .B2(new_n296), .ZN(new_n556));
  AOI211_X1 g370(.A(KEYINPUT25), .B(G902), .C1(new_n553), .C2(new_n554), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n399), .B1(G234), .B2(new_n296), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G902), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n558), .A2(new_n559), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n529), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n310), .A2(new_n416), .A3(KEYINPUT91), .A4(new_n470), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n473), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(G101), .ZN(G3));
  OAI21_X1  g379(.A(G472), .B1(new_n511), .B2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n517), .A2(new_n512), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n569), .A2(new_n561), .A3(new_n470), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n298), .A2(new_n571), .A3(new_n305), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(KEYINPUT92), .B(new_n188), .C1(new_n286), .C2(new_n297), .ZN(new_n574));
  INV_X1    g388(.A(new_n309), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT33), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n404), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n406), .A2(G902), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n400), .B1(new_n387), .B2(new_n395), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT93), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n403), .A2(KEYINPUT94), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n387), .A2(new_n395), .A3(new_n584), .A4(new_n400), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(KEYINPUT33), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n579), .B(new_n580), .C1(new_n582), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT95), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT93), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n581), .B(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n583), .A2(KEYINPUT33), .A3(new_n585), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT95), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n579), .A4(new_n580), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n405), .A2(new_n406), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n588), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n351), .A2(new_n354), .B1(G475), .B2(new_n358), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n570), .A2(new_n415), .A3(new_n577), .A4(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT34), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G104), .ZN(G6));
  AOI21_X1  g416(.A(new_n408), .B1(G475), .B2(new_n358), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n604));
  AND4_X1   g418(.A1(new_n353), .A2(new_n348), .A3(new_n349), .A4(new_n296), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n353), .B1(new_n352), .B2(new_n296), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n351), .A2(KEYINPUT96), .A3(new_n354), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n577), .A2(new_n603), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n414), .B(KEYINPUT97), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n570), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT98), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT35), .B(G107), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NAND2_X1  g430(.A1(new_n555), .A2(new_n296), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT25), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n555), .A2(new_n530), .A3(new_n296), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n559), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n549), .A2(KEYINPUT36), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(new_n543), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n560), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n473), .A2(new_n563), .A3(new_n569), .A4(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n625), .B(KEYINPUT37), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G110), .ZN(G12));
  INV_X1    g441(.A(G900), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n410), .B1(new_n411), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n607), .A2(new_n608), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n603), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n529), .A2(new_n470), .ZN(new_n633));
  AND4_X1   g447(.A1(new_n575), .A2(new_n624), .A3(new_n572), .A4(new_n574), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G128), .ZN(G30));
  XOR2_X1   g450(.A(new_n629), .B(KEYINPUT39), .Z(new_n637));
  NAND2_X1  g451(.A1(new_n470), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n638), .A2(KEYINPUT40), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(KEYINPUT40), .ZN(new_n640));
  NOR4_X1   g454(.A1(new_n639), .A2(new_n640), .A3(new_n309), .A4(new_n624), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n306), .B(KEYINPUT99), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT38), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n519), .A2(new_n496), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n524), .A2(new_n488), .A3(new_n497), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n296), .ZN(new_n648));
  OAI21_X1  g462(.A(G472), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n514), .A2(new_n518), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n598), .A2(new_n408), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n641), .A2(new_n644), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G143), .ZN(G45));
  OAI21_X1  g467(.A(new_n359), .B1(new_n605), .B2(new_n606), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n596), .A2(new_n654), .A3(new_n630), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n634), .A2(new_n529), .A3(new_n655), .A4(new_n470), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n633), .A2(KEYINPUT100), .A3(new_n634), .A4(new_n655), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G146), .ZN(G48));
  OAI21_X1  g475(.A(new_n296), .B1(new_n453), .B2(new_n458), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G469), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n417), .A3(new_n459), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n573), .A2(new_n576), .A3(new_n664), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n561), .A2(new_n596), .A3(new_n654), .A4(new_n415), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n529), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT101), .A4(new_n529), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT41), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G113), .ZN(G15));
  NOR2_X1   g487(.A1(new_n664), .A2(new_n611), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n610), .A2(new_n562), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G116), .ZN(G18));
  NAND4_X1  g490(.A1(new_n665), .A2(new_n529), .A3(new_n416), .A4(new_n624), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G119), .ZN(G21));
  NAND2_X1  g492(.A1(new_n566), .A2(KEYINPUT102), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n523), .A2(new_n524), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n504), .B1(new_n680), .B2(new_n496), .ZN(new_n681));
  INV_X1    g495(.A(new_n507), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n512), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n684), .B(G472), .C1(new_n511), .C2(G902), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n561), .A2(new_n679), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n577), .A2(new_n651), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n674), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G122), .ZN(G24));
  INV_X1    g503(.A(new_n665), .ZN(new_n690));
  INV_X1    g504(.A(new_n655), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n679), .A2(new_n624), .A3(new_n683), .A4(new_n685), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G125), .ZN(G27));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n698));
  INV_X1    g512(.A(new_n461), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n465), .A2(G469), .A3(new_n466), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n459), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n418), .A2(new_n309), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n701), .A2(new_n298), .A3(new_n305), .A4(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n529), .B(new_n561), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n698), .B1(new_n706), .B2(new_n691), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n703), .B(KEYINPUT104), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n562), .A2(new_n709), .A3(KEYINPUT105), .A4(new_n655), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n561), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT106), .B1(new_n514), .B2(new_n518), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(KEYINPUT106), .B2(new_n514), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n712), .B1(new_n714), .B2(new_n528), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(KEYINPUT42), .A3(new_n655), .A4(new_n709), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G131), .ZN(G33));
  NAND3_X1  g532(.A1(new_n632), .A2(new_n562), .A3(new_n709), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G134), .ZN(G36));
  NAND2_X1  g534(.A1(new_n598), .A2(new_n596), .ZN(new_n721));
  NAND2_X1  g535(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n722));
  OR2_X1    g536(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n598), .A2(new_n596), .A3(KEYINPUT43), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n721), .A2(KEYINPUT109), .A3(new_n722), .A4(new_n723), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n726), .A2(KEYINPUT110), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n729), .A2(new_n568), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n731), .A2(new_n732), .B1(new_n620), .B2(new_n623), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT111), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n730), .A2(new_n733), .A3(new_n737), .A4(KEYINPUT44), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n306), .A2(new_n309), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n465), .A2(KEYINPUT45), .A3(new_n466), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n467), .A2(new_n468), .ZN(new_n744));
  OAI211_X1 g558(.A(G469), .B(new_n743), .C1(new_n744), .C2(KEYINPUT45), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n699), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n699), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n459), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n417), .A3(new_n637), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT107), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n735), .B2(new_n734), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n736), .A2(new_n738), .A3(KEYINPUT112), .A4(new_n739), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n742), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  NAND2_X1  g570(.A1(new_n750), .A2(new_n417), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n750), .A2(KEYINPUT47), .A3(new_n417), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n655), .A2(new_n739), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n762), .A2(new_n529), .A3(new_n561), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT113), .Z(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  NOR2_X1   g580(.A1(new_n650), .A2(new_n712), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n663), .A2(new_n459), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT49), .Z(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n769), .A3(new_n702), .ZN(new_n770));
  OR3_X1    g584(.A1(new_n644), .A2(new_n721), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n624), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n417), .A2(new_n650), .A3(new_n772), .A4(new_n701), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n630), .A3(new_n687), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n696), .A2(new_n660), .A3(new_n635), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n693), .B(KEYINPUT103), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n778), .B1(new_n779), .B2(new_n692), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(KEYINPUT52), .A3(new_n660), .A4(new_n774), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n709), .A2(new_n655), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n408), .A2(new_n359), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n739), .A2(new_n624), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n788), .A2(new_n633), .A3(new_n631), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n719), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n786), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(new_n717), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n307), .A2(new_n309), .A3(new_n611), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n596), .A2(new_n654), .A3(KEYINPUT114), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT114), .B1(new_n596), .B2(new_n654), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT115), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n794), .B(new_n799), .C1(new_n795), .C2(new_n796), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n570), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n654), .A2(new_n408), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT116), .Z(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n570), .A3(new_n794), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n801), .A2(new_n804), .A3(new_n625), .A4(new_n564), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n671), .A2(new_n688), .A3(new_n675), .A4(new_n677), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n782), .A2(new_n793), .A3(KEYINPUT53), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n564), .A2(new_n801), .A3(new_n804), .A4(new_n625), .ZN(new_n811));
  INV_X1    g625(.A(new_n806), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n812), .A3(new_n792), .A4(new_n717), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT118), .A3(KEYINPUT53), .A4(new_n782), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n813), .A2(KEYINPUT117), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n782), .B1(new_n813), .B2(KEYINPUT117), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT54), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n777), .A2(new_n781), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n817), .B1(new_n823), .B2(new_n813), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n808), .ZN(new_n826));
  OAI211_X1 g640(.A(KEYINPUT119), .B(new_n817), .C1(new_n823), .C2(new_n813), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n768), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n410), .A2(new_n307), .A3(new_n831), .A4(new_n702), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n767), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT121), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(KEYINPUT121), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n599), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n831), .A2(new_n418), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n759), .A2(new_n760), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n731), .A2(new_n410), .A3(new_n686), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n739), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT120), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n842), .A2(KEYINPUT120), .ZN(new_n844));
  INV_X1    g658(.A(new_n664), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n643), .A2(new_n309), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n843), .B(new_n844), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n731), .A2(new_n832), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n779), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n834), .A2(new_n598), .A3(new_n597), .A4(new_n835), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n841), .A2(new_n848), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n846), .A2(new_n843), .A3(new_n847), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n837), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n409), .A2(G953), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n852), .A2(new_n853), .A3(new_n837), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n822), .A2(new_n830), .A3(new_n836), .A4(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n840), .A2(new_n665), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n849), .A2(new_n715), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT48), .Z(new_n862));
  NOR3_X1   g676(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(G952), .A2(G953), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n771), .B1(new_n863), .B2(new_n864), .ZN(G75));
  NAND2_X1  g679(.A1(new_n290), .A2(new_n292), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n294), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT55), .Z(new_n868));
  NAND3_X1  g682(.A1(new_n826), .A2(G902), .A3(new_n827), .ZN(new_n869));
  INV_X1    g683(.A(G210), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n868), .B1(new_n871), .B2(KEYINPUT56), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n314), .A2(G952), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n826), .A2(KEYINPUT122), .A3(G902), .A4(new_n827), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n188), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n868), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n877), .A2(new_n188), .A3(new_n879), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT56), .B1(new_n883), .B2(KEYINPUT123), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n875), .B1(new_n882), .B2(new_n884), .ZN(G51));
  NAND2_X1  g699(.A1(new_n699), .A2(KEYINPUT57), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n828), .A2(new_n829), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT54), .B1(new_n826), .B2(new_n827), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n699), .A2(KEYINPUT57), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n889), .A2(new_n890), .B1(new_n458), .B2(new_n453), .ZN(new_n891));
  INV_X1    g705(.A(new_n745), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n877), .A2(new_n892), .A3(new_n879), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n873), .B1(new_n891), .B2(new_n893), .ZN(G54));
  NAND4_X1  g708(.A1(new_n877), .A2(KEYINPUT58), .A3(G475), .A4(new_n879), .ZN(new_n895));
  INV_X1    g709(.A(new_n348), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n873), .ZN(G60));
  NAND2_X1  g713(.A1(new_n592), .A2(new_n579), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n888), .B1(KEYINPUT54), .B2(new_n821), .ZN(new_n901));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT59), .Z(new_n903));
  OAI21_X1  g717(.A(new_n900), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n900), .ZN(new_n905));
  INV_X1    g719(.A(new_n903), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n905), .B(new_n906), .C1(new_n887), .C2(new_n888), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n904), .A2(new_n874), .A3(new_n907), .ZN(G63));
  AND2_X1   g722(.A1(new_n826), .A2(new_n827), .ZN(new_n909));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT60), .Z(new_n911));
  NAND4_X1  g725(.A1(new_n909), .A2(KEYINPUT124), .A3(new_n622), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n826), .A2(new_n827), .A3(new_n911), .ZN(new_n913));
  INV_X1    g727(.A(new_n555), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n873), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n826), .A2(new_n622), .A3(new_n827), .A4(new_n911), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n912), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G66));
  INV_X1    g735(.A(G224), .ZN(new_n922));
  OAI21_X1  g736(.A(G953), .B1(new_n413), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n314), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n807), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n866), .B1(G898), .B2(new_n314), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT125), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n925), .B(new_n927), .ZN(G69));
  NAND2_X1  g742(.A1(new_n924), .A2(G227), .ZN(new_n929));
  INV_X1    g743(.A(new_n752), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n687), .A3(new_n715), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n717), .A2(new_n719), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT127), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n761), .B2(new_n764), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n780), .A2(new_n660), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n755), .A2(KEYINPUT126), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT126), .B1(new_n755), .B2(new_n935), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n931), .B(new_n934), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n929), .B1(new_n938), .B2(new_n924), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n500), .A2(new_n501), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n326), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n924), .A2(new_n628), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n935), .A2(new_n652), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n803), .A2(new_n796), .A3(new_n795), .ZN(new_n948));
  INV_X1    g762(.A(new_n638), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n562), .A3(new_n949), .A4(new_n739), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n755), .A2(new_n947), .A3(new_n765), .A4(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n929), .B(new_n941), .C1(new_n951), .C2(new_n924), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n943), .A2(new_n944), .A3(new_n952), .ZN(G72));
  NAND2_X1  g767(.A1(G472), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT63), .Z(new_n955));
  INV_X1    g769(.A(new_n807), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n646), .ZN(new_n958));
  INV_X1    g772(.A(new_n520), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n821), .A2(new_n959), .A3(new_n645), .A4(new_n955), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n874), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n955), .B1(new_n938), .B2(new_n956), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n520), .B2(new_n962), .ZN(G57));
endmodule


