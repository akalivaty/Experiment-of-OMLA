

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745;

  XNOR2_X1 U373 ( .A(n577), .B(n576), .ZN(n743) );
  BUF_X1 U374 ( .A(n516), .Z(n477) );
  NAND2_X1 U375 ( .A1(n354), .A2(n390), .ZN(n542) );
  AND2_X1 U376 ( .A1(n422), .A2(G224), .ZN(n423) );
  INV_X1 U377 ( .A(KEYINPUT64), .ZN(n360) );
  XNOR2_X1 U378 ( .A(n427), .B(n428), .ZN(n434) );
  NAND2_X1 U379 ( .A1(n471), .A2(n687), .ZN(n692) );
  NOR2_X1 U380 ( .A1(n692), .A2(n690), .ZN(n473) );
  XOR2_X1 U381 ( .A(G104), .B(G107), .Z(n351) );
  OR2_X2 U382 ( .A1(n544), .A2(n543), .ZN(n547) );
  NOR2_X2 U383 ( .A1(n630), .A2(n578), .ZN(n579) );
  XNOR2_X2 U384 ( .A(n563), .B(KEYINPUT35), .ZN(n630) );
  NAND2_X1 U385 ( .A1(n636), .A2(n744), .ZN(n485) );
  NAND2_X1 U386 ( .A1(n583), .A2(n565), .ZN(n568) );
  INV_X1 U387 ( .A(n542), .ZN(n588) );
  INV_X1 U388 ( .A(n534), .ZN(n543) );
  AND2_X1 U389 ( .A1(n601), .A2(n600), .ZN(n606) );
  INV_X1 U390 ( .A(n352), .ZN(n664) );
  AND2_X1 U391 ( .A1(n421), .A2(n420), .ZN(n505) );
  OR2_X1 U392 ( .A1(n477), .A2(n489), .ZN(n419) );
  BUF_X1 U393 ( .A(n477), .Z(n677) );
  XNOR2_X1 U394 ( .A(n527), .B(n526), .ZN(n534) );
  OR2_X1 U395 ( .A1(n648), .A2(G902), .ZN(n400) );
  XNOR2_X1 U396 ( .A(n360), .B(G953), .ZN(n422) );
  XOR2_X1 U397 ( .A(G146), .B(G125), .Z(n424) );
  XNOR2_X2 U398 ( .A(n598), .B(n353), .ZN(n352) );
  XOR2_X1 U399 ( .A(n597), .B(KEYINPUT45), .Z(n353) );
  XNOR2_X2 U400 ( .A(n620), .B(G146), .ZN(n413) );
  NOR2_X1 U401 ( .A1(n602), .A2(n665), .ZN(n603) );
  NAND2_X1 U402 ( .A1(n448), .A2(G221), .ZN(n374) );
  XNOR2_X1 U403 ( .A(n566), .B(KEYINPUT22), .ZN(n567) );
  BUF_X1 U404 ( .A(n422), .Z(n622) );
  XNOR2_X1 U405 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U406 ( .A(n429), .B(KEYINPUT16), .ZN(n430) );
  AND2_X2 U407 ( .A1(n606), .A2(n670), .ZN(n652) );
  NOR2_X1 U408 ( .A1(n622), .A2(G952), .ZN(n659) );
  XOR2_X1 U409 ( .A(n387), .B(n386), .Z(n354) );
  XOR2_X1 U410 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n355) );
  XNOR2_X2 U411 ( .A(n400), .B(n399), .ZN(n527) );
  NOR2_X1 U412 ( .A1(n533), .A2(n537), .ZN(n525) );
  AND2_X1 U413 ( .A1(n475), .A2(n588), .ZN(n356) );
  INV_X1 U414 ( .A(KEYINPUT107), .ZN(n522) );
  XNOR2_X1 U415 ( .A(n667), .B(n666), .ZN(n668) );
  BUF_X1 U416 ( .A(n607), .Z(n608) );
  BUF_X1 U417 ( .A(n617), .Z(n663) );
  BUF_X1 U418 ( .A(n652), .Z(n646) );
  BUF_X1 U419 ( .A(n534), .Z(n585) );
  INV_X1 U420 ( .A(n659), .ZN(n612) );
  NAND2_X1 U421 ( .A1(G234), .A2(G237), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n357), .B(KEYINPUT14), .ZN(n358) );
  XNOR2_X1 U423 ( .A(KEYINPUT76), .B(n358), .ZN(n365) );
  NAND2_X1 U424 ( .A1(n365), .A2(G902), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n359), .B(KEYINPUT92), .ZN(n550) );
  NOR2_X1 U426 ( .A1(n550), .A2(n622), .ZN(n362) );
  INV_X1 U427 ( .A(KEYINPUT105), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n364) );
  INV_X1 U429 ( .A(G900), .ZN(n363) );
  NAND2_X1 U430 ( .A1(n364), .A2(n363), .ZN(n367) );
  NAND2_X1 U431 ( .A1(G952), .A2(n365), .ZN(n702) );
  NOR2_X1 U432 ( .A1(G953), .A2(n702), .ZN(n366) );
  XOR2_X1 U433 ( .A(KEYINPUT90), .B(n366), .Z(n552) );
  NAND2_X1 U434 ( .A1(n367), .A2(n552), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n368), .B(KEYINPUT82), .ZN(n475) );
  NAND2_X1 U436 ( .A1(n422), .A2(G234), .ZN(n370) );
  INV_X1 U437 ( .A(KEYINPUT8), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n448) );
  XNOR2_X1 U439 ( .A(G110), .B(KEYINPUT23), .ZN(n372) );
  XNOR2_X1 U440 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n371) );
  XNOR2_X1 U441 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n374), .B(n373), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n424), .B(KEYINPUT10), .ZN(n619) );
  INV_X1 U444 ( .A(n619), .ZN(n378) );
  XNOR2_X1 U445 ( .A(G128), .B(G119), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n375), .B(KEYINPUT96), .ZN(n376) );
  XNOR2_X1 U447 ( .A(G137), .B(G140), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n376), .B(n393), .ZN(n377) );
  XNOR2_X1 U449 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U450 ( .A(n380), .B(n379), .ZN(n639) );
  INV_X1 U451 ( .A(G902), .ZN(n465) );
  NAND2_X1 U452 ( .A1(n639), .A2(n465), .ZN(n387) );
  XNOR2_X1 U453 ( .A(G902), .B(KEYINPUT89), .ZN(n381) );
  XNOR2_X1 U454 ( .A(n381), .B(KEYINPUT15), .ZN(n600) );
  INV_X1 U455 ( .A(n600), .ZN(n435) );
  NAND2_X1 U456 ( .A1(G234), .A2(n435), .ZN(n382) );
  XNOR2_X1 U457 ( .A(KEYINPUT20), .B(n382), .ZN(n388) );
  NAND2_X1 U458 ( .A1(n388), .A2(G217), .ZN(n385) );
  XOR2_X1 U459 ( .A(KEYINPUT80), .B(KEYINPUT25), .Z(n383) );
  XNOR2_X1 U460 ( .A(n383), .B(KEYINPUT97), .ZN(n384) );
  XNOR2_X1 U461 ( .A(n385), .B(n384), .ZN(n386) );
  NAND2_X1 U462 ( .A1(G221), .A2(n388), .ZN(n389) );
  XNOR2_X1 U463 ( .A(n389), .B(KEYINPUT21), .ZN(n674) );
  XNOR2_X1 U464 ( .A(n674), .B(KEYINPUT98), .ZN(n564) );
  INV_X1 U465 ( .A(n564), .ZN(n390) );
  XNOR2_X2 U466 ( .A(KEYINPUT67), .B(G143), .ZN(n391) );
  XNOR2_X2 U467 ( .A(n391), .B(G128), .ZN(n447) );
  XNOR2_X2 U468 ( .A(n447), .B(KEYINPUT4), .ZN(n428) );
  XNOR2_X1 U469 ( .A(G134), .B(G131), .ZN(n392) );
  XNOR2_X2 U470 ( .A(n428), .B(n392), .ZN(n620) );
  XNOR2_X1 U471 ( .A(KEYINPUT94), .B(n393), .ZN(n618) );
  XNOR2_X1 U472 ( .A(G101), .B(G110), .ZN(n394) );
  XNOR2_X1 U473 ( .A(n351), .B(n394), .ZN(n431) );
  XOR2_X1 U474 ( .A(n618), .B(n431), .Z(n396) );
  NAND2_X1 U475 ( .A1(n622), .A2(G227), .ZN(n395) );
  XNOR2_X1 U476 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U477 ( .A(n413), .B(n397), .ZN(n648) );
  INV_X1 U478 ( .A(KEYINPUT70), .ZN(n398) );
  XNOR2_X1 U479 ( .A(n398), .B(G469), .ZN(n399) );
  INV_X1 U480 ( .A(n527), .ZN(n401) );
  NAND2_X1 U481 ( .A1(n356), .A2(n401), .ZN(n403) );
  INV_X1 U482 ( .A(KEYINPUT78), .ZN(n402) );
  XNOR2_X1 U483 ( .A(n403), .B(n402), .ZN(n421) );
  XNOR2_X1 U484 ( .A(G116), .B(G113), .ZN(n404) );
  XNOR2_X1 U485 ( .A(n404), .B(KEYINPUT71), .ZN(n406) );
  XOR2_X1 U486 ( .A(KEYINPUT3), .B(G119), .Z(n405) );
  XNOR2_X1 U487 ( .A(n406), .B(n405), .ZN(n432) );
  NOR2_X1 U488 ( .A1(G953), .A2(G237), .ZN(n453) );
  NAND2_X1 U489 ( .A1(n453), .A2(G210), .ZN(n408) );
  INV_X1 U490 ( .A(G137), .ZN(n407) );
  XNOR2_X1 U491 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U492 ( .A(KEYINPUT5), .B(G101), .ZN(n409) );
  XNOR2_X1 U493 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U494 ( .A(n432), .B(n411), .ZN(n412) );
  XNOR2_X1 U495 ( .A(n413), .B(n412), .ZN(n607) );
  OR2_X2 U496 ( .A1(n607), .A2(G902), .ZN(n415) );
  INV_X1 U497 ( .A(G472), .ZN(n414) );
  XNOR2_X2 U498 ( .A(n415), .B(n414), .ZN(n516) );
  INV_X1 U499 ( .A(G237), .ZN(n416) );
  NAND2_X1 U500 ( .A1(n465), .A2(n416), .ZN(n436) );
  NAND2_X1 U501 ( .A1(n436), .A2(G214), .ZN(n687) );
  INV_X1 U502 ( .A(n687), .ZN(n489) );
  INV_X1 U503 ( .A(KEYINPUT108), .ZN(n417) );
  XNOR2_X1 U504 ( .A(n417), .B(KEYINPUT30), .ZN(n418) );
  XNOR2_X1 U505 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U506 ( .A(n423), .B(KEYINPUT18), .ZN(n426) );
  XOR2_X1 U507 ( .A(n424), .B(KEYINPUT17), .Z(n425) );
  XNOR2_X1 U508 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U509 ( .A(KEYINPUT75), .B(G122), .Z(n429) );
  XNOR2_X1 U510 ( .A(n433), .B(n432), .ZN(n739) );
  XNOR2_X1 U511 ( .A(n434), .B(n739), .ZN(n656) );
  NAND2_X1 U512 ( .A1(n656), .A2(n435), .ZN(n438) );
  NAND2_X1 U513 ( .A1(n436), .A2(G210), .ZN(n437) );
  XNOR2_X2 U514 ( .A(n438), .B(n437), .ZN(n537) );
  XNOR2_X1 U515 ( .A(n537), .B(KEYINPUT38), .ZN(n471) );
  NAND2_X1 U516 ( .A1(n505), .A2(n471), .ZN(n440) );
  XNOR2_X1 U517 ( .A(KEYINPUT86), .B(KEYINPUT39), .ZN(n439) );
  XNOR2_X1 U518 ( .A(n440), .B(n439), .ZN(n539) );
  XNOR2_X1 U519 ( .A(G116), .B(G134), .ZN(n441) );
  XNOR2_X1 U520 ( .A(n441), .B(G122), .ZN(n445) );
  XOR2_X1 U521 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n443) );
  XNOR2_X1 U522 ( .A(G107), .B(KEYINPUT101), .ZN(n442) );
  XNOR2_X1 U523 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U524 ( .A(n445), .B(n444), .Z(n446) );
  XNOR2_X1 U525 ( .A(n447), .B(n446), .ZN(n450) );
  AND2_X1 U526 ( .A1(n448), .A2(G217), .ZN(n449) );
  XNOR2_X1 U527 ( .A(n450), .B(n449), .ZN(n644) );
  NAND2_X1 U528 ( .A1(n644), .A2(n465), .ZN(n452) );
  XNOR2_X1 U529 ( .A(KEYINPUT102), .B(G478), .ZN(n451) );
  XNOR2_X1 U530 ( .A(n452), .B(n451), .ZN(n502) );
  INV_X1 U531 ( .A(n502), .ZN(n486) );
  XOR2_X1 U532 ( .A(G131), .B(G140), .Z(n455) );
  NAND2_X1 U533 ( .A1(G214), .A2(n453), .ZN(n454) );
  XNOR2_X1 U534 ( .A(n455), .B(n454), .ZN(n463) );
  XOR2_X1 U535 ( .A(G122), .B(G104), .Z(n457) );
  XNOR2_X1 U536 ( .A(G113), .B(G143), .ZN(n456) );
  XNOR2_X1 U537 ( .A(n457), .B(n456), .ZN(n461) );
  XOR2_X1 U538 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n459) );
  XNOR2_X1 U539 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n458) );
  XNOR2_X1 U540 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U541 ( .A(n461), .B(n460), .Z(n462) );
  XNOR2_X1 U542 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U543 ( .A(n464), .B(n619), .ZN(n631) );
  NAND2_X1 U544 ( .A1(n631), .A2(n465), .ZN(n467) );
  XOR2_X1 U545 ( .A(KEYINPUT13), .B(G475), .Z(n466) );
  XNOR2_X1 U546 ( .A(n467), .B(n466), .ZN(n503) );
  NAND2_X1 U547 ( .A1(n486), .A2(n503), .ZN(n520) );
  INV_X1 U548 ( .A(n520), .ZN(n468) );
  NAND2_X1 U549 ( .A1(n539), .A2(n468), .ZN(n470) );
  XNOR2_X1 U550 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n469) );
  XNOR2_X2 U551 ( .A(n470), .B(n469), .ZN(n636) );
  OR2_X1 U552 ( .A1(n502), .A2(n503), .ZN(n690) );
  XNOR2_X1 U553 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n472) );
  XNOR2_X1 U554 ( .A(n473), .B(n472), .ZN(n672) );
  INV_X1 U555 ( .A(n674), .ZN(n474) );
  AND2_X1 U556 ( .A1(n475), .A2(n474), .ZN(n476) );
  INV_X1 U557 ( .A(n354), .ZN(n675) );
  NAND2_X1 U558 ( .A1(n476), .A2(n675), .ZN(n517) );
  OR2_X1 U559 ( .A1(n517), .A2(n677), .ZN(n479) );
  INV_X1 U560 ( .A(KEYINPUT28), .ZN(n478) );
  XNOR2_X1 U561 ( .A(n479), .B(n478), .ZN(n481) );
  XNOR2_X1 U562 ( .A(n527), .B(KEYINPUT109), .ZN(n480) );
  NAND2_X1 U563 ( .A1(n481), .A2(n480), .ZN(n494) );
  INV_X1 U564 ( .A(n494), .ZN(n482) );
  NAND2_X1 U565 ( .A1(n672), .A2(n482), .ZN(n483) );
  XNOR2_X1 U566 ( .A(n483), .B(KEYINPUT42), .ZN(n744) );
  XNOR2_X1 U567 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n484) );
  XNOR2_X1 U568 ( .A(n485), .B(n484), .ZN(n514) );
  INV_X1 U569 ( .A(KEYINPUT83), .ZN(n488) );
  OR2_X1 U570 ( .A1(n486), .A2(n503), .ZN(n730) );
  NAND2_X1 U571 ( .A1(n730), .A2(n520), .ZN(n592) );
  INV_X1 U572 ( .A(n592), .ZN(n693) );
  NOR2_X1 U573 ( .A1(KEYINPUT69), .A2(n693), .ZN(n497) );
  INV_X1 U574 ( .A(n497), .ZN(n487) );
  NAND2_X1 U575 ( .A1(n488), .A2(n487), .ZN(n495) );
  NOR2_X2 U576 ( .A1(n537), .A2(n489), .ZN(n491) );
  XNOR2_X1 U577 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n490) );
  XNOR2_X1 U578 ( .A(n491), .B(n490), .ZN(n554) );
  BUF_X1 U579 ( .A(n554), .Z(n492) );
  INV_X1 U580 ( .A(n492), .ZN(n493) );
  NOR2_X1 U581 ( .A1(n494), .A2(n493), .ZN(n724) );
  AND2_X1 U582 ( .A1(n495), .A2(n724), .ZN(n496) );
  NAND2_X1 U583 ( .A1(n496), .A2(KEYINPUT47), .ZN(n501) );
  NAND2_X1 U584 ( .A1(n497), .A2(n724), .ZN(n499) );
  INV_X1 U585 ( .A(KEYINPUT47), .ZN(n498) );
  NAND2_X1 U586 ( .A1(n499), .A2(n498), .ZN(n500) );
  NAND2_X1 U587 ( .A1(n501), .A2(n500), .ZN(n512) );
  NAND2_X1 U588 ( .A1(n503), .A2(n502), .ZN(n560) );
  NOR2_X1 U589 ( .A1(n537), .A2(n560), .ZN(n504) );
  AND2_X1 U590 ( .A1(n505), .A2(n504), .ZN(n722) );
  INV_X1 U591 ( .A(n722), .ZN(n508) );
  NAND2_X1 U592 ( .A1(n693), .A2(KEYINPUT47), .ZN(n506) );
  NAND2_X1 U593 ( .A1(KEYINPUT83), .A2(n506), .ZN(n507) );
  NAND2_X1 U594 ( .A1(n508), .A2(n507), .ZN(n510) );
  NAND2_X1 U595 ( .A1(n722), .A2(KEYINPUT83), .ZN(n509) );
  NAND2_X1 U596 ( .A1(n510), .A2(n509), .ZN(n511) );
  AND2_X1 U597 ( .A1(n512), .A2(n511), .ZN(n513) );
  AND2_X1 U598 ( .A1(n514), .A2(n513), .ZN(n530) );
  XNOR2_X1 U599 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n515) );
  XNOR2_X1 U600 ( .A(n516), .B(n515), .ZN(n573) );
  OR2_X2 U601 ( .A1(n573), .A2(n517), .ZN(n518) );
  XNOR2_X1 U602 ( .A(n518), .B(KEYINPUT106), .ZN(n521) );
  INV_X1 U603 ( .A(KEYINPUT104), .ZN(n519) );
  XNOR2_X1 U604 ( .A(n520), .B(n519), .ZN(n723) );
  INV_X1 U605 ( .A(n723), .ZN(n727) );
  NOR2_X2 U606 ( .A1(n521), .A2(n727), .ZN(n523) );
  XNOR2_X1 U607 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U608 ( .A1(n524), .A2(n687), .ZN(n533) );
  XNOR2_X1 U609 ( .A(n525), .B(KEYINPUT36), .ZN(n528) );
  INV_X1 U610 ( .A(KEYINPUT1), .ZN(n526) );
  NAND2_X1 U611 ( .A1(n528), .A2(n585), .ZN(n529) );
  XNOR2_X2 U612 ( .A(n529), .B(KEYINPUT112), .ZN(n637) );
  NAND2_X1 U613 ( .A1(n530), .A2(n637), .ZN(n532) );
  INV_X1 U614 ( .A(KEYINPUT48), .ZN(n531) );
  XNOR2_X1 U615 ( .A(n532), .B(n531), .ZN(n541) );
  INV_X1 U616 ( .A(n533), .ZN(n535) );
  NAND2_X1 U617 ( .A1(n535), .A2(n543), .ZN(n536) );
  XNOR2_X1 U618 ( .A(n536), .B(KEYINPUT43), .ZN(n538) );
  AND2_X1 U619 ( .A1(n538), .A2(n537), .ZN(n732) );
  INV_X1 U620 ( .A(n730), .ZN(n719) );
  AND2_X1 U621 ( .A1(n539), .A2(n719), .ZN(n615) );
  NOR2_X1 U622 ( .A1(n732), .A2(n615), .ZN(n540) );
  NAND2_X2 U623 ( .A1(n541), .A2(n540), .ZN(n602) );
  XNOR2_X2 U624 ( .A(n602), .B(KEYINPUT85), .ZN(n617) );
  OR2_X1 U625 ( .A1(n573), .A2(n542), .ZN(n544) );
  INV_X1 U626 ( .A(KEYINPUT72), .ZN(n545) );
  XNOR2_X1 U627 ( .A(n545), .B(KEYINPUT33), .ZN(n546) );
  XNOR2_X2 U628 ( .A(n547), .B(n546), .ZN(n704) );
  INV_X1 U629 ( .A(n704), .ZN(n557) );
  INV_X1 U630 ( .A(G953), .ZN(n548) );
  NOR2_X1 U631 ( .A1(n548), .A2(G898), .ZN(n549) );
  XNOR2_X1 U632 ( .A(n549), .B(KEYINPUT91), .ZN(n740) );
  NOR2_X1 U633 ( .A1(n550), .A2(n740), .ZN(n551) );
  XNOR2_X1 U634 ( .A(KEYINPUT93), .B(n551), .ZN(n553) );
  NAND2_X1 U635 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U636 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X2 U637 ( .A(n556), .B(n355), .ZN(n583) );
  NAND2_X1 U638 ( .A1(n557), .A2(n583), .ZN(n559) );
  INV_X1 U639 ( .A(KEYINPUT34), .ZN(n558) );
  XNOR2_X1 U640 ( .A(n559), .B(n558), .ZN(n562) );
  XNOR2_X1 U641 ( .A(n560), .B(KEYINPUT81), .ZN(n561) );
  NAND2_X1 U642 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U643 ( .A1(n564), .A2(n690), .ZN(n565) );
  XNOR2_X1 U644 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n566) );
  XNOR2_X2 U645 ( .A(n568), .B(n567), .ZN(n580) );
  AND2_X1 U646 ( .A1(n543), .A2(n677), .ZN(n569) );
  NAND2_X1 U647 ( .A1(n580), .A2(n569), .ZN(n571) );
  INV_X1 U648 ( .A(KEYINPUT68), .ZN(n570) );
  XNOR2_X1 U649 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n572), .A2(n675), .ZN(n629) );
  NAND2_X1 U651 ( .A1(n580), .A2(n585), .ZN(n575) );
  NAND2_X1 U652 ( .A1(n573), .A2(n675), .ZN(n574) );
  NOR2_X2 U653 ( .A1(n575), .A2(n574), .ZN(n577) );
  INV_X1 U654 ( .A(KEYINPUT32), .ZN(n576) );
  NAND2_X1 U655 ( .A1(n629), .A2(n743), .ZN(n578) );
  XNOR2_X1 U656 ( .A(n579), .B(KEYINPUT44), .ZN(n596) );
  AND2_X1 U657 ( .A1(n580), .A2(n543), .ZN(n582) );
  AND2_X1 U658 ( .A1(n573), .A2(n354), .ZN(n581) );
  NAND2_X1 U659 ( .A1(n582), .A2(n581), .ZN(n616) );
  INV_X1 U660 ( .A(n583), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n677), .A2(n542), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n682) );
  OR2_X1 U663 ( .A1(n591), .A2(n682), .ZN(n587) );
  INV_X1 U664 ( .A(KEYINPUT31), .ZN(n586) );
  XNOR2_X1 U665 ( .A(n587), .B(n586), .ZN(n729) );
  NAND2_X1 U666 ( .A1(n677), .A2(n588), .ZN(n589) );
  OR2_X1 U667 ( .A1(n589), .A2(n527), .ZN(n590) );
  OR2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n715) );
  NAND2_X1 U669 ( .A1(n729), .A2(n715), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n594) );
  AND2_X1 U671 ( .A1(n616), .A2(n594), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n598) );
  INV_X1 U673 ( .A(KEYINPUT66), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n617), .A2(n352), .ZN(n599) );
  INV_X1 U675 ( .A(KEYINPUT2), .ZN(n665) );
  NAND2_X1 U676 ( .A1(n599), .A2(n665), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n352), .A2(n603), .ZN(n605) );
  INV_X1 U678 ( .A(KEYINPUT77), .ZN(n604) );
  XNOR2_X2 U679 ( .A(n605), .B(n604), .ZN(n670) );
  NAND2_X1 U680 ( .A1(n652), .A2(G472), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n608), .B(KEYINPUT62), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n611) );
  INV_X1 U683 ( .A(n611), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n614), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U686 ( .A(G134), .B(n615), .Z(G36) );
  XNOR2_X1 U687 ( .A(n616), .B(G101), .ZN(G3) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(n621) );
  XNOR2_X1 U689 ( .A(n621), .B(n620), .ZN(n624) );
  XNOR2_X1 U690 ( .A(n663), .B(n624), .ZN(n623) );
  NAND2_X1 U691 ( .A1(n623), .A2(n622), .ZN(n628) );
  XOR2_X1 U692 ( .A(G227), .B(n624), .Z(n625) );
  NAND2_X1 U693 ( .A1(n625), .A2(G900), .ZN(n626) );
  NAND2_X1 U694 ( .A1(G953), .A2(n626), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n628), .A2(n627), .ZN(G72) );
  XNOR2_X1 U696 ( .A(n629), .B(G110), .ZN(G12) );
  XOR2_X1 U697 ( .A(G122), .B(n630), .Z(G24) );
  NAND2_X1 U698 ( .A1(n652), .A2(G475), .ZN(n633) );
  XNOR2_X1 U699 ( .A(n631), .B(KEYINPUT59), .ZN(n632) );
  XNOR2_X1 U700 ( .A(n633), .B(n632), .ZN(n634) );
  NOR2_X2 U701 ( .A1(n634), .A2(n659), .ZN(n635) );
  XNOR2_X1 U702 ( .A(n635), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U703 ( .A(n636), .B(G131), .ZN(G33) );
  XNOR2_X1 U704 ( .A(G125), .B(KEYINPUT37), .ZN(n638) );
  XOR2_X1 U705 ( .A(n638), .B(n637), .Z(G27) );
  NAND2_X1 U706 ( .A1(n646), .A2(G217), .ZN(n641) );
  XOR2_X1 U707 ( .A(KEYINPUT124), .B(n639), .Z(n640) );
  XNOR2_X1 U708 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X1 U709 ( .A1(n642), .A2(n659), .ZN(G66) );
  NAND2_X1 U710 ( .A1(n652), .A2(G478), .ZN(n643) );
  XOR2_X1 U711 ( .A(n644), .B(n643), .Z(n645) );
  NOR2_X1 U712 ( .A1(n645), .A2(n659), .ZN(G63) );
  NAND2_X1 U713 ( .A1(n646), .A2(G469), .ZN(n650) );
  XOR2_X1 U714 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n647) );
  XNOR2_X1 U715 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X1 U717 ( .A1(n651), .A2(n659), .ZN(G54) );
  NAND2_X1 U718 ( .A1(n652), .A2(G210), .ZN(n658) );
  XOR2_X1 U719 ( .A(KEYINPUT55), .B(KEYINPUT87), .Z(n654) );
  XNOR2_X1 U720 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U722 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U723 ( .A(n658), .B(n657), .ZN(n660) );
  NOR2_X2 U724 ( .A1(n660), .A2(n659), .ZN(n662) );
  XOR2_X1 U725 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n661) );
  XNOR2_X1 U726 ( .A(n662), .B(n661), .ZN(G51) );
  NOR2_X1 U727 ( .A1(n663), .A2(KEYINPUT2), .ZN(n669) );
  NAND2_X1 U728 ( .A1(n664), .A2(n665), .ZN(n667) );
  INV_X1 U729 ( .A(KEYINPUT84), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n669), .A2(n668), .ZN(n671) );
  NAND2_X1 U731 ( .A1(n671), .A2(n670), .ZN(n709) );
  NAND2_X1 U732 ( .A1(n543), .A2(n542), .ZN(n673) );
  XNOR2_X1 U733 ( .A(n673), .B(KEYINPUT50), .ZN(n681) );
  NAND2_X1 U734 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U735 ( .A(KEYINPUT49), .B(n676), .Z(n678) );
  NAND2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U737 ( .A(KEYINPUT114), .B(n679), .Z(n680) );
  NAND2_X1 U738 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U739 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U740 ( .A(KEYINPUT51), .B(n684), .Z(n685) );
  NAND2_X1 U741 ( .A1(n672), .A2(n685), .ZN(n686) );
  XNOR2_X1 U742 ( .A(n686), .B(KEYINPUT115), .ZN(n699) );
  NOR2_X1 U743 ( .A1(n471), .A2(n687), .ZN(n688) );
  XNOR2_X1 U744 ( .A(n688), .B(KEYINPUT116), .ZN(n689) );
  NOR2_X1 U745 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U746 ( .A(KEYINPUT117), .B(n691), .Z(n695) );
  NOR2_X1 U747 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U748 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U749 ( .A(KEYINPUT118), .B(n696), .ZN(n697) );
  NOR2_X1 U750 ( .A1(n697), .A2(n704), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U752 ( .A(n700), .B(KEYINPUT119), .Z(n701) );
  XNOR2_X1 U753 ( .A(KEYINPUT52), .B(n701), .ZN(n703) );
  NOR2_X1 U754 ( .A1(n703), .A2(n702), .ZN(n707) );
  INV_X1 U755 ( .A(n672), .ZN(n705) );
  NOR2_X1 U756 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U757 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U758 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U759 ( .A(n710), .B(KEYINPUT120), .ZN(n711) );
  NOR2_X1 U760 ( .A1(n711), .A2(G953), .ZN(n713) );
  XOR2_X1 U761 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n712) );
  XNOR2_X1 U762 ( .A(n713), .B(n712), .ZN(G75) );
  NOR2_X1 U763 ( .A1(n715), .A2(n727), .ZN(n714) );
  XOR2_X1 U764 ( .A(G104), .B(n714), .Z(G6) );
  NOR2_X1 U765 ( .A1(n715), .A2(n730), .ZN(n717) );
  XNOR2_X1 U766 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n716) );
  XNOR2_X1 U767 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U768 ( .A(G107), .B(n718), .ZN(G9) );
  XOR2_X1 U769 ( .A(G128), .B(KEYINPUT29), .Z(n721) );
  NAND2_X1 U770 ( .A1(n724), .A2(n719), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n721), .B(n720), .ZN(G30) );
  XOR2_X1 U772 ( .A(G143), .B(n722), .Z(G45) );
  XOR2_X1 U773 ( .A(G146), .B(KEYINPUT113), .Z(n726) );
  NAND2_X1 U774 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U775 ( .A(n726), .B(n725), .ZN(G48) );
  NOR2_X1 U776 ( .A1(n727), .A2(n729), .ZN(n728) );
  XOR2_X1 U777 ( .A(G113), .B(n728), .Z(G15) );
  NOR2_X1 U778 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U779 ( .A(G116), .B(n731), .Z(G18) );
  XOR2_X1 U780 ( .A(G140), .B(n732), .Z(G42) );
  NOR2_X1 U781 ( .A1(n664), .A2(G953), .ZN(n733) );
  XNOR2_X1 U782 ( .A(n733), .B(KEYINPUT125), .ZN(n737) );
  NAND2_X1 U783 ( .A1(G953), .A2(G224), .ZN(n734) );
  XNOR2_X1 U784 ( .A(KEYINPUT61), .B(n734), .ZN(n735) );
  NAND2_X1 U785 ( .A1(n735), .A2(G898), .ZN(n736) );
  NAND2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n738), .B(KEYINPUT126), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U789 ( .A(n742), .B(n741), .Z(G69) );
  XNOR2_X1 U790 ( .A(n743), .B(G119), .ZN(G21) );
  XOR2_X1 U791 ( .A(G137), .B(n744), .Z(n745) );
  XNOR2_X1 U792 ( .A(KEYINPUT127), .B(n745), .ZN(G39) );
endmodule

