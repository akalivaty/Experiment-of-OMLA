//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1193, new_n1194, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1240, new_n1241, new_n1242, new_n1243;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n215), .C1(G58), .C2(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G1), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n220), .B(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n223), .A2(new_n218), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT0), .Z(new_n230));
  NOR3_X1   g0030(.A1(new_n222), .A2(new_n225), .A3(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n208), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n207), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(KEYINPUT72), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n211), .A2(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n217), .A2(G13), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  NAND2_X1  g0051(.A1(new_n218), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n218), .A2(new_n254), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n248), .B1(new_n252), .B2(new_n253), .C1(new_n202), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n224), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT71), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT11), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT71), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n259), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT11), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n258), .B1(new_n217), .B2(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G68), .ZN(new_n267));
  AND4_X1   g0067(.A1(new_n251), .A2(new_n262), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT13), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  OAI211_X1 g0073(.A(G226), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(G232), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G97), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT68), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT68), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G33), .A3(G97), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n274), .A2(new_n275), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n217), .B1(G41), .B2(G45), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT65), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n282), .A2(KEYINPUT65), .A3(new_n285), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G238), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n290), .A2(KEYINPUT69), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT69), .B1(new_n290), .B2(new_n293), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n270), .B(new_n284), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n284), .B1(new_n294), .B2(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT13), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT69), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n282), .A2(KEYINPUT65), .A3(new_n285), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT65), .B1(new_n282), .B2(new_n285), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n302), .A2(new_n303), .A3(new_n212), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n301), .B1(new_n304), .B2(new_n292), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n290), .A2(KEYINPUT69), .A3(new_n293), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n307), .A2(KEYINPUT70), .A3(new_n270), .A4(new_n284), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n298), .A2(new_n300), .A3(new_n308), .A4(G179), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT75), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n270), .B1(new_n307), .B2(new_n284), .ZN(new_n311));
  INV_X1    g0111(.A(new_n284), .ZN(new_n312));
  AOI211_X1 g0112(.A(KEYINPUT13), .B(new_n312), .C1(new_n305), .C2(new_n306), .ZN(new_n313));
  OAI21_X1  g0113(.A(G169), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT14), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n269), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n298), .A2(new_n300), .A3(new_n308), .A4(G190), .ZN(new_n317));
  OAI21_X1  g0117(.A(G200), .B1(new_n311), .B2(new_n313), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(new_n268), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT73), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n317), .A2(new_n318), .A3(new_n268), .A4(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n320), .A2(KEYINPUT74), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT74), .B1(new_n320), .B2(new_n322), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n302), .A2(new_n303), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G226), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n272), .A2(new_n273), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(G1698), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(G222), .B1(G77), .B2(new_n328), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT3), .B(G33), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G223), .A3(G1698), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n293), .B(new_n327), .C1(new_n333), .C2(new_n282), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(G200), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT67), .A2(KEYINPUT9), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n226), .A2(new_n218), .A3(G1), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n202), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n266), .A2(G50), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT8), .B(G58), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n342), .A2(new_n252), .B1(new_n343), .B2(new_n255), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(G20), .B2(new_n203), .ZN(new_n345));
  INV_X1    g0145(.A(new_n258), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n340), .B(new_n341), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(KEYINPUT67), .A2(KEYINPUT9), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n338), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OR3_X1    g0149(.A1(new_n347), .A2(new_n338), .A3(new_n348), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n336), .A2(new_n337), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT10), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT7), .B1(new_n328), .B2(new_n218), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NOR4_X1   g0154(.A1(new_n272), .A2(new_n273), .A3(new_n354), .A4(G20), .ZN(new_n355));
  OAI21_X1  g0155(.A(G68), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT76), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G58), .A2(G68), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT77), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G58), .B2(G68), .ZN(new_n361));
  INV_X1    g0161(.A(new_n255), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n361), .A2(G20), .B1(G159), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(KEYINPUT76), .B(G68), .C1(new_n353), .C2(new_n355), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n358), .A2(new_n363), .A3(KEYINPUT16), .A4(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT77), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n359), .B(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n201), .ZN(new_n369));
  INV_X1    g0169(.A(G159), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n369), .A2(new_n218), .B1(new_n370), .B2(new_n255), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n354), .B1(new_n331), .B2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n328), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n211), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n366), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n365), .A2(new_n258), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n339), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n342), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n266), .B2(new_n342), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(G226), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n381));
  OAI211_X1 g0181(.A(G223), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n382));
  INV_X1    g0182(.A(G87), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n381), .B(new_n382), .C1(new_n254), .C2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n292), .B1(new_n384), .B2(new_n283), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n282), .A2(G232), .A3(new_n285), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n385), .A2(G179), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G169), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n385), .B2(new_n386), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n380), .A2(KEYINPUT18), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT18), .B1(new_n380), .B2(new_n391), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n385), .A2(new_n335), .A3(new_n386), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n384), .A2(new_n283), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n397), .A2(new_n293), .A3(new_n386), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n398), .B2(G200), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n376), .A2(new_n399), .A3(new_n379), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT17), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n352), .A2(new_n395), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n334), .A2(new_n388), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(new_n347), .C1(G179), .C2(new_n334), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT66), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n331), .A2(G232), .A3(new_n271), .ZN(new_n407));
  INV_X1    g0207(.A(G107), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n331), .A2(G1698), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n407), .B1(new_n408), .B2(new_n331), .C1(new_n409), .C2(new_n212), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n283), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n326), .A2(G244), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n293), .A3(new_n412), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n413), .A2(G179), .ZN(new_n414));
  INV_X1    g0214(.A(new_n342), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n362), .B1(G20), .B2(G77), .ZN(new_n416));
  XOR2_X1   g0216(.A(KEYINPUT15), .B(G87), .Z(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n218), .A3(G33), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n346), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n377), .A2(G77), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n266), .A2(G77), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n413), .A2(new_n388), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n414), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n413), .A2(G200), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(new_n422), .C1(new_n335), .C2(new_n413), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n406), .A2(new_n428), .ZN(new_n429));
  AND4_X1   g0229(.A1(new_n316), .A2(new_n325), .A3(new_n403), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G283), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(new_n218), .C1(G33), .C2(new_n213), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n207), .A2(G20), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n258), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT20), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n433), .A2(KEYINPUT20), .A3(new_n258), .A4(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n249), .A2(new_n434), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n254), .A2(G1), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n339), .A2(new_n258), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n442), .B2(G116), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n388), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(G264), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n331), .A2(KEYINPUT80), .A3(G264), .A4(G1698), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n329), .A2(G257), .B1(G303), .B2(new_n328), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n282), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  INV_X1    g0252(.A(G41), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT5), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(KEYINPUT78), .B2(G41), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n454), .A2(new_n456), .A3(new_n458), .A4(G274), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT79), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n454), .A2(new_n456), .A3(new_n458), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n461), .A2(new_n282), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G270), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n444), .B1(new_n451), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT21), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n447), .A2(new_n448), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n331), .A2(new_n271), .ZN(new_n469));
  INV_X1    g0269(.A(G303), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n469), .A2(new_n214), .B1(new_n470), .B2(new_n331), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n283), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n473), .A2(new_n474), .B1(new_n462), .B2(G270), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n439), .A2(new_n443), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n472), .A2(new_n475), .A3(new_n476), .A4(G179), .ZN(new_n477));
  OAI211_X1 g0277(.A(KEYINPUT21), .B(new_n444), .C1(new_n451), .C2(new_n464), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n467), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n331), .A2(new_n218), .A3(G68), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT19), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n252), .B2(new_n213), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n277), .A2(new_n279), .ZN(new_n483));
  AOI21_X1  g0283(.A(G20), .B1(new_n483), .B2(KEYINPUT19), .ZN(new_n484));
  NOR3_X1   g0284(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n480), .B(new_n482), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n417), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n486), .A2(new_n258), .B1(new_n339), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n442), .A2(new_n417), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(G238), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n491));
  OAI211_X1 g0291(.A(G244), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n491), .B(new_n492), .C1(new_n254), .C2(new_n207), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n283), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n217), .A2(G45), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n291), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n282), .A2(G250), .A3(new_n495), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n388), .ZN(new_n500));
  INV_X1    g0300(.A(new_n498), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n496), .B(new_n501), .C1(new_n493), .C2(new_n283), .ZN(new_n502));
  INV_X1    g0302(.A(G179), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n490), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(G190), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n499), .A2(G200), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n442), .A2(G87), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n488), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n475), .A2(new_n472), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n335), .ZN(new_n512));
  INV_X1    g0312(.A(G200), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n475), .B2(new_n472), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n512), .A2(new_n476), .A3(new_n514), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n479), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT24), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT22), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n218), .B(G87), .C1(new_n272), .C2(new_n273), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(KEYINPUT82), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT82), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n521), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT82), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n519), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(new_n522), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n408), .A2(KEYINPUT23), .A3(G20), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT23), .B1(new_n408), .B2(G20), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n532), .A2(new_n533), .B1(new_n207), .B2(new_n252), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n517), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  AOI211_X1 g0336(.A(KEYINPUT24), .B(new_n534), .C1(new_n525), .C2(new_n530), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n258), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n339), .A2(new_n408), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n539), .B(KEYINPUT25), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(G107), .B2(new_n442), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n331), .A2(G250), .A3(new_n271), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n409), .C2(new_n214), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n283), .B1(new_n462), .B2(G264), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n460), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n513), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n283), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n462), .A2(G264), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n548), .A2(new_n335), .A3(new_n460), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT83), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT83), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n545), .A2(new_n552), .A3(new_n335), .A4(new_n460), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n547), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n538), .A2(new_n541), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G244), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n331), .A2(G250), .A3(G1698), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n432), .B1(new_n556), .B2(new_n557), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n283), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n462), .A2(G257), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n460), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n377), .A2(G97), .ZN(new_n566));
  OAI21_X1  g0366(.A(G107), .B1(new_n353), .B2(new_n355), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n362), .A2(G77), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n213), .A2(new_n408), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n408), .A2(KEYINPUT6), .A3(G97), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n567), .B(new_n568), .C1(new_n218), .C2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n566), .B1(new_n575), .B2(new_n258), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n442), .A2(G97), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n562), .A2(G190), .A3(new_n460), .A4(new_n563), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n565), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n566), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n408), .B1(new_n372), .B2(new_n373), .ZN(new_n581));
  INV_X1    g0381(.A(new_n568), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n218), .B1(new_n572), .B2(new_n573), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n580), .B(new_n577), .C1(new_n584), .C2(new_n346), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n564), .A2(new_n388), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n562), .A2(new_n503), .A3(new_n460), .A4(new_n563), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n546), .A2(new_n388), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n545), .A2(new_n503), .A3(new_n460), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n523), .A2(new_n524), .A3(new_n519), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n529), .B1(new_n528), .B2(new_n522), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n535), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT24), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n531), .A2(new_n517), .A3(new_n535), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n346), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n541), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n593), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n516), .A2(new_n555), .A3(new_n589), .A4(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n431), .A2(new_n602), .ZN(G372));
  NAND2_X1  g0403(.A1(new_n320), .A2(new_n322), .ZN(new_n604));
  INV_X1    g0404(.A(new_n425), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n606), .A2(new_n316), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT17), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n400), .B(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n395), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n406), .B1(new_n610), .B2(new_n352), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n478), .A2(new_n477), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT21), .B1(new_n511), .B2(new_n444), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n467), .A2(KEYINPUT85), .A3(new_n477), .A4(new_n478), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n592), .B1(new_n538), .B2(new_n541), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n612), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT84), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n502), .B2(new_n513), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n499), .A2(KEYINPUT84), .A3(G200), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n506), .A2(new_n488), .A3(new_n508), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n488), .A2(new_n489), .B1(new_n388), .B2(new_n499), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(new_n504), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n555), .A2(new_n589), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n601), .A2(KEYINPUT86), .A3(new_n616), .A4(new_n617), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n620), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT87), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n588), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n488), .A2(new_n508), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n506), .A3(new_n622), .A4(new_n623), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n633), .A2(new_n635), .A3(new_n636), .A4(new_n505), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT26), .B1(new_n510), .B2(new_n588), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n505), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT88), .A4(new_n505), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n620), .A2(new_n628), .A3(new_n629), .A4(KEYINPUT87), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n632), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n611), .B1(new_n431), .B2(new_n646), .ZN(G369));
  NOR2_X1   g0447(.A1(new_n226), .A2(G20), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n217), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n476), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n616), .B2(new_n617), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n479), .A2(new_n515), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT89), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n654), .B1(new_n599), .B2(new_n600), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n619), .B1(new_n662), .B2(new_n555), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n601), .A2(new_n654), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n479), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n654), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(G399));
  NOR2_X1   g0470(.A1(new_n227), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n485), .A2(new_n207), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n223), .B2(new_n672), .ZN(new_n676));
  XOR2_X1   g0476(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n677));
  XNOR2_X1  g0477(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  INV_X1    g0479(.A(new_n654), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n645), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n622), .A2(new_n623), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n506), .A2(new_n488), .A3(new_n508), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n505), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT26), .B1(new_n684), .B2(new_n588), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n633), .A2(new_n636), .A3(new_n509), .A4(new_n505), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n505), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT92), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n601), .A2(new_n667), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n628), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT92), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n685), .A2(new_n686), .A3(new_n691), .A4(new_n505), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n680), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n681), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n511), .A2(new_n503), .ZN(new_n697));
  INV_X1    g0497(.A(new_n564), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n545), .A3(new_n698), .A4(new_n502), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT91), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT30), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n511), .A2(new_n564), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n703), .A2(new_n503), .A3(new_n546), .A4(new_n499), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n699), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n654), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT31), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n708), .B(KEYINPUT31), .C1(new_n602), .C2(new_n654), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n696), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n678), .B1(new_n714), .B2(G1), .ZN(G364));
  NOR2_X1   g0515(.A1(G13), .A2(G33), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n658), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n217), .B1(new_n648), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n671), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n224), .B1(G20), .B2(new_n388), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n242), .A2(G45), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n227), .A2(new_n331), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n726), .B(new_n727), .C1(G45), .C2(new_n223), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n228), .A2(G355), .A3(new_n331), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G116), .B2(new_n228), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT93), .Z(new_n731));
  AOI21_X1  g0531(.A(new_n725), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n335), .A2(G20), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT96), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n735), .A2(G179), .A3(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G159), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT32), .Z(new_n738));
  NOR2_X1   g0538(.A1(new_n513), .A2(G179), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n408), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n218), .A2(new_n335), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n745), .A2(new_n503), .A3(G200), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G58), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n331), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n745), .A2(new_n740), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n383), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n218), .A2(new_n503), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(new_n335), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n218), .B1(new_n755), .B2(G190), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n754), .A2(new_n211), .B1(new_n756), .B2(new_n213), .ZN(new_n757));
  NOR4_X1   g0557(.A1(new_n743), .A2(new_n749), .A3(new_n752), .A4(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n335), .A2(new_n513), .A3(G20), .A4(G179), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G77), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n753), .A2(G190), .A3(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT95), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n765), .A2(KEYINPUT95), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G50), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n738), .A2(new_n758), .A3(new_n764), .A4(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n331), .B1(new_n746), .B2(G322), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT33), .B(G317), .Z(new_n774));
  OAI221_X1 g0574(.A(new_n773), .B1(new_n470), .B2(new_n751), .C1(new_n754), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G326), .B2(new_n770), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n736), .A2(G329), .B1(new_n741), .B2(G283), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n762), .ZN(new_n779));
  INV_X1    g0579(.A(G294), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n756), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n772), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n732), .B1(new_n782), .B2(new_n723), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n719), .A2(new_n722), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n722), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n660), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n659), .A2(G330), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(G396));
  INV_X1    g0588(.A(new_n713), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n423), .A2(new_n654), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n425), .A2(new_n427), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT100), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n645), .A2(new_n680), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n793), .B1(new_n425), .B2(new_n680), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n645), .B2(new_n680), .ZN(new_n798));
  OR3_X1    g0598(.A1(new_n789), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n789), .B1(new_n796), .B2(new_n798), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n799), .A2(new_n785), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n723), .A2(new_n716), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n785), .B1(new_n253), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT97), .ZN(new_n804));
  INV_X1    g0604(.A(new_n756), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n328), .B1(new_n805), .B2(G58), .ZN(new_n806));
  INV_X1    g0606(.A(new_n736), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n742), .B2(new_n211), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n754), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n763), .A2(G159), .B1(G150), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  INV_X1    g0612(.A(G143), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(new_n812), .B2(new_n769), .C1(new_n813), .C2(new_n747), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT34), .Z(new_n815));
  AOI211_X1 g0615(.A(new_n809), .B(new_n815), .C1(G50), .C2(new_n750), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n751), .A2(new_n408), .B1(new_n756), .B2(new_n213), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n331), .B(new_n817), .C1(G294), .C2(new_n746), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n818), .B1(new_n470), .B2(new_n769), .C1(new_n778), .C2(new_n807), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n762), .A2(new_n207), .B1(new_n820), .B2(new_n754), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT98), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n742), .A2(new_n383), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n819), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT99), .Z(new_n826));
  INV_X1    g0626(.A(new_n723), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n804), .B1(new_n717), .B2(new_n797), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n801), .A2(new_n828), .ZN(G384));
  INV_X1    g0629(.A(KEYINPUT35), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n218), .B(new_n224), .C1(new_n574), .C2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n831), .B(G116), .C1(new_n830), .C2(new_n574), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT36), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n368), .A2(new_n253), .A3(new_n223), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT101), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n211), .A2(G50), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n226), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n217), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT102), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n605), .A2(new_n680), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n795), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  INV_X1    g0642(.A(new_n652), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n380), .B1(new_n391), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT37), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n844), .A2(new_n845), .A3(new_n400), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n358), .A2(new_n363), .A3(new_n364), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n366), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n258), .A3(new_n365), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n849), .A2(new_n379), .B1(new_n390), .B2(new_n652), .ZN(new_n850));
  INV_X1    g0650(.A(new_n400), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT37), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n401), .B1(new_n393), .B2(new_n392), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n652), .B1(new_n849), .B2(new_n379), .ZN(new_n854));
  AOI221_X4 g0654(.A(new_n842), .B1(new_n846), .B2(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n852), .A2(new_n846), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT38), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n310), .A2(new_n315), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n323), .B2(new_n324), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n269), .A2(new_n654), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n320), .B2(new_n322), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n316), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n841), .A2(new_n859), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n395), .A2(new_n843), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT103), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n652), .B1(new_n376), .B2(new_n379), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n394), .B2(new_n609), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n390), .A2(new_n652), .B1(new_n376), .B2(new_n379), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n875), .A2(new_n851), .A3(KEYINPUT37), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n845), .B1(new_n844), .B2(new_n400), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT105), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n875), .B2(new_n851), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT105), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n846), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n874), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n856), .A2(KEYINPUT38), .A3(new_n857), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT39), .B1(new_n855), .B2(new_n858), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT106), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n884), .A2(new_n890), .A3(new_n885), .A4(new_n886), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n316), .A2(new_n654), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n868), .A2(new_n895), .A3(new_n870), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n872), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n696), .A2(new_n430), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n611), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n709), .A2(new_n710), .A3(new_n797), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n867), .A2(new_n859), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n884), .A2(new_n886), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n867), .A2(KEYINPUT40), .A3(new_n901), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n431), .A2(new_n711), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n907), .B(new_n908), .Z(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(new_n712), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n900), .B(new_n910), .Z(new_n911));
  NOR2_X1   g0711(.A1(new_n648), .A2(new_n217), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n839), .B1(new_n911), .B2(new_n912), .ZN(G367));
  INV_X1    g0713(.A(new_n727), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n238), .A2(new_n914), .B1(new_n228), .B2(new_n487), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n722), .B1(new_n915), .B2(new_n725), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT111), .ZN(new_n917));
  INV_X1    g0717(.A(new_n718), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n634), .A2(new_n680), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n626), .A3(new_n504), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n684), .B2(new_n919), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n810), .A2(G159), .B1(new_n805), .B2(G68), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n328), .B1(new_n750), .B2(G58), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(new_n769), .C2(new_n813), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n741), .A2(G77), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n925), .B1(new_n202), .B2(new_n762), .C1(new_n807), .C2(new_n812), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n924), .B(new_n926), .C1(G150), .C2(new_n746), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n331), .B1(new_n805), .B2(G107), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n928), .B1(new_n780), .B2(new_n754), .C1(new_n769), .C2(new_n778), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n750), .A2(G116), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT46), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n763), .A2(G283), .B1(new_n741), .B2(G97), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n736), .A2(G317), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n929), .B(new_n934), .C1(G303), .C2(new_n746), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT47), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n917), .B1(new_n918), .B2(new_n921), .C1(new_n937), .C2(new_n827), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n665), .A2(new_n668), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n585), .A2(new_n654), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n589), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT42), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n669), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT42), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n664), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n942), .B1(new_n588), .B2(new_n654), .C1(new_n945), .C2(new_n941), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT107), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n633), .A2(new_n654), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n941), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n666), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n952), .B(new_n953), .C1(KEYINPUT108), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(KEYINPUT108), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n943), .A2(new_n956), .B1(KEYINPUT109), .B2(KEYINPUT44), .ZN(new_n961));
  NOR2_X1   g0761(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT110), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n669), .A2(new_n955), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT45), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n661), .A3(new_n665), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n964), .A2(new_n666), .A3(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n665), .B(new_n668), .Z(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(new_n660), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n714), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n714), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n671), .B(KEYINPUT41), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n721), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n938), .B1(new_n960), .B2(new_n977), .ZN(G387));
  OR2_X1    g0778(.A1(new_n972), .A2(new_n714), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(new_n671), .A3(new_n973), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n972), .A2(new_n721), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n342), .A2(KEYINPUT50), .A3(G50), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n673), .B1(G68), .B2(G77), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT50), .B1(new_n342), .B2(G50), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n457), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n914), .B1(new_n235), .B2(G45), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n674), .A2(new_n227), .A3(new_n328), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n227), .A2(new_n408), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n725), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n736), .A2(G326), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n763), .A2(G303), .B1(G317), .B2(new_n746), .ZN(new_n992));
  INV_X1    g0792(.A(G322), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n778), .B2(new_n754), .C1(new_n993), .C2(new_n769), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT48), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n820), .B2(new_n756), .C1(new_n780), .C2(new_n751), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT49), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n331), .B(new_n991), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n997), .B2(new_n996), .C1(new_n207), .C2(new_n742), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n751), .A2(new_n253), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n342), .B2(new_n754), .C1(new_n487), .C2(new_n756), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n331), .B1(new_n202), .B2(new_n747), .C1(new_n769), .C2(new_n370), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n742), .A2(new_n213), .B1(new_n211), .B2(new_n762), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n343), .B2(new_n807), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n990), .B1(new_n1007), .B2(new_n723), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n722), .C1(new_n665), .C2(new_n918), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n980), .A2(new_n981), .A3(new_n1009), .ZN(G393));
  AOI21_X1  g0810(.A(new_n672), .B1(new_n970), .B2(new_n973), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n974), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n970), .A2(KEYINPUT112), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT112), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n968), .B2(new_n969), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n721), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n770), .A2(G317), .B1(G311), .B2(new_n746), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT114), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT52), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n331), .B1(new_n810), .B2(G303), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n207), .B2(new_n756), .C1(new_n820), .C2(new_n751), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n743), .B(new_n1021), .C1(G322), .C2(new_n736), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1019), .B(new_n1022), .C1(new_n780), .C2(new_n762), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n742), .A2(new_n383), .B1(new_n342), .B2(new_n762), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n756), .A2(new_n253), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G50), .B2(new_n810), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1026), .B(new_n331), .C1(new_n211), .C2(new_n751), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n769), .A2(new_n343), .B1(new_n370), .B2(new_n747), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT51), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1024), .B(new_n1027), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n1029), .B2(new_n1028), .C1(new_n813), .C2(new_n807), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1023), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n785), .B1(new_n1032), .B2(new_n723), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n724), .B1(new_n213), .B2(new_n228), .C1(new_n245), .C2(new_n914), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT113), .Z(new_n1035));
  OAI211_X1 g0835(.A(new_n1033), .B(new_n1035), .C1(new_n918), .C2(new_n955), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1012), .A2(new_n1016), .A3(new_n1036), .ZN(G390));
  AOI22_X1  g0837(.A1(new_n861), .A2(new_n863), .B1(new_n316), .B2(new_n865), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n709), .A2(new_n710), .A3(G330), .A4(new_n797), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n893), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n841), .A2(new_n867), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n892), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n905), .A2(new_n1041), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n693), .A2(new_n680), .A3(new_n794), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT115), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n1046), .A3(new_n840), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1046), .B1(new_n1045), .B2(new_n840), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1044), .B1(new_n1050), .B2(new_n867), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1040), .B1(new_n1043), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1045), .A2(new_n840), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT115), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n867), .A3(new_n1047), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n1041), .A3(new_n905), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1039), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n867), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1038), .B1(new_n795), .B2(new_n840), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1059), .A2(new_n893), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1056), .B(new_n1058), .C1(new_n892), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1052), .A2(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n325), .A2(new_n429), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n711), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n403), .A2(new_n316), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1063), .A2(G330), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n898), .A2(new_n611), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n841), .B1(new_n1069), .B2(new_n1040), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1058), .B(new_n1068), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1067), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1072), .A2(KEYINPUT116), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(KEYINPUT116), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1062), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1052), .A2(new_n1061), .A3(new_n1072), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n671), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1052), .A2(new_n721), .A3(new_n1061), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT54), .B(G143), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n762), .A2(new_n1079), .B1(new_n812), .B2(new_n754), .ZN(new_n1080));
  OR3_X1    g0880(.A1(new_n751), .A2(KEYINPUT53), .A3(new_n343), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT53), .B1(new_n751), .B2(new_n343), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(new_n370), .C2(new_n756), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1080), .B(new_n1083), .C1(G128), .C2(new_n770), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n328), .B1(new_n736), .B2(G125), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n202), .B2(new_n742), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT117), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1084), .B(new_n1087), .C1(new_n808), .C2(new_n747), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n770), .A2(G283), .B1(G97), .B2(new_n763), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n408), .B2(new_n754), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT118), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n807), .A2(new_n780), .B1(new_n742), .B2(new_n211), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(new_n1025), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n331), .B(new_n752), .C1(G116), .C2(new_n746), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1092), .A2(new_n1093), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n827), .B1(new_n1088), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n342), .B2(new_n802), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n722), .B(new_n1099), .C1(new_n892), .C2(new_n717), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1077), .A2(new_n1078), .A3(new_n1100), .ZN(G378));
  AOI211_X1 g0901(.A(KEYINPUT103), .B(new_n869), .C1(new_n1059), .C2(new_n859), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n895), .B1(new_n868), .B2(new_n870), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT56), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n352), .A2(new_n405), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n347), .A3(new_n843), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT55), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n347), .A2(new_n843), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n352), .A2(new_n405), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1108), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1105), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1113), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n1111), .A3(KEYINPUT56), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1117), .A2(new_n904), .A3(G330), .A4(new_n906), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n855), .A2(new_n858), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n709), .A2(new_n710), .A3(new_n797), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1038), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(G330), .B(new_n906), .C1(new_n1121), .C2(KEYINPUT40), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1104), .A2(new_n894), .A3(new_n1118), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1118), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n897), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1067), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1076), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1128), .A2(new_n1130), .A3(KEYINPUT57), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n671), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1123), .A2(new_n716), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n802), .A2(new_n202), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n453), .B(new_n328), .C1(new_n747), .C2(new_n408), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1001), .B1(new_n211), .B2(new_n756), .C1(new_n213), .C2(new_n754), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(G116), .C2(new_n770), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n763), .A2(new_n417), .B1(new_n741), .B2(G58), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n820), .C2(new_n807), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT58), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n202), .B1(new_n272), .B2(G41), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n762), .A2(new_n812), .B1(new_n808), .B2(new_n754), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n746), .A2(G128), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n751), .A2(new_n1079), .B1(new_n343), .B2(new_n756), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n770), .B2(G125), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT59), .Z(new_n1151));
  AOI21_X1  g0951(.A(G41), .B1(new_n736), .B2(G124), .ZN(new_n1152));
  AOI21_X1  g0952(.A(G33), .B1(new_n741), .B2(G159), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1143), .A2(new_n1144), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n785), .B1(new_n1155), .B2(new_n723), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1136), .A2(new_n1137), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n1128), .B2(new_n721), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1135), .A2(new_n1159), .ZN(G375));
  NAND3_X1  g0960(.A1(new_n1067), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n976), .B(new_n1161), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT120), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n720), .B(KEYINPUT121), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G128), .A2(new_n736), .B1(new_n763), .B2(G150), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n756), .A2(new_n202), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n754), .A2(new_n1079), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(G137), .C2(new_n746), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1167), .B(new_n1170), .C1(new_n808), .C2(new_n769), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n328), .B1(new_n741), .B2(G58), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT123), .Z(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G159), .C2(new_n750), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n810), .A2(G116), .B1(new_n805), .B2(new_n417), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n331), .B1(new_n746), .B2(G283), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n769), .C2(new_n780), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n925), .B1(new_n408), .B2(new_n762), .C1(new_n807), .C2(new_n470), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(G97), .C2(new_n750), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1174), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1180), .A2(new_n827), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1038), .B2(new_n716), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n785), .B1(new_n211), .B2(new_n802), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT122), .Z(new_n1184));
  AOI21_X1  g0984(.A(new_n1166), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT124), .Z(new_n1186));
  NAND2_X1  g0986(.A1(new_n1163), .A2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT125), .Z(G381));
  NOR3_X1   g0988(.A1(G381), .A2(G384), .A3(G387), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(G375), .A2(G378), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(G407));
  INV_X1    g0992(.A(G213), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1190), .B2(new_n653), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(G407), .A2(new_n1194), .ZN(G409));
  NOR2_X1   g0995(.A1(new_n1193), .A2(G343), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1135), .A2(G378), .A3(new_n1159), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT126), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT126), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1135), .A2(G378), .A3(new_n1199), .A4(new_n1159), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1130), .A2(new_n976), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1128), .B1(new_n1202), .B2(new_n1164), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G378), .B1(new_n1157), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1196), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT127), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1161), .A2(new_n1207), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n672), .B(new_n1072), .C1(new_n1208), .C2(KEYINPUT60), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(KEYINPUT60), .B2(new_n1208), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1186), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(new_n801), .A3(new_n828), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1186), .A2(new_n1210), .A3(G384), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1196), .A2(G2897), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1214), .B(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT63), .B1(new_n1206), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1214), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1206), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT61), .ZN(new_n1221));
  XOR2_X1   g1021(.A(G393), .B(G396), .Z(new_n1222));
  AND2_X1   g1022(.A1(G390), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G390), .A2(new_n1222), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n938), .C1(new_n977), .C2(new_n960), .ZN(new_n1226));
  OAI21_X1  g1026(.A(G387), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1204), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1229), .A2(new_n1196), .A3(new_n1214), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1228), .B1(new_n1230), .B2(KEYINPUT63), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1220), .A2(new_n1221), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1221), .B1(new_n1206), .B2(new_n1216), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT62), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1206), .B2(new_n1218), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1229), .A2(KEYINPUT62), .A3(new_n1196), .A4(new_n1214), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1233), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1228), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1232), .B1(new_n1237), .B2(new_n1238), .ZN(G405));
  INV_X1    g1039(.A(G378), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G375), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1201), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(new_n1218), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(new_n1228), .ZN(G402));
endmodule


