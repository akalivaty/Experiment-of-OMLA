//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n638, new_n639,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G235), .A3(G237), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(G2106), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT69), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT69), .B1(new_n465), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n464), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(KEYINPUT70), .A3(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n472), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n482), .B(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G101), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n483), .A2(KEYINPUT3), .A3(new_n484), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n494), .A2(new_n462), .A3(G137), .A4(new_n465), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G101), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT72), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n499), .B2(new_n490), .ZN(new_n500));
  INV_X1    g075(.A(new_n495), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT73), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n463), .A2(new_n481), .B1(new_n496), .B2(new_n502), .ZN(G160));
  AND2_X1   g078(.A1(new_n494), .A2(new_n465), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n486), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT74), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n504), .A2(new_n507), .A3(new_n486), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G136), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT75), .ZN(new_n511));
  OAI221_X1 g086(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n462), .C2(G112), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n504), .A2(new_n463), .ZN(new_n513));
  INV_X1    g088(.A(G124), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n511), .A2(new_n515), .ZN(G162));
  NOR2_X1   g091(.A1(new_n468), .A2(new_n469), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(G138), .A3(new_n462), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT77), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n494), .A2(new_n462), .A3(G138), .A4(new_n465), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT4), .ZN(new_n522));
  INV_X1    g097(.A(new_n461), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G138), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT77), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n478), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n520), .A2(new_n522), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n531));
  INV_X1    g106(.A(G114), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n531), .B1(new_n532), .B2(G2105), .ZN(new_n533));
  AND2_X1   g108(.A1(G126), .A2(G2105), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n533), .B1(new_n504), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(G164));
  XNOR2_X1  g112(.A(KEYINPUT5), .B(G543), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT6), .B(G651), .Z(new_n540));
  OAI21_X1  g115(.A(KEYINPUT78), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n538), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g119(.A1(new_n539), .A2(KEYINPUT78), .A3(new_n540), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(G303));
  INV_X1    g121(.A(G303), .ZN(G166));
  INV_X1    g122(.A(KEYINPUT80), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT6), .B(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT80), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n549), .A2(G543), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G51), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n538), .B(KEYINPUT79), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n555), .A2(G63), .A3(G651), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n538), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n540), .ZN(new_n559));
  NAND3_X1  g134(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT7), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n560), .A2(KEYINPUT7), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n559), .A2(G89), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n554), .B1(new_n553), .B2(new_n556), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT82), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n553), .A2(new_n556), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT81), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n568), .A2(new_n569), .A3(new_n557), .A4(new_n563), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G168));
  NAND2_X1  g146(.A1(new_n552), .A2(G52), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n559), .A2(G90), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n555), .A2(G64), .ZN(new_n575));
  NAND2_X1  g150(.A1(G77), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n542), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(G171));
  NAND2_X1  g153(.A1(G68), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n538), .B(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G56), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT83), .B(G81), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n552), .A2(G43), .B1(new_n559), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G860), .ZN(G153));
  AND3_X1   g164(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G36), .ZN(G176));
  NAND2_X1  g166(.A1(G1), .A2(G3), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT8), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(G188));
  NAND4_X1  g169(.A1(new_n549), .A2(G53), .A3(G543), .A4(new_n551), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT9), .ZN(new_n596));
  NAND2_X1  g171(.A1(G78), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G65), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n558), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(new_n559), .B2(G91), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(G299));
  INV_X1    g176(.A(G171), .ZN(G301));
  INV_X1    g177(.A(G168), .ZN(G286));
  OAI21_X1  g178(.A(G651), .B1(new_n555), .B2(G74), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT84), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n552), .A2(G49), .B1(G87), .B2(new_n559), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n607), .B(G651), .C1(new_n555), .C2(G74), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(G288));
  AOI22_X1  g184(.A1(new_n538), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(new_n542), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n538), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(new_n540), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT85), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(G305));
  NAND2_X1  g191(.A1(G72), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G60), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n581), .B2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n542), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(new_n619), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n552), .A2(G47), .B1(G85), .B2(new_n559), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(G290));
  AOI22_X1  g199(.A1(new_n538), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n625), .A2(new_n542), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(new_n552), .B2(G54), .ZN(new_n627));
  AND3_X1   g202(.A1(new_n550), .A2(new_n538), .A3(G92), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT10), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G171), .B2(new_n631), .ZN(G284));
  OAI21_X1  g208(.A(new_n632), .B1(G171), .B2(new_n631), .ZN(G321));
  NOR2_X1   g209(.A1(G299), .A2(G868), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g211(.A(new_n635), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g212(.A(new_n630), .ZN(new_n638));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n638), .B1(new_n639), .B2(G860), .ZN(G148));
  NAND2_X1  g215(.A1(new_n587), .A2(new_n631), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n630), .A2(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(new_n631), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g219(.A1(new_n509), .A2(G135), .ZN(new_n645));
  OAI221_X1 g220(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n462), .C2(G111), .ZN(new_n646));
  INV_X1    g221(.A(G123), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n513), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(G2096), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(G2096), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n499), .A2(new_n490), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(new_n478), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT12), .Z(new_n655));
  XOR2_X1   g230(.A(KEYINPUT87), .B(KEYINPUT13), .Z(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n652), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(G156));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT14), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2451), .B(G2454), .Z(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G14), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(G401));
  INV_X1    g252(.A(KEYINPUT18), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(KEYINPUT17), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n681), .B2(KEYINPUT18), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT90), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2096), .B(G2100), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT19), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  OR3_X1    g275(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n696), .A2(new_n700), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n696), .A2(new_n699), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT20), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G1981), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(G1981), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n693), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n709), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n711), .A2(new_n707), .A3(G1986), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n710), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n715), .B1(new_n710), .B2(new_n712), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n692), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n710), .A2(new_n712), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(new_n714), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n721), .A2(new_n716), .A3(new_n691), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n722), .ZN(G229));
  XNOR2_X1  g298(.A(KEYINPUT94), .B(KEYINPUT36), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n615), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G6), .B2(G16), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT32), .B(G1981), .Z(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n726), .B(new_n728), .C1(G6), .C2(G16), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G22), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G166), .B2(new_n732), .ZN(new_n734));
  INV_X1    g309(.A(G1971), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(G1971), .B(new_n733), .C1(G166), .C2(new_n732), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n730), .A2(new_n731), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n732), .A2(G23), .ZN(new_n739));
  INV_X1    g314(.A(G288), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n732), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT33), .B(G1976), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n725), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT93), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G290), .A2(new_n732), .ZN(new_n747));
  NOR2_X1   g322(.A1(G16), .A2(G24), .ZN(new_n748));
  OR3_X1    g323(.A1(new_n747), .A2(new_n693), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G25), .ZN(new_n751));
  OAI221_X1 g326(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n462), .C2(G107), .ZN(new_n752));
  INV_X1    g327(.A(G119), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n513), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n509), .B2(G131), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n751), .B1(new_n755), .B2(new_n750), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT35), .B(G1991), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n756), .B(new_n757), .Z(new_n758));
  OAI21_X1  g333(.A(new_n693), .B1(new_n747), .B2(new_n748), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n749), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n738), .A2(new_n725), .A3(new_n743), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n760), .B(new_n761), .C1(new_n744), .C2(KEYINPUT93), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n724), .B1(new_n746), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n738), .A2(new_n743), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n725), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n761), .A2(new_n760), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT36), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(KEYINPUT94), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n766), .A2(new_n767), .A3(new_n769), .A4(new_n745), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n750), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n750), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(KEYINPUT29), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(KEYINPUT29), .ZN(new_n776));
  OAI21_X1  g351(.A(G2090), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n773), .A2(KEYINPUT29), .ZN(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n778), .A2(new_n779), .A3(new_n774), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n732), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n732), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT101), .B(G1966), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AND3_X1   g359(.A1(new_n777), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n750), .A2(G33), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n509), .A2(G139), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT25), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  INV_X1    g365(.A(G127), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n517), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n789), .B1(new_n463), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n786), .B1(new_n794), .B2(G29), .ZN(new_n795));
  INV_X1    g370(.A(G2072), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT97), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n750), .A2(G32), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT26), .Z(new_n801));
  INV_X1    g376(.A(G129), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n513), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n509), .B2(G141), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n653), .A2(G105), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT99), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n799), .B1(new_n808), .B2(new_n750), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT27), .B(G1996), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(G160), .A2(G29), .ZN(new_n813));
  INV_X1    g388(.A(G34), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(KEYINPUT24), .ZN(new_n815));
  AOI21_X1  g390(.A(G29), .B1(new_n814), .B2(KEYINPUT24), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(KEYINPUT98), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(KEYINPUT98), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G2084), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n795), .A2(new_n796), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n798), .A2(new_n812), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  INV_X1    g402(.A(G1961), .ZN(new_n828));
  NAND2_X1  g403(.A1(G301), .A2(G16), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n732), .A2(G5), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n650), .A2(new_n750), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT31), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(G11), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(G11), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT30), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(G28), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n750), .B1(new_n836), .B2(G28), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n834), .B(new_n835), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n831), .A2(new_n832), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G19), .ZN(new_n841));
  OR3_X1    g416(.A1(new_n841), .A2(KEYINPUT95), .A3(G16), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT95), .B1(new_n841), .B2(G16), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n842), .B(new_n843), .C1(new_n588), .C2(new_n732), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(G1341), .Z(new_n845));
  NAND3_X1  g420(.A1(new_n829), .A2(new_n828), .A3(new_n830), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n732), .A2(G4), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n638), .B2(new_n732), .ZN(new_n848));
  INV_X1    g423(.A(G1348), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n840), .A2(new_n845), .A3(new_n846), .A4(new_n850), .ZN(new_n851));
  OAI221_X1 g426(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n462), .C2(G116), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n504), .A2(G128), .A3(new_n463), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n509), .A2(KEYINPUT96), .A3(G140), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT96), .B1(new_n509), .B2(G140), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G29), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n750), .A2(G26), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT28), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G2067), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n809), .A2(new_n811), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n750), .A2(G27), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(G164), .B2(new_n750), .ZN(new_n864));
  INV_X1    g439(.A(G2078), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT102), .B(KEYINPUT23), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n732), .A2(G20), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G299), .B2(G16), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G1956), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n819), .A2(new_n820), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n862), .A2(new_n866), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n851), .A2(new_n861), .A3(new_n873), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n785), .A2(new_n826), .A3(new_n827), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n771), .A2(new_n875), .ZN(G311));
  OAI21_X1  g451(.A(KEYINPUT103), .B1(new_n771), .B2(new_n875), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n826), .A3(new_n827), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n777), .A2(new_n780), .A3(new_n784), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n770), .A4(new_n763), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n877), .A2(new_n882), .ZN(G150));
  NAND2_X1  g458(.A1(G80), .A2(G543), .ZN(new_n884));
  INV_X1    g459(.A(G67), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n581), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(G651), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n552), .A2(G55), .B1(G93), .B2(new_n559), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT104), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n588), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n587), .A2(new_n889), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n630), .A2(new_n639), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n895), .B(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT39), .ZN(new_n900));
  AOI21_X1  g475(.A(G860), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n900), .B2(new_n899), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT106), .Z(new_n903));
  NAND2_X1  g478(.A1(new_n891), .A2(new_n892), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G860), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(KEYINPUT37), .Z(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(G145));
  XNOR2_X1  g482(.A(new_n807), .B(new_n794), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n509), .A2(G142), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n504), .A2(G130), .A3(new_n463), .ZN(new_n910));
  OAI21_X1  g485(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT109), .Z(new_n912));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n462), .A2(G118), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n917), .A2(new_n655), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n655), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n908), .B(new_n920), .Z(new_n921));
  AND3_X1   g496(.A1(new_n530), .A2(KEYINPUT107), .A3(new_n535), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT107), .B1(new_n530), .B2(new_n535), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n856), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n755), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n856), .A2(new_n924), .ZN(new_n927));
  INV_X1    g502(.A(new_n755), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n856), .A2(new_n924), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n921), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n908), .B(new_n920), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n926), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n649), .B(G160), .Z(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(G162), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT110), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n932), .A2(new_n934), .A3(new_n940), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n935), .B2(new_n938), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n942), .A2(KEYINPUT40), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT40), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(G395));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n904), .B2(new_n631), .ZN(new_n948));
  OR3_X1    g523(.A1(new_n893), .A2(new_n642), .A3(new_n894), .ZN(new_n949));
  AND2_X1   g524(.A1(G299), .A2(new_n630), .ZN(new_n950));
  NOR2_X1   g525(.A1(G299), .A2(new_n630), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n642), .B1(new_n893), .B2(new_n894), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT111), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n949), .A2(new_n956), .A3(new_n952), .A4(new_n953), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n949), .A2(new_n953), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n638), .A2(new_n596), .A3(new_n600), .ZN(new_n960));
  NAND2_X1  g535(.A1(G299), .A2(new_n630), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n960), .A2(KEYINPUT41), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT41), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n959), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n959), .B2(new_n964), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n958), .B(KEYINPUT113), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(G290), .B(new_n615), .ZN(new_n970));
  XNOR2_X1  g545(.A(G288), .B(G303), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n971), .ZN(new_n973));
  INV_X1    g548(.A(G290), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(new_n615), .ZN(new_n975));
  NOR2_X1   g550(.A1(G290), .A2(G305), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT42), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n969), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n968), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n966), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT113), .B1(new_n982), .B2(new_n958), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n978), .B(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n967), .A2(new_n968), .ZN(new_n988));
  INV_X1    g563(.A(new_n958), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n986), .B(new_n987), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G868), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n948), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n969), .A3(new_n979), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n994), .A2(new_n947), .A3(G868), .A4(new_n990), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n992), .A2(new_n995), .ZN(G295));
  AND2_X1   g571(.A1(new_n992), .A2(new_n995), .ZN(G331));
  NAND3_X1  g572(.A1(new_n566), .A2(new_n570), .A3(G301), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(G301), .B1(new_n566), .B2(new_n570), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n999), .A2(new_n1000), .B1(new_n893), .B2(new_n894), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1000), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1002), .A2(new_n895), .A3(new_n998), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1001), .A2(new_n1003), .A3(new_n952), .ZN(new_n1004));
  INV_X1    g579(.A(new_n964), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n978), .ZN(new_n1008));
  AOI21_X1  g583(.A(G37), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n978), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1001), .A2(new_n1003), .A3(new_n952), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1008), .B(new_n1014), .C1(new_n1015), .C2(new_n1005), .ZN(new_n1016));
  INV_X1    g591(.A(G37), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1012), .A2(new_n1016), .A3(new_n1011), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT115), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1012), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1013), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(KEYINPUT44), .A3(new_n1018), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(G397));
  NAND2_X1  g601(.A1(new_n496), .A2(new_n502), .ZN(new_n1027));
  INV_X1    g602(.A(G125), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n476), .B2(new_n477), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n480), .B1(new_n1029), .B2(KEYINPUT70), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n470), .A2(new_n471), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n463), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1027), .A2(new_n1032), .A3(G40), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n530), .B2(new_n535), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n740), .A2(G1976), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(G8), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT52), .ZN(new_n1038));
  INV_X1    g613(.A(G1384), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n536), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1027), .A2(new_n1032), .A3(G40), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n614), .A2(G1981), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n611), .A2(new_n613), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1035), .A2(new_n1036), .A3(G8), .A4(new_n1056), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1038), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1041), .B1(new_n1060), .B2(new_n1040), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT107), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n536), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n530), .A2(KEYINPUT107), .A3(new_n535), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(KEYINPUT45), .A3(new_n1039), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n735), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1040), .A2(KEYINPUT50), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1034), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1068), .A2(new_n779), .A3(new_n1033), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1059), .B1(new_n1072), .B2(G8), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1971), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1034), .A2(new_n1069), .ZN(new_n1075));
  AOI211_X1 g650(.A(KEYINPUT50), .B(G1384), .C1(new_n530), .C2(new_n535), .ZN(new_n1076));
  NOR4_X1   g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n1041), .A4(G2090), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1059), .B(G8), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(G303), .A2(G8), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT55), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1058), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT120), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1084), .B(new_n1058), .C1(new_n1073), .C2(new_n1081), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1080), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1086), .B(G8), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(G160), .B(G40), .C1(new_n1034), .C2(KEYINPUT45), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1034), .A2(KEYINPUT45), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n783), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1068), .A2(new_n820), .A3(new_n1033), .A4(new_n1070), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1043), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G168), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT63), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1088), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1083), .A2(new_n1085), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(G8), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1080), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n1058), .A3(new_n1087), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1095), .B1(new_n1100), .B2(new_n1094), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1088), .A2(new_n1058), .ZN(new_n1103));
  AOI211_X1 g678(.A(G1976), .B(G288), .C1(new_n1044), .C2(new_n1053), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1049), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1044), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1091), .A2(G168), .A3(new_n1092), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1043), .B1(KEYINPUT122), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(KEYINPUT122), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1108), .B(new_n1110), .C1(KEYINPUT122), .C2(new_n1109), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1093), .A2(G286), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1111), .A2(new_n1112), .B1(G286), .B2(new_n1093), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(KEYINPUT62), .A3(new_n1114), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1061), .A2(new_n865), .A3(new_n1065), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(G160), .B(G40), .C1(new_n1034), .C2(new_n1069), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n828), .B1(new_n1125), .B2(new_n1076), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1123), .A2(G2078), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1061), .B(new_n1128), .C1(new_n1060), .C2(new_n1040), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(new_n1100), .A3(G301), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1107), .B1(new_n1121), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT57), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(KEYINPUT57), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(G299), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1136), .B1(G299), .B2(new_n1134), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1061), .A2(new_n1065), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1956), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1125), .B2(new_n1076), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n849), .B1(new_n1125), .B2(new_n1076), .ZN(new_n1145));
  INV_X1    g720(.A(G2067), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1042), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n630), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1141), .A2(new_n1143), .A3(new_n1139), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1144), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1139), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1153), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n1155));
  INV_X1    g730(.A(G1996), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1061), .A2(new_n1156), .A3(new_n1065), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT58), .B(G1341), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n1035), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1155), .B1(new_n1160), .B2(new_n588), .ZN(new_n1161));
  AOI211_X1 g736(.A(KEYINPUT59), .B(new_n587), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1154), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1141), .A2(new_n1143), .A3(new_n1139), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n1144), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1167), .A2(KEYINPUT60), .A3(new_n638), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n630), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n638), .A2(KEYINPUT60), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1145), .A2(new_n1147), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1166), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1150), .B1(new_n1163), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT45), .B1(new_n924), .B2(new_n1039), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1065), .A2(new_n1033), .A3(new_n1128), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1124), .B(new_n1126), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(G171), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT123), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1180), .A3(G171), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1127), .A2(G301), .A3(new_n1129), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1179), .A2(KEYINPUT54), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT54), .ZN(new_n1184));
  AOI21_X1  g759(.A(G301), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1177), .A2(G171), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1100), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1174), .A2(new_n1183), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1102), .A2(new_n1132), .A3(new_n1189), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1175), .A2(new_n1033), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1191), .A2(new_n693), .A3(new_n974), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1191), .A2(G1986), .A3(G290), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT116), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n856), .B(new_n1146), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT117), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n807), .B(new_n1156), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n755), .B(new_n757), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1195), .B1(new_n1191), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1190), .A2(new_n1202), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n1196), .A2(KEYINPUT117), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1196), .A2(KEYINPUT117), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1191), .B1(new_n1206), .B2(new_n807), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT47), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1191), .A2(new_n1156), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT46), .ZN(new_n1210));
  AND3_X1   g785(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1208), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1201), .A2(new_n1191), .ZN(new_n1213));
  XOR2_X1   g788(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1214));
  XOR2_X1   g789(.A(new_n1192), .B(new_n1214), .Z(new_n1215));
  OAI22_X1  g790(.A1(new_n1211), .A2(new_n1212), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1191), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n928), .A2(new_n757), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT124), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1204), .A2(new_n1219), .A3(new_n1205), .A4(new_n1199), .ZN(new_n1220));
  OR2_X1    g795(.A1(new_n856), .A2(G2067), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1217), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1216), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1203), .A2(new_n1225), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g801(.A(G319), .B1(new_n675), .B2(new_n676), .ZN(new_n1228));
  NOR2_X1   g802(.A1(G227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n719), .A2(new_n1229), .A3(new_n722), .ZN(new_n1230));
  OR2_X1    g804(.A1(new_n1230), .A2(KEYINPUT127), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n1230), .A2(KEYINPUT127), .ZN(new_n1232));
  AOI22_X1  g806(.A1(new_n942), .A2(new_n943), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1233), .A2(new_n1022), .ZN(G225));
  INV_X1    g808(.A(G225), .ZN(G308));
endmodule


