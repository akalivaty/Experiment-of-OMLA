//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1124,
    new_n1125, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(KEYINPUT3), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n468), .A2(G137), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n471), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n471), .B2(new_n478), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G125), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n477), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n476), .B1(G2105), .B2(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n468), .A2(new_n471), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT72), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n486), .A2(new_n469), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT73), .B1(G100), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NOR3_X1   g068(.A1(KEYINPUT73), .A2(G100), .A3(G2105), .ZN(new_n494));
  OAI221_X1 g069(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n489), .A2(new_n496), .ZN(G162));
  OAI211_X1 g072(.A(G138), .B(new_n469), .C1(new_n480), .C2(new_n481), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n468), .A2(new_n471), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT74), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n468), .A2(new_n504), .A3(new_n471), .A4(new_n501), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT4), .A2(G138), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n468), .A2(new_n469), .A3(new_n471), .A4(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(G102), .A2(G2105), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n509), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n500), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n514), .A2(new_n515), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT5), .B(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n519), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n523), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT75), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n518), .A2(G51), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n533), .A2(new_n534), .A3(new_n536), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(new_n518), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n523), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT77), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(KEYINPUT77), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT5), .B(G543), .Z(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n543), .A2(new_n544), .B1(G651), .B2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n526), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n546), .A2(new_n516), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G81), .B1(new_n518), .B2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT78), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n518), .A2(G53), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n546), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n552), .B2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n552), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n518), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n552), .A2(G86), .B1(new_n518), .B2(G48), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n546), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n578), .A2(KEYINPUT79), .A3(G651), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n522), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n526), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n575), .A2(new_n579), .A3(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n518), .A2(G47), .ZN(new_n584));
  XOR2_X1   g159(.A(KEYINPUT80), .B(G85), .Z(new_n585));
  AOI22_X1  g160(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n523), .B2(new_n585), .C1(new_n526), .C2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n522), .A2(G66), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT82), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n526), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(G54), .B2(new_n518), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n552), .A2(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G299), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G168), .B2(new_n603), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(G168), .B2(new_n603), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n554), .A2(new_n603), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n599), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g187(.A1(new_n480), .A2(new_n481), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n466), .A2(new_n467), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n613), .A2(new_n469), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT84), .B(G2100), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n487), .A2(G135), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n490), .A2(G123), .ZN(new_n622));
  NOR3_X1   g197(.A1(new_n469), .A2(KEYINPUT85), .A3(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT85), .B1(new_n469), .B2(G111), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(G2104), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n619), .A2(new_n620), .A3(new_n628), .ZN(G156));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n633), .B(new_n639), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(G14), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n641), .ZN(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n646), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n647), .B2(new_n648), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT87), .Z(new_n654));
  XOR2_X1   g229(.A(new_n648), .B(KEYINPUT17), .Z(new_n655));
  AOI21_X1  g230(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n654), .B1(new_n646), .B2(new_n655), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n656), .B1(new_n657), .B2(new_n647), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n662), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G22), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G166), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1971), .ZN(new_n682));
  OR2_X1    g257(.A1(G6), .A2(G16), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G305), .B2(new_n679), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  AOI21_X1  g260(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(G16), .A2(G23), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT92), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G288), .B2(new_n679), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT33), .ZN(new_n690));
  INV_X1    g265(.A(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n686), .B(new_n692), .C1(new_n684), .C2(new_n685), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT34), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G25), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n490), .A2(G119), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(G95), .A2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n700), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n487), .A2(G131), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n696), .B1(new_n705), .B2(new_n695), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT91), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n708), .ZN(new_n710));
  MUX2_X1   g285(.A(G24), .B(G290), .S(G16), .Z(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(G1986), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n694), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT36), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n695), .A2(G35), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G162), .B2(new_n695), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G2090), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n627), .A2(new_n695), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT97), .Z(new_n722));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n723), .A2(G28), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n695), .B1(new_n723), .B2(G28), .ZN(new_n725));
  AND2_X1   g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  NOR2_X1   g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n555), .A2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G16), .B2(G19), .ZN(new_n730));
  INV_X1    g305(.A(G1341), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n722), .B(new_n732), .C1(new_n731), .C2(new_n730), .ZN(new_n733));
  NOR2_X1   g308(.A1(G5), .A2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT98), .Z(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G171), .B2(G16), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT95), .B(G2067), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n695), .A2(G26), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT28), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n487), .A2(G140), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n490), .A2(G128), .ZN(new_n742));
  OAI21_X1  g317(.A(KEYINPUT94), .B1(G104), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(KEYINPUT94), .A2(G104), .A3(G2105), .ZN(new_n745));
  OAI221_X1 g320(.A(G2104), .B1(G116), .B2(new_n469), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n741), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n740), .B1(new_n748), .B2(new_n695), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n737), .A2(G1961), .B1(new_n738), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n733), .A2(new_n750), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n737), .A2(G1961), .B1(new_n738), .B2(new_n749), .ZN(new_n752));
  NOR2_X1   g327(.A1(G160), .A2(new_n695), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n695), .B1(KEYINPUT24), .B2(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(KEYINPUT24), .B2(G34), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2084), .ZN(new_n757));
  AND3_X1   g332(.A1(new_n751), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n679), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n679), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1966), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n512), .A2(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n695), .A2(G27), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n761), .B1(G2078), .B2(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n758), .B(new_n766), .C1(G2078), .C2(new_n765), .ZN(new_n767));
  NOR2_X1   g342(.A1(G4), .A2(G16), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n600), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT93), .B(G1348), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n695), .A2(G32), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n487), .A2(G141), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n490), .A2(G129), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT26), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  AOI22_X1  g353(.A1(G105), .A2(new_n473), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n773), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n772), .B1(new_n781), .B2(new_n695), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT27), .B(G1996), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n679), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT23), .ZN(new_n786));
  INV_X1    g361(.A(G299), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n679), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1956), .Z(new_n789));
  OR2_X1    g364(.A1(new_n782), .A2(new_n783), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n771), .A2(new_n784), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n695), .A2(G33), .ZN(new_n792));
  NAND2_X1  g367(.A1(G115), .A2(G2104), .ZN(new_n793));
  INV_X1    g368(.A(G127), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n482), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n469), .B1(new_n795), .B2(KEYINPUT96), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(KEYINPUT96), .B2(new_n795), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT25), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n487), .B2(G139), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n792), .B1(new_n802), .B2(new_n695), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2072), .ZN(new_n804));
  OR4_X1    g379(.A1(new_n720), .A2(new_n767), .A3(new_n791), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n715), .A2(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  AOI22_X1  g382(.A1(new_n552), .A2(G93), .B1(new_n518), .B2(G55), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT100), .Z(new_n809));
  AOI22_X1  g384(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(new_n526), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT101), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT101), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n809), .A2(new_n814), .A3(new_n811), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n813), .A2(new_n554), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n812), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n817), .A2(new_n814), .A3(new_n555), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n600), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n823));
  AOI21_X1  g398(.A(G860), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n812), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G145));
  XNOR2_X1  g403(.A(KEYINPUT104), .B(G37), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n512), .B(new_n747), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n703), .B(KEYINPUT90), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n801), .A2(new_n780), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n802), .A2(new_n781), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n833), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(new_n705), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n831), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n487), .A2(G142), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n490), .A2(G130), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n469), .A2(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n616), .B(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n835), .A2(new_n837), .A3(new_n831), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n839), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  INV_X1    g423(.A(new_n846), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(new_n838), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(G162), .B(new_n627), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G160), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n856), .A2(new_n847), .A3(new_n850), .A4(new_n851), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n830), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n860), .B(new_n862), .ZN(G395));
  AOI21_X1  g438(.A(new_n787), .B1(new_n595), .B2(new_n598), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n595), .A2(new_n787), .A3(new_n598), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT41), .B1(new_n868), .B2(new_n864), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(new_n870), .A3(new_n866), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT107), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n867), .B2(KEYINPUT41), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n819), .B(new_n610), .ZN(new_n876));
  MUX2_X1   g451(.A(new_n867), .B(new_n875), .S(new_n876), .Z(new_n877));
  XOR2_X1   g452(.A(G305), .B(G290), .Z(new_n878));
  XNOR2_X1  g453(.A(G166), .B(G288), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT42), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n877), .A2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(G868), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(G868), .B2(new_n817), .ZN(G295));
  OAI21_X1  g462(.A(new_n886), .B1(G868), .B2(new_n817), .ZN(G331));
  XNOR2_X1  g463(.A(G171), .B(G286), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n816), .A2(new_n889), .A3(new_n818), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n816), .B2(new_n818), .ZN(new_n892));
  OAI22_X1  g467(.A1(new_n872), .A2(new_n874), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n894), .A2(new_n865), .A3(new_n866), .A4(new_n890), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n895), .A3(new_n882), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n880), .A2(KEYINPUT108), .A3(new_n881), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT108), .B1(new_n880), .B2(new_n881), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n893), .B2(new_n895), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n894), .A2(new_n890), .B1(new_n869), .B2(new_n871), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n891), .A2(new_n892), .A3(new_n867), .ZN(new_n906));
  OAI22_X1  g481(.A1(new_n905), .A2(new_n906), .B1(new_n899), .B2(new_n900), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n907), .A2(new_n896), .A3(new_n908), .A4(new_n829), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n896), .A3(new_n829), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n898), .A2(KEYINPUT43), .A3(new_n902), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n910), .B1(new_n917), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g493(.A(G1384), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n512), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n472), .A2(G40), .A3(new_n474), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n484), .B2(G2105), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n925));
  XNOR2_X1  g500(.A(KEYINPUT56), .B(G2072), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n922), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT118), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT45), .B1(new_n512), .B2(new_n919), .ZN(new_n929));
  INV_X1    g504(.A(new_n924), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT118), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n925), .A4(new_n926), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n563), .A2(new_n567), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n563), .B2(new_n567), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n512), .A2(new_n939), .A3(new_n919), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT115), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n920), .A2(KEYINPUT50), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT115), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n512), .A2(new_n943), .A3(new_n939), .A4(new_n919), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n941), .A2(new_n942), .A3(new_n924), .A4(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(KEYINPUT116), .B(G1956), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n938), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n934), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n938), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n934), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT119), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n508), .A2(new_n510), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n499), .B2(new_n498), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n954), .B2(new_n506), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n924), .B1(new_n955), .B2(new_n939), .ZN(new_n956));
  INV_X1    g531(.A(new_n940), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n930), .B1(new_n920), .B2(KEYINPUT50), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(KEYINPUT119), .A3(new_n940), .ZN(new_n960));
  INV_X1    g535(.A(G1348), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G2067), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n955), .A2(new_n963), .A3(new_n924), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n599), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n948), .B1(new_n951), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT121), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n934), .A2(new_n950), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n968), .A2(new_n938), .B1(new_n934), .B2(new_n947), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n969), .B2(KEYINPUT61), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT61), .ZN(new_n971));
  INV_X1    g546(.A(new_n948), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT121), .B(new_n971), .C1(new_n972), .C2(new_n951), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n938), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT122), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n948), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n934), .A2(KEYINPUT122), .A3(new_n947), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n975), .A2(new_n977), .A3(KEYINPUT61), .A4(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n962), .A2(KEYINPUT60), .A3(new_n964), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n599), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n962), .A2(new_n964), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT60), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n962), .A2(KEYINPUT60), .A3(new_n600), .A4(new_n964), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n955), .A2(new_n924), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT58), .B(G1341), .Z(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT120), .B(G1996), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n555), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT59), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n979), .A2(new_n986), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n966), .B1(new_n974), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1961), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n958), .A2(new_n960), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G2078), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n931), .A2(new_n999), .A3(new_n925), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(G171), .B(KEYINPUT54), .Z(new_n1006));
  NAND2_X1  g581(.A1(new_n484), .A2(KEYINPUT123), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n484), .A2(KEYINPUT123), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(new_n469), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n923), .B(new_n929), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(KEYINPUT124), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n925), .A2(KEYINPUT53), .A3(new_n999), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n1010), .B2(KEYINPUT124), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1006), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1005), .A2(new_n1006), .B1(new_n1014), .B2(new_n1003), .ZN(new_n1015));
  INV_X1    g590(.A(G1966), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n990), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2084), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n959), .A2(new_n1018), .A3(new_n940), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(G168), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G8), .ZN(new_n1021));
  AOI21_X1  g596(.A(G168), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT51), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1024), .A3(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n571), .A2(new_n573), .A3(G1976), .A4(new_n572), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n987), .A2(G8), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT52), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n691), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n987), .A2(new_n1029), .A3(G8), .A4(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n987), .A2(G8), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n579), .A2(new_n582), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G1981), .ZN(new_n1038));
  INV_X1    g613(.A(G305), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(G305), .A2(new_n1037), .A3(G1981), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT49), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1035), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(KEYINPUT114), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(KEYINPUT114), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  INV_X1    g623(.A(G1971), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n990), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G2090), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n959), .A2(new_n1051), .A3(new_n941), .A4(new_n944), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1048), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G166), .A2(new_n1048), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT55), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1034), .B(new_n1047), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n959), .A2(KEYINPUT110), .A3(new_n1051), .A4(new_n940), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n940), .A2(new_n1051), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n956), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1050), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(G8), .A3(new_n1055), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT111), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1061), .A2(new_n1064), .A3(G8), .A4(new_n1055), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1056), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1015), .A2(new_n1026), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n996), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1023), .A2(new_n1069), .A3(new_n1025), .ZN(new_n1070));
  AOI21_X1  g645(.A(G301), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1066), .A2(new_n1070), .A3(KEYINPUT125), .A4(new_n1071), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1034), .A2(new_n1047), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1079));
  NOR2_X1   g654(.A1(G286), .A2(new_n1048), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT63), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1055), .B2(new_n1053), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1078), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1034), .A2(new_n1047), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1055), .B1(new_n1061), .B2(G8), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT63), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(G305), .A2(G1981), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G288), .A2(G1976), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1047), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1091), .B2(new_n1035), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1085), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1068), .A2(new_n1077), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n922), .A2(new_n930), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n832), .A2(new_n708), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n832), .A2(new_n708), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n747), .B(new_n963), .ZN(new_n1098));
  INV_X1    g673(.A(G1996), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n780), .B(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(G290), .B(G1986), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1095), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1094), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n1096), .A2(new_n1105), .B1(G2067), .B2(new_n747), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1095), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1107), .B(KEYINPUT126), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1101), .A2(new_n1095), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G290), .A2(G1986), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1095), .A2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1111), .B(KEYINPUT127), .Z(new_n1112));
  OAI21_X1  g687(.A(new_n1109), .B1(KEYINPUT48), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(KEYINPUT48), .B2(new_n1112), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1115), .A2(KEYINPUT46), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(KEYINPUT46), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1098), .A2(new_n781), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1116), .A2(new_n1117), .B1(new_n1095), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT47), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1108), .A2(new_n1114), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1104), .A2(new_n1121), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g697(.A(new_n860), .ZN(new_n1124));
  NAND2_X1  g698(.A1(new_n903), .A2(new_n909), .ZN(new_n1125));
  INV_X1    g699(.A(G319), .ZN(new_n1126));
  NOR4_X1   g700(.A1(G229), .A2(new_n1126), .A3(G401), .A4(G227), .ZN(new_n1127));
  AND3_X1   g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(G308));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(G225));
endmodule


