

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769;

  XNOR2_X1 U375 ( .A(n576), .B(KEYINPUT38), .ZN(n685) );
  NOR2_X2 U376 ( .A1(n640), .A2(n742), .ZN(n641) );
  NOR2_X2 U377 ( .A1(n646), .A2(n742), .ZN(n648) );
  NOR2_X2 U378 ( .A1(n655), .A2(n742), .ZN(n657) );
  XNOR2_X2 U379 ( .A(n414), .B(KEYINPUT41), .ZN(n726) );
  XNOR2_X1 U380 ( .A(G122), .B(G113), .ZN(n426) );
  XNOR2_X1 U381 ( .A(n532), .B(n531), .ZN(n591) );
  XNOR2_X1 U382 ( .A(n413), .B(n540), .ZN(n570) );
  XNOR2_X1 U383 ( .A(n416), .B(n550), .ZN(n568) );
  XNOR2_X1 U384 ( .A(n373), .B(KEYINPUT33), .ZN(n727) );
  NAND2_X1 U385 ( .A1(n415), .A2(n537), .ZN(n414) );
  NOR2_X1 U386 ( .A1(n739), .A2(G902), .ZN(n516) );
  XNOR2_X1 U387 ( .A(n419), .B(n418), .ZN(n739) );
  XNOR2_X1 U388 ( .A(n420), .B(n510), .ZN(n419) );
  XNOR2_X1 U389 ( .A(n363), .B(G119), .ZN(n498) );
  XNOR2_X1 U390 ( .A(n424), .B(G110), .ZN(n490) );
  XNOR2_X1 U391 ( .A(n426), .B(G104), .ZN(n467) );
  INV_X2 U392 ( .A(G953), .ZN(n760) );
  XNOR2_X1 U393 ( .A(G101), .B(KEYINPUT3), .ZN(n363) );
  XNOR2_X1 U394 ( .A(KEYINPUT69), .B(KEYINPUT88), .ZN(n424) );
  XNOR2_X2 U395 ( .A(n389), .B(KEYINPUT32), .ZN(n610) );
  XNOR2_X1 U396 ( .A(n390), .B(G143), .ZN(n448) );
  INV_X1 U397 ( .A(G128), .ZN(n390) );
  NAND2_X1 U398 ( .A1(n410), .A2(n501), .ZN(n409) );
  INV_X1 U399 ( .A(G469), .ZN(n410) );
  XNOR2_X1 U400 ( .A(n485), .B(n484), .ZN(n499) );
  XNOR2_X1 U401 ( .A(n541), .B(KEYINPUT64), .ZN(n555) );
  XNOR2_X1 U402 ( .A(n616), .B(n544), .ZN(n417) );
  XNOR2_X1 U403 ( .A(n477), .B(n476), .ZN(n557) );
  XNOR2_X1 U404 ( .A(n461), .B(n460), .ZN(n558) );
  NOR2_X1 U405 ( .A1(n394), .A2(KEYINPUT44), .ZN(n393) );
  XNOR2_X1 U406 ( .A(G137), .B(G113), .ZN(n496) );
  NAND2_X1 U407 ( .A1(n494), .A2(G210), .ZN(n380) );
  XNOR2_X1 U408 ( .A(n379), .B(G146), .ZN(n378) );
  INV_X1 U409 ( .A(G116), .ZN(n379) );
  NOR2_X1 U410 ( .A1(G953), .A2(G237), .ZN(n494) );
  XNOR2_X1 U411 ( .A(n716), .B(KEYINPUT70), .ZN(n371) );
  XNOR2_X1 U412 ( .A(G146), .B(G125), .ZN(n470) );
  XNOR2_X1 U413 ( .A(n448), .B(KEYINPUT4), .ZN(n485) );
  NAND2_X1 U414 ( .A1(G234), .A2(G237), .ZN(n441) );
  XNOR2_X1 U415 ( .A(n365), .B(n364), .ZN(n415) );
  INV_X1 U416 ( .A(KEYINPUT106), .ZN(n364) );
  NAND2_X1 U417 ( .A1(n685), .A2(n684), .ZN(n365) );
  BUF_X1 U418 ( .A(n555), .Z(n698) );
  XNOR2_X1 U419 ( .A(n382), .B(G472), .ZN(n556) );
  XNOR2_X1 U420 ( .A(n507), .B(n421), .ZN(n420) );
  XNOR2_X1 U421 ( .A(n509), .B(n506), .ZN(n421) );
  XNOR2_X1 U422 ( .A(G119), .B(G128), .ZN(n502) );
  XOR2_X1 U423 ( .A(KEYINPUT24), .B(G110), .Z(n503) );
  XNOR2_X1 U424 ( .A(G116), .B(G107), .ZN(n455) );
  XNOR2_X1 U425 ( .A(G122), .B(KEYINPUT98), .ZN(n447) );
  XNOR2_X1 U426 ( .A(n392), .B(n391), .ZN(n559) );
  INV_X1 U427 ( .A(KEYINPUT34), .ZN(n391) );
  OR2_X1 U428 ( .A1(n652), .A2(n630), .ZN(n439) );
  NAND2_X1 U429 ( .A1(n543), .A2(n542), .ZN(n616) );
  XNOR2_X1 U430 ( .A(n483), .B(n482), .ZN(n625) );
  OR2_X1 U431 ( .A1(n613), .A2(n481), .ZN(n483) );
  XNOR2_X1 U432 ( .A(n556), .B(KEYINPUT6), .ZN(n622) );
  NAND2_X1 U433 ( .A1(n406), .A2(n411), .ZN(n399) );
  AND2_X1 U434 ( .A1(n404), .A2(n401), .ZN(n400) );
  NAND2_X1 U435 ( .A1(G902), .A2(G469), .ZN(n412) );
  XNOR2_X1 U436 ( .A(n376), .B(KEYINPUT45), .ZN(n632) );
  NAND2_X1 U437 ( .A1(n375), .A2(n374), .ZN(n376) );
  NAND2_X1 U438 ( .A1(n356), .A2(n395), .ZN(n374) );
  XNOR2_X1 U439 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n430) );
  NAND2_X1 U440 ( .A1(n608), .A2(n423), .ZN(n633) );
  INV_X1 U441 ( .A(G237), .ZN(n436) );
  NAND2_X1 U442 ( .A1(KEYINPUT1), .A2(n403), .ZN(n402) );
  INV_X1 U443 ( .A(n409), .ZN(n403) );
  XNOR2_X1 U444 ( .A(n381), .B(n377), .ZN(n500) );
  XNOR2_X1 U445 ( .A(n380), .B(n378), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n498), .B(n497), .ZN(n381) );
  XNOR2_X1 U447 ( .A(KEYINPUT67), .B(KEYINPUT16), .ZN(n425) );
  BUF_X1 U448 ( .A(n632), .Z(n750) );
  XNOR2_X1 U449 ( .A(G131), .B(KEYINPUT12), .ZN(n462) );
  XOR2_X1 U450 ( .A(KEYINPUT11), .B(KEYINPUT93), .Z(n463) );
  XNOR2_X1 U451 ( .A(n499), .B(n486), .ZN(n756) );
  XOR2_X1 U452 ( .A(G101), .B(G104), .Z(n488) );
  NAND2_X2 U453 ( .A1(n366), .A2(n631), .ZN(n635) );
  XNOR2_X1 U454 ( .A(n368), .B(n367), .ZN(n366) );
  INV_X1 U455 ( .A(KEYINPUT81), .ZN(n367) );
  BUF_X1 U456 ( .A(n716), .Z(n759) );
  NAND2_X1 U457 ( .A1(n372), .A2(n563), .ZN(n373) );
  NOR2_X1 U458 ( .A1(n698), .A2(n622), .ZN(n372) );
  XNOR2_X1 U459 ( .A(n386), .B(KEYINPUT0), .ZN(n613) );
  XNOR2_X1 U460 ( .A(n388), .B(n387), .ZN(n530) );
  INV_X1 U461 ( .A(KEYINPUT19), .ZN(n387) );
  NOR2_X1 U462 ( .A1(n576), .A2(n536), .ZN(n388) );
  XNOR2_X1 U463 ( .A(n508), .B(n758), .ZN(n418) );
  XNOR2_X1 U464 ( .A(n459), .B(n458), .ZN(n735) );
  AND2_X1 U465 ( .A1(n639), .A2(G953), .ZN(n742) );
  XNOR2_X1 U466 ( .A(n562), .B(n561), .ZN(n611) );
  AND2_X1 U467 ( .A1(n417), .A2(n549), .ZN(n594) );
  AND2_X1 U468 ( .A1(n575), .A2(n383), .ZN(n354) );
  AND2_X1 U469 ( .A1(n635), .A2(n724), .ZN(n355) );
  XNOR2_X1 U470 ( .A(G137), .B(G140), .ZN(n505) );
  XNOR2_X1 U471 ( .A(n633), .B(KEYINPUT83), .ZN(n716) );
  AND2_X1 U472 ( .A1(n610), .A2(n393), .ZN(n356) );
  INV_X1 U473 ( .A(KEYINPUT1), .ZN(n407) );
  AND2_X1 U474 ( .A1(n397), .A2(KEYINPUT44), .ZN(n357) );
  INV_X1 U475 ( .A(n563), .ZN(n697) );
  NAND2_X1 U476 ( .A1(n400), .A2(n399), .ZN(n563) );
  AND2_X1 U477 ( .A1(n724), .A2(G475), .ZN(n358) );
  AND2_X1 U478 ( .A1(n724), .A2(G472), .ZN(n359) );
  AND2_X1 U479 ( .A1(n724), .A2(G210), .ZN(n360) );
  INV_X1 U480 ( .A(n576), .ZN(n383) );
  NOR2_X1 U481 ( .A1(n566), .A2(n565), .ZN(n361) );
  AND2_X1 U482 ( .A1(n549), .A2(n685), .ZN(n362) );
  INV_X1 U483 ( .A(n415), .ZN(n682) );
  NAND2_X1 U484 ( .A1(n371), .A2(n369), .ZN(n368) );
  XNOR2_X1 U485 ( .A(n629), .B(n370), .ZN(n369) );
  INV_X1 U486 ( .A(KEYINPUT82), .ZN(n370) );
  NOR2_X1 U487 ( .A1(n698), .A2(n697), .ZN(n612) );
  NAND2_X1 U488 ( .A1(n727), .A2(n617), .ZN(n392) );
  NOR2_X1 U489 ( .A1(n385), .A2(n357), .ZN(n375) );
  NOR2_X1 U490 ( .A1(n573), .A2(n622), .ZN(n574) );
  NAND2_X1 U491 ( .A1(n643), .A2(n501), .ZN(n382) );
  NAND2_X1 U492 ( .A1(n384), .A2(n575), .ZN(n603) );
  NAND2_X1 U493 ( .A1(n384), .A2(n354), .ZN(n578) );
  NOR2_X1 U494 ( .A1(n676), .A2(n536), .ZN(n384) );
  NAND2_X1 U495 ( .A1(n396), .A2(n628), .ZN(n385) );
  NAND2_X1 U496 ( .A1(n530), .A2(n446), .ZN(n386) );
  INV_X1 U497 ( .A(n625), .ZN(n567) );
  NAND2_X1 U498 ( .A1(n625), .A2(n361), .ZN(n389) );
  NAND2_X1 U499 ( .A1(n610), .A2(n609), .ZN(n397) );
  INV_X1 U500 ( .A(n609), .ZN(n394) );
  INV_X1 U501 ( .A(n611), .ZN(n395) );
  NAND2_X1 U502 ( .A1(n611), .A2(KEYINPUT44), .ZN(n396) );
  NAND2_X1 U503 ( .A1(n398), .A2(n412), .ZN(n405) );
  NAND2_X1 U504 ( .A1(n663), .A2(G469), .ZN(n398) );
  AND2_X1 U505 ( .A1(n408), .A2(n407), .ZN(n406) );
  OR2_X1 U506 ( .A1(n663), .A2(n409), .ZN(n408) );
  INV_X1 U507 ( .A(n405), .ZN(n411) );
  OR2_X1 U508 ( .A1(n663), .A2(n402), .ZN(n401) );
  NAND2_X1 U509 ( .A1(n405), .A2(KEYINPUT1), .ZN(n404) );
  NAND2_X1 U510 ( .A1(n411), .A2(n408), .ZN(n542) );
  NAND2_X1 U511 ( .A1(n726), .A2(n538), .ZN(n413) );
  XNOR2_X2 U512 ( .A(n439), .B(n438), .ZN(n576) );
  NAND2_X1 U513 ( .A1(n635), .A2(n358), .ZN(n638) );
  NAND2_X1 U514 ( .A1(n635), .A2(n359), .ZN(n645) );
  NAND2_X1 U515 ( .A1(n635), .A2(n360), .ZN(n654) );
  NAND2_X1 U516 ( .A1(n417), .A2(n362), .ZN(n416) );
  XNOR2_X1 U517 ( .A(n602), .B(n601), .ZN(n608) );
  XNOR2_X2 U518 ( .A(n516), .B(n515), .ZN(n694) );
  XOR2_X1 U519 ( .A(n592), .B(KEYINPUT74), .Z(n422) );
  AND2_X1 U520 ( .A1(n767), .A2(n607), .ZN(n423) );
  INV_X1 U521 ( .A(KEYINPUT5), .ZN(n495) );
  INV_X1 U522 ( .A(KEYINPUT48), .ZN(n601) );
  XNOR2_X1 U523 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U524 ( .A(KEYINPUT79), .ZN(n506) );
  INV_X1 U525 ( .A(KEYINPUT23), .ZN(n509) );
  NOR2_X1 U526 ( .A1(n573), .A2(n525), .ZN(n526) );
  XNOR2_X1 U527 ( .A(n457), .B(n456), .ZN(n458) );
  INV_X1 U528 ( .A(KEYINPUT104), .ZN(n544) );
  XNOR2_X1 U529 ( .A(n490), .B(n498), .ZN(n429) );
  XNOR2_X1 U530 ( .A(n455), .B(n425), .ZN(n427) );
  XNOR2_X1 U531 ( .A(n427), .B(n467), .ZN(n428) );
  XNOR2_X1 U532 ( .A(n429), .B(n428), .ZN(n743) );
  XNOR2_X1 U533 ( .A(n470), .B(n430), .ZN(n433) );
  NAND2_X1 U534 ( .A1(n760), .A2(G224), .ZN(n431) );
  XNOR2_X1 U535 ( .A(n431), .B(KEYINPUT89), .ZN(n432) );
  XNOR2_X1 U536 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U537 ( .A(n485), .B(n434), .ZN(n435) );
  XNOR2_X1 U538 ( .A(n743), .B(n435), .ZN(n652) );
  XNOR2_X1 U539 ( .A(G902), .B(KEYINPUT15), .ZN(n478) );
  INV_X1 U540 ( .A(n478), .ZN(n630) );
  INV_X1 U541 ( .A(G902), .ZN(n501) );
  NAND2_X1 U542 ( .A1(n501), .A2(n436), .ZN(n440) );
  NAND2_X1 U543 ( .A1(n440), .A2(G210), .ZN(n437) );
  XNOR2_X1 U544 ( .A(n437), .B(KEYINPUT90), .ZN(n438) );
  NAND2_X1 U545 ( .A1(n440), .A2(G214), .ZN(n684) );
  INV_X1 U546 ( .A(n684), .ZN(n536) );
  XNOR2_X1 U547 ( .A(n441), .B(KEYINPUT14), .ZN(n442) );
  XNOR2_X1 U548 ( .A(KEYINPUT68), .B(n442), .ZN(n443) );
  NAND2_X1 U549 ( .A1(G952), .A2(n443), .ZN(n714) );
  OR2_X1 U550 ( .A1(n714), .A2(G953), .ZN(n521) );
  NAND2_X1 U551 ( .A1(n443), .A2(G902), .ZN(n519) );
  NOR2_X1 U552 ( .A1(G898), .A2(n760), .ZN(n444) );
  XNOR2_X1 U553 ( .A(KEYINPUT91), .B(n444), .ZN(n744) );
  OR2_X1 U554 ( .A1(n519), .A2(n744), .ZN(n445) );
  NAND2_X1 U555 ( .A1(n521), .A2(n445), .ZN(n446) );
  XNOR2_X1 U556 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U557 ( .A(KEYINPUT97), .B(KEYINPUT9), .Z(n450) );
  XNOR2_X1 U558 ( .A(KEYINPUT99), .B(KEYINPUT7), .ZN(n449) );
  XNOR2_X1 U559 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U560 ( .A(n452), .B(n451), .Z(n459) );
  NAND2_X1 U561 ( .A1(n760), .A2(G234), .ZN(n454) );
  XNOR2_X1 U562 ( .A(KEYINPUT8), .B(KEYINPUT65), .ZN(n453) );
  XNOR2_X1 U563 ( .A(n454), .B(n453), .ZN(n504) );
  NAND2_X1 U564 ( .A1(G217), .A2(n504), .ZN(n457) );
  XNOR2_X1 U565 ( .A(n455), .B(G134), .ZN(n456) );
  NAND2_X1 U566 ( .A1(n735), .A2(n501), .ZN(n461) );
  INV_X1 U567 ( .A(G478), .ZN(n460) );
  XNOR2_X1 U568 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U569 ( .A(n464), .B(KEYINPUT94), .Z(n466) );
  XNOR2_X1 U570 ( .A(G143), .B(G140), .ZN(n465) );
  XNOR2_X1 U571 ( .A(n466), .B(n465), .ZN(n473) );
  INV_X1 U572 ( .A(n467), .ZN(n469) );
  NAND2_X1 U573 ( .A1(G214), .A2(n494), .ZN(n468) );
  XNOR2_X1 U574 ( .A(n469), .B(n468), .ZN(n471) );
  XNOR2_X1 U575 ( .A(n470), .B(KEYINPUT10), .ZN(n758) );
  XNOR2_X1 U576 ( .A(n471), .B(n758), .ZN(n472) );
  XNOR2_X1 U577 ( .A(n473), .B(n472), .ZN(n636) );
  NAND2_X1 U578 ( .A1(n636), .A2(n501), .ZN(n477) );
  XOR2_X1 U579 ( .A(KEYINPUT13), .B(KEYINPUT95), .Z(n475) );
  XNOR2_X1 U580 ( .A(KEYINPUT96), .B(G475), .ZN(n474) );
  XNOR2_X1 U581 ( .A(n475), .B(n474), .ZN(n476) );
  AND2_X1 U582 ( .A1(n558), .A2(n557), .ZN(n537) );
  NAND2_X1 U583 ( .A1(n478), .A2(G234), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n479), .B(KEYINPUT20), .ZN(n511) );
  AND2_X1 U585 ( .A1(n511), .A2(G221), .ZN(n480) );
  XNOR2_X1 U586 ( .A(n480), .B(KEYINPUT21), .ZN(n693) );
  NAND2_X1 U587 ( .A1(n537), .A2(n693), .ZN(n481) );
  INV_X1 U588 ( .A(KEYINPUT22), .ZN(n482) );
  XNOR2_X1 U589 ( .A(G134), .B(G131), .ZN(n484) );
  INV_X1 U590 ( .A(n505), .ZN(n486) );
  NAND2_X1 U591 ( .A1(G227), .A2(n760), .ZN(n487) );
  XNOR2_X1 U592 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U593 ( .A(n489), .B(G107), .Z(n492) );
  XNOR2_X1 U594 ( .A(n490), .B(G146), .ZN(n491) );
  XNOR2_X1 U595 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U596 ( .A(n756), .B(n493), .ZN(n663) );
  XNOR2_X1 U597 ( .A(n500), .B(n499), .ZN(n643) );
  INV_X1 U598 ( .A(n556), .ZN(n525) );
  INV_X1 U599 ( .A(n525), .ZN(n701) );
  XNOR2_X1 U600 ( .A(n503), .B(n502), .ZN(n510) );
  NAND2_X1 U601 ( .A1(G221), .A2(n504), .ZN(n508) );
  XNOR2_X1 U602 ( .A(n505), .B(KEYINPUT72), .ZN(n507) );
  XOR2_X1 U603 ( .A(KEYINPUT25), .B(KEYINPUT92), .Z(n513) );
  NAND2_X1 U604 ( .A1(n511), .A2(G217), .ZN(n512) );
  XNOR2_X1 U605 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U606 ( .A(n514), .B(KEYINPUT71), .ZN(n515) );
  NOR2_X1 U607 ( .A1(n701), .A2(n694), .ZN(n517) );
  NAND2_X1 U608 ( .A1(n697), .A2(n517), .ZN(n518) );
  OR2_X1 U609 ( .A1(n567), .A2(n518), .ZN(n609) );
  XNOR2_X1 U610 ( .A(n609), .B(G110), .ZN(G12) );
  XNOR2_X1 U611 ( .A(G128), .B(KEYINPUT29), .ZN(n535) );
  OR2_X1 U612 ( .A1(n760), .A2(n519), .ZN(n520) );
  NOR2_X1 U613 ( .A1(G900), .A2(n520), .ZN(n523) );
  INV_X1 U614 ( .A(n521), .ZN(n522) );
  NOR2_X1 U615 ( .A1(n523), .A2(n522), .ZN(n546) );
  NOR2_X1 U616 ( .A1(n694), .A2(n546), .ZN(n524) );
  NAND2_X1 U617 ( .A1(n524), .A2(n693), .ZN(n573) );
  XNOR2_X1 U618 ( .A(n526), .B(KEYINPUT28), .ZN(n529) );
  INV_X1 U619 ( .A(KEYINPUT105), .ZN(n527) );
  XNOR2_X1 U620 ( .A(n542), .B(n527), .ZN(n528) );
  AND2_X1 U621 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U622 ( .A1(n538), .A2(n530), .ZN(n532) );
  INV_X1 U623 ( .A(KEYINPUT76), .ZN(n531) );
  INV_X1 U624 ( .A(n558), .ZN(n533) );
  NAND2_X1 U625 ( .A1(n533), .A2(n557), .ZN(n680) );
  INV_X1 U626 ( .A(n680), .ZN(n582) );
  NAND2_X1 U627 ( .A1(n591), .A2(n582), .ZN(n534) );
  XOR2_X1 U628 ( .A(n535), .B(n534), .Z(G30) );
  INV_X1 U629 ( .A(n537), .ZN(n686) );
  INV_X1 U630 ( .A(KEYINPUT107), .ZN(n539) );
  XNOR2_X1 U631 ( .A(n539), .B(KEYINPUT42), .ZN(n540) );
  XNOR2_X1 U632 ( .A(n570), .B(G137), .ZN(G39) );
  NAND2_X1 U633 ( .A1(n694), .A2(n693), .ZN(n541) );
  INV_X1 U634 ( .A(n555), .ZN(n543) );
  NAND2_X1 U635 ( .A1(n556), .A2(n684), .ZN(n545) );
  XOR2_X1 U636 ( .A(KEYINPUT30), .B(n545), .Z(n548) );
  INV_X1 U637 ( .A(n546), .ZN(n547) );
  AND2_X1 U638 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U639 ( .A(KEYINPUT66), .B(KEYINPUT39), .ZN(n550) );
  NAND2_X1 U640 ( .A1(n568), .A2(n582), .ZN(n607) );
  XNOR2_X1 U641 ( .A(n607), .B(G134), .ZN(G36) );
  INV_X1 U642 ( .A(n591), .ZN(n584) );
  INV_X1 U643 ( .A(n557), .ZN(n551) );
  NAND2_X1 U644 ( .A1(n551), .A2(n558), .ZN(n553) );
  INV_X1 U645 ( .A(KEYINPUT100), .ZN(n552) );
  XNOR2_X1 U646 ( .A(n553), .B(n552), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT101), .ZN(n676) );
  NOR2_X1 U648 ( .A1(n584), .A2(n676), .ZN(n554) );
  XOR2_X1 U649 ( .A(G146), .B(n554), .Z(G48) );
  INV_X1 U650 ( .A(n613), .ZN(n617) );
  OR2_X1 U651 ( .A1(n558), .A2(n557), .ZN(n592) );
  NAND2_X1 U652 ( .A1(n559), .A2(n422), .ZN(n562) );
  INV_X1 U653 ( .A(KEYINPUT73), .ZN(n560) );
  XNOR2_X1 U654 ( .A(n560), .B(KEYINPUT35), .ZN(n561) );
  XOR2_X1 U655 ( .A(n611), .B(G122), .Z(G24) );
  XNOR2_X1 U656 ( .A(n622), .B(KEYINPUT75), .ZN(n566) );
  INV_X1 U657 ( .A(n694), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U659 ( .A(n610), .B(G119), .ZN(G21) );
  NAND2_X1 U660 ( .A1(n568), .A2(n583), .ZN(n569) );
  XNOR2_X1 U661 ( .A(n569), .B(KEYINPUT40), .ZN(n658) );
  NAND2_X1 U662 ( .A1(n658), .A2(n570), .ZN(n572) );
  INV_X1 U663 ( .A(KEYINPUT46), .ZN(n571) );
  XNOR2_X1 U664 ( .A(n572), .B(n571), .ZN(n600) );
  XNOR2_X1 U665 ( .A(KEYINPUT102), .B(n574), .ZN(n575) );
  XNOR2_X1 U666 ( .A(KEYINPUT85), .B(KEYINPUT36), .ZN(n577) );
  XNOR2_X1 U667 ( .A(n578), .B(n577), .ZN(n579) );
  NAND2_X1 U668 ( .A1(n579), .A2(n563), .ZN(n581) );
  INV_X1 U669 ( .A(KEYINPUT108), .ZN(n580) );
  XNOR2_X1 U670 ( .A(n581), .B(n580), .ZN(n768) );
  OR2_X1 U671 ( .A1(n583), .A2(n582), .ZN(n619) );
  INV_X1 U672 ( .A(n619), .ZN(n683) );
  OR2_X1 U673 ( .A1(n584), .A2(n683), .ZN(n585) );
  NAND2_X1 U674 ( .A1(n585), .A2(KEYINPUT47), .ZN(n597) );
  OR2_X1 U675 ( .A1(n619), .A2(KEYINPUT78), .ZN(n589) );
  INV_X1 U676 ( .A(KEYINPUT78), .ZN(n586) );
  NOR2_X1 U677 ( .A1(n586), .A2(KEYINPUT47), .ZN(n587) );
  NAND2_X1 U678 ( .A1(n619), .A2(n587), .ZN(n588) );
  NAND2_X1 U679 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U680 ( .A1(n591), .A2(n590), .ZN(n595) );
  NOR2_X1 U681 ( .A1(n592), .A2(n576), .ZN(n593) );
  NAND2_X1 U682 ( .A1(n594), .A2(n593), .ZN(n675) );
  AND2_X1 U683 ( .A1(n595), .A2(n675), .ZN(n596) );
  NAND2_X1 U684 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U685 ( .A1(n768), .A2(n598), .ZN(n599) );
  NAND2_X1 U686 ( .A1(n600), .A2(n599), .ZN(n602) );
  NOR2_X1 U687 ( .A1(n563), .A2(n603), .ZN(n604) );
  XNOR2_X1 U688 ( .A(n604), .B(KEYINPUT43), .ZN(n605) );
  NOR2_X1 U689 ( .A1(n605), .A2(n383), .ZN(n606) );
  XNOR2_X1 U690 ( .A(n606), .B(KEYINPUT103), .ZN(n767) );
  NAND2_X1 U691 ( .A1(n612), .A2(n701), .ZN(n706) );
  OR2_X1 U692 ( .A1(n706), .A2(n613), .ZN(n615) );
  INV_X1 U693 ( .A(KEYINPUT31), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n615), .B(n614), .ZN(n679) );
  NOR2_X1 U695 ( .A1(n616), .A2(n701), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n670) );
  NAND2_X1 U697 ( .A1(n679), .A2(n670), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n619), .B(KEYINPUT78), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n622), .A2(n694), .ZN(n623) );
  NOR2_X1 U701 ( .A1(n623), .A2(n563), .ZN(n624) );
  AND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n667) );
  INV_X1 U703 ( .A(n667), .ZN(n626) );
  AND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n632), .A2(n630), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(KEYINPUT2), .ZN(n631) );
  INV_X1 U707 ( .A(KEYINPUT2), .ZN(n717) );
  NOR2_X1 U708 ( .A1(n633), .A2(n717), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n750), .A2(n634), .ZN(n724) );
  XNOR2_X1 U710 ( .A(n636), .B(KEYINPUT59), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(n640) );
  INV_X1 U712 ( .A(G952), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n641), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U714 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U717 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(G57) );
  XNOR2_X1 U719 ( .A(KEYINPUT86), .B(KEYINPUT54), .ZN(n650) );
  XNOR2_X1 U720 ( .A(KEYINPUT55), .B(KEYINPUT77), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U724 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n656) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(G51) );
  XNOR2_X1 U726 ( .A(G131), .B(KEYINPUT127), .ZN(n659) );
  XOR2_X1 U727 ( .A(n659), .B(n658), .Z(G33) );
  NAND2_X1 U728 ( .A1(n355), .A2(G469), .ZN(n665) );
  XNOR2_X1 U729 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n661) );
  XNOR2_X1 U730 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U734 ( .A1(n666), .A2(n742), .ZN(G54) );
  XOR2_X1 U735 ( .A(G101), .B(n667), .Z(G3) );
  NOR2_X1 U736 ( .A1(n676), .A2(n670), .ZN(n668) );
  XOR2_X1 U737 ( .A(KEYINPUT110), .B(n668), .Z(n669) );
  XNOR2_X1 U738 ( .A(G104), .B(n669), .ZN(G6) );
  NOR2_X1 U739 ( .A1(n670), .A2(n680), .ZN(n674) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n672) );
  XNOR2_X1 U741 ( .A(G107), .B(KEYINPUT26), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(G9) );
  XNOR2_X1 U744 ( .A(G143), .B(n675), .ZN(G45) );
  NOR2_X1 U745 ( .A1(n676), .A2(n679), .ZN(n677) );
  XOR2_X1 U746 ( .A(KEYINPUT112), .B(n677), .Z(n678) );
  XNOR2_X1 U747 ( .A(G113), .B(n678), .ZN(G15) );
  NOR2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U749 ( .A(G116), .B(n681), .Z(G18) );
  OR2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n690) );
  NOR2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U753 ( .A(n688), .B(KEYINPUT115), .ZN(n689) );
  NAND2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U755 ( .A1(n727), .A2(n691), .ZN(n692) );
  XOR2_X1 U756 ( .A(KEYINPUT116), .B(n692), .Z(n711) );
  NOR2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U758 ( .A(KEYINPUT49), .B(n695), .Z(n696) );
  XNOR2_X1 U759 ( .A(KEYINPUT113), .B(n696), .ZN(n704) );
  XOR2_X1 U760 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n700) );
  NAND2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U762 ( .A(n700), .B(n699), .ZN(n702) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U766 ( .A(KEYINPUT51), .B(n707), .ZN(n709) );
  INV_X1 U767 ( .A(n726), .ZN(n708) );
  NOR2_X1 U768 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U770 ( .A(n712), .B(KEYINPUT52), .ZN(n713) );
  NOR2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U772 ( .A(KEYINPUT117), .B(n715), .ZN(n733) );
  NAND2_X1 U773 ( .A1(n750), .A2(n759), .ZN(n718) );
  NAND2_X1 U774 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U775 ( .A1(n719), .A2(KEYINPUT80), .ZN(n723) );
  NOR2_X1 U776 ( .A1(KEYINPUT2), .A2(KEYINPUT80), .ZN(n720) );
  NAND2_X1 U777 ( .A1(n750), .A2(n720), .ZN(n721) );
  OR2_X1 U778 ( .A1(n721), .A2(n759), .ZN(n722) );
  NAND2_X1 U779 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U780 ( .A1(n725), .A2(n724), .ZN(n731) );
  NAND2_X1 U781 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U782 ( .A(KEYINPUT118), .B(n728), .Z(n729) );
  NOR2_X1 U783 ( .A1(n729), .A2(G953), .ZN(n730) );
  AND2_X1 U784 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U785 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U786 ( .A(KEYINPUT53), .B(n734), .Z(G75) );
  NAND2_X1 U787 ( .A1(n355), .A2(G478), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n735), .B(KEYINPUT121), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U790 ( .A1(n742), .A2(n738), .ZN(G63) );
  NAND2_X1 U791 ( .A1(n355), .A2(G217), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n742), .A2(n741), .ZN(G66) );
  XNOR2_X1 U794 ( .A(n743), .B(KEYINPUT125), .ZN(n745) );
  NAND2_X1 U795 ( .A1(n745), .A2(n744), .ZN(n755) );
  NAND2_X1 U796 ( .A1(G224), .A2(G953), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n746), .B(KEYINPUT122), .ZN(n747) );
  XNOR2_X1 U798 ( .A(KEYINPUT61), .B(n747), .ZN(n748) );
  NAND2_X1 U799 ( .A1(n748), .A2(G898), .ZN(n749) );
  XNOR2_X1 U800 ( .A(KEYINPUT123), .B(n749), .ZN(n753) );
  NAND2_X1 U801 ( .A1(n750), .A2(n760), .ZN(n751) );
  XOR2_X1 U802 ( .A(KEYINPUT124), .B(n751), .Z(n752) );
  NOR2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U804 ( .A(n755), .B(n754), .ZN(G69) );
  XNOR2_X1 U805 ( .A(n756), .B(KEYINPUT126), .ZN(n757) );
  XOR2_X1 U806 ( .A(n758), .B(n757), .Z(n762) );
  XOR2_X1 U807 ( .A(n762), .B(n759), .Z(n761) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(n766) );
  XNOR2_X1 U809 ( .A(G227), .B(n762), .ZN(n763) );
  NAND2_X1 U810 ( .A1(n763), .A2(G900), .ZN(n764) );
  NAND2_X1 U811 ( .A1(G953), .A2(n764), .ZN(n765) );
  NAND2_X1 U812 ( .A1(n766), .A2(n765), .ZN(G72) );
  XNOR2_X1 U813 ( .A(G140), .B(n767), .ZN(G42) );
  XNOR2_X1 U814 ( .A(G125), .B(KEYINPUT37), .ZN(n769) );
  XNOR2_X1 U815 ( .A(n769), .B(n768), .ZN(G27) );
endmodule

