

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U552 ( .A1(n530), .A2(G2104), .ZN(n887) );
  NOR2_X2 U553 ( .A1(G164), .A2(G1384), .ZN(n734) );
  NOR2_X2 U554 ( .A1(n542), .A2(n541), .ZN(G164) );
  XNOR2_X1 U555 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U556 ( .A(KEYINPUT103), .B(n831), .Z(n520) );
  NOR2_X1 U557 ( .A1(n809), .A2(n808), .ZN(n521) );
  INV_X1 U558 ( .A(KEYINPUT64), .ZN(n759) );
  XNOR2_X1 U559 ( .A(n740), .B(KEYINPUT99), .ZN(n741) );
  XNOR2_X1 U560 ( .A(n742), .B(n741), .ZN(n743) );
  AND2_X1 U561 ( .A1(G160), .A2(G40), .ZN(n735) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XNOR2_X1 U563 ( .A(KEYINPUT65), .B(KEYINPUT66), .ZN(n523) );
  NOR2_X1 U564 ( .A1(G651), .A2(n663), .ZN(n657) );
  AND2_X1 U565 ( .A1(G2104), .A2(G101), .ZN(n522) );
  NAND2_X1 U566 ( .A1(n522), .A2(n530), .ZN(n524) );
  XNOR2_X1 U567 ( .A(n525), .B(KEYINPUT23), .ZN(n527) );
  AND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NAND2_X1 U569 ( .A1(G113), .A2(n883), .ZN(n526) );
  NAND2_X1 U570 ( .A1(n527), .A2(n526), .ZN(n534) );
  XOR2_X1 U571 ( .A(KEYINPUT17), .B(n528), .Z(n529) );
  BUF_X2 U572 ( .A(n529), .Z(n888) );
  NAND2_X1 U573 ( .A1(G137), .A2(n888), .ZN(n532) );
  INV_X1 U574 ( .A(G2105), .ZN(n530) );
  NOR2_X4 U575 ( .A1(G2104), .A2(n530), .ZN(n884) );
  NAND2_X1 U576 ( .A1(G125), .A2(n884), .ZN(n531) );
  NAND2_X1 U577 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X2 U578 ( .A1(n534), .A2(n533), .ZN(G160) );
  NAND2_X1 U579 ( .A1(G102), .A2(n887), .ZN(n535) );
  XNOR2_X1 U580 ( .A(n535), .B(KEYINPUT88), .ZN(n538) );
  NAND2_X1 U581 ( .A1(G126), .A2(n884), .ZN(n536) );
  XOR2_X1 U582 ( .A(KEYINPUT87), .B(n536), .Z(n537) );
  NAND2_X1 U583 ( .A1(n538), .A2(n537), .ZN(n542) );
  NAND2_X1 U584 ( .A1(G114), .A2(n883), .ZN(n540) );
  NAND2_X1 U585 ( .A1(G138), .A2(n888), .ZN(n539) );
  NAND2_X1 U586 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U587 ( .A(G2443), .B(G2446), .Z(n544) );
  XNOR2_X1 U588 ( .A(G2427), .B(G2451), .ZN(n543) );
  XNOR2_X1 U589 ( .A(n544), .B(n543), .ZN(n550) );
  XOR2_X1 U590 ( .A(G2430), .B(G2454), .Z(n546) );
  XNOR2_X1 U591 ( .A(G1348), .B(G1341), .ZN(n545) );
  XNOR2_X1 U592 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U593 ( .A(G2435), .B(G2438), .Z(n547) );
  XNOR2_X1 U594 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U595 ( .A(n550), .B(n549), .Z(n551) );
  AND2_X1 U596 ( .A1(G14), .A2(n551), .ZN(G401) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U598 ( .A1(G99), .A2(n887), .ZN(n552) );
  XNOR2_X1 U599 ( .A(n552), .B(KEYINPUT74), .ZN(n556) );
  XOR2_X1 U600 ( .A(KEYINPUT18), .B(KEYINPUT73), .Z(n554) );
  NAND2_X1 U601 ( .A1(G123), .A2(n884), .ZN(n553) );
  XNOR2_X1 U602 ( .A(n554), .B(n553), .ZN(n555) );
  NAND2_X1 U603 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U604 ( .A1(G111), .A2(n883), .ZN(n558) );
  NAND2_X1 U605 ( .A1(G135), .A2(n888), .ZN(n557) );
  NAND2_X1 U606 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U607 ( .A1(n560), .A2(n559), .ZN(n1003) );
  XNOR2_X1 U608 ( .A(n1003), .B(G2096), .ZN(n561) );
  XNOR2_X1 U609 ( .A(n561), .B(KEYINPUT75), .ZN(n562) );
  OR2_X1 U610 ( .A1(G2100), .A2(n562), .ZN(G156) );
  INV_X1 U611 ( .A(G651), .ZN(n567) );
  NOR2_X1 U612 ( .A1(G543), .A2(n567), .ZN(n564) );
  XNOR2_X1 U613 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n563) );
  XNOR2_X1 U614 ( .A(n564), .B(n563), .ZN(n661) );
  NAND2_X1 U615 ( .A1(G65), .A2(n661), .ZN(n566) );
  XOR2_X1 U616 ( .A(KEYINPUT0), .B(G543), .Z(n663) );
  NAND2_X1 U617 ( .A1(G53), .A2(n657), .ZN(n565) );
  NAND2_X1 U618 ( .A1(n566), .A2(n565), .ZN(n571) );
  NOR2_X1 U619 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U620 ( .A1(G91), .A2(n645), .ZN(n569) );
  NOR2_X1 U621 ( .A1(n663), .A2(n567), .ZN(n650) );
  NAND2_X1 U622 ( .A1(G78), .A2(n650), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U624 ( .A1(n571), .A2(n570), .ZN(n771) );
  INV_X1 U625 ( .A(n771), .ZN(G299) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  NAND2_X1 U627 ( .A1(G64), .A2(n661), .ZN(n573) );
  NAND2_X1 U628 ( .A1(G52), .A2(n657), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n573), .A2(n572), .ZN(n580) );
  NAND2_X1 U630 ( .A1(n645), .A2(G90), .ZN(n574) );
  XNOR2_X1 U631 ( .A(KEYINPUT69), .B(n574), .ZN(n577) );
  NAND2_X1 U632 ( .A1(n650), .A2(G77), .ZN(n575) );
  XOR2_X1 U633 ( .A(KEYINPUT70), .B(n575), .Z(n576) );
  NOR2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U635 ( .A(n578), .B(KEYINPUT9), .ZN(n579) );
  NOR2_X1 U636 ( .A1(n580), .A2(n579), .ZN(G171) );
  INV_X1 U637 ( .A(G171), .ZN(G301) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U639 ( .A(n581), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U640 ( .A(G223), .ZN(n834) );
  NAND2_X1 U641 ( .A1(n834), .A2(G567), .ZN(n582) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  NAND2_X1 U643 ( .A1(G56), .A2(n661), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(n583), .Z(n589) );
  NAND2_X1 U645 ( .A1(n645), .A2(G81), .ZN(n584) );
  XNOR2_X1 U646 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G68), .A2(n650), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U649 ( .A(KEYINPUT13), .B(n587), .Z(n588) );
  NOR2_X1 U650 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U651 ( .A1(n657), .A2(G43), .ZN(n590) );
  NAND2_X1 U652 ( .A1(n591), .A2(n590), .ZN(n949) );
  INV_X1 U653 ( .A(G860), .ZN(n616) );
  OR2_X1 U654 ( .A1(n949), .A2(n616), .ZN(G153) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U656 ( .A1(G66), .A2(n661), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G92), .A2(n645), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U659 ( .A1(G79), .A2(n650), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G54), .A2(n657), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n598), .Z(n622) );
  INV_X1 U664 ( .A(n622), .ZN(n948) );
  INV_X1 U665 ( .A(G868), .ZN(n612) );
  NAND2_X1 U666 ( .A1(n948), .A2(n612), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U668 ( .A1(n645), .A2(G89), .ZN(n601) );
  XNOR2_X1 U669 ( .A(n601), .B(KEYINPUT4), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G76), .A2(n650), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U672 ( .A(KEYINPUT5), .B(n604), .ZN(n610) );
  NAND2_X1 U673 ( .A1(n657), .A2(G51), .ZN(n605) );
  XOR2_X1 U674 ( .A(KEYINPUT71), .B(n605), .Z(n607) );
  NAND2_X1 U675 ( .A1(n661), .A2(G63), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U677 ( .A(KEYINPUT6), .B(n608), .Z(n609) );
  NAND2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U679 ( .A(KEYINPUT7), .B(n611), .ZN(G168) );
  XOR2_X1 U680 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U681 ( .A1(G286), .A2(n612), .ZN(n614) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n613) );
  NOR2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U684 ( .A(KEYINPUT72), .B(n615), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n616), .A2(G559), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n617), .A2(n622), .ZN(n618) );
  XNOR2_X1 U687 ( .A(n618), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G868), .A2(n949), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n622), .A2(G868), .ZN(n619) );
  NOR2_X1 U690 ( .A1(G559), .A2(n619), .ZN(n620) );
  NOR2_X1 U691 ( .A1(n621), .A2(n620), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G559), .A2(n622), .ZN(n623) );
  XNOR2_X1 U693 ( .A(n949), .B(n623), .ZN(n676) );
  NOR2_X1 U694 ( .A1(n676), .A2(G860), .ZN(n630) );
  NAND2_X1 U695 ( .A1(G67), .A2(n661), .ZN(n625) );
  NAND2_X1 U696 ( .A1(G55), .A2(n657), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U698 ( .A1(G93), .A2(n645), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G80), .A2(n650), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U701 ( .A1(n629), .A2(n628), .ZN(n670) );
  XNOR2_X1 U702 ( .A(n630), .B(n670), .ZN(G145) );
  NAND2_X1 U703 ( .A1(G62), .A2(n661), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G50), .A2(n657), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U706 ( .A(KEYINPUT81), .B(n633), .ZN(n637) );
  NAND2_X1 U707 ( .A1(G88), .A2(n645), .ZN(n635) );
  NAND2_X1 U708 ( .A1(G75), .A2(n650), .ZN(n634) );
  AND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n637), .A2(n636), .ZN(G303) );
  INV_X1 U711 ( .A(G303), .ZN(G166) );
  NAND2_X1 U712 ( .A1(n645), .A2(G85), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n661), .A2(G60), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U715 ( .A1(G72), .A2(n650), .ZN(n641) );
  NAND2_X1 U716 ( .A1(G47), .A2(n657), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U719 ( .A(KEYINPUT68), .B(n644), .Z(G290) );
  NAND2_X1 U720 ( .A1(n645), .A2(G86), .ZN(n646) );
  XNOR2_X1 U721 ( .A(n646), .B(KEYINPUT78), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G61), .A2(n661), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U724 ( .A(KEYINPUT79), .B(n649), .ZN(n656) );
  NAND2_X1 U725 ( .A1(G73), .A2(n650), .ZN(n651) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n651), .Z(n654) );
  NAND2_X1 U727 ( .A1(n657), .A2(G48), .ZN(n652) );
  XOR2_X1 U728 ( .A(KEYINPUT80), .B(n652), .Z(n653) );
  NOR2_X1 U729 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(G305) );
  NAND2_X1 U731 ( .A1(G49), .A2(n657), .ZN(n659) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n662), .B(KEYINPUT76), .ZN(n665) );
  NAND2_X1 U736 ( .A1(G87), .A2(n663), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U738 ( .A(KEYINPUT77), .B(n666), .Z(G288) );
  NOR2_X1 U739 ( .A1(G868), .A2(n670), .ZN(n667) );
  XOR2_X1 U740 ( .A(n667), .B(KEYINPUT84), .Z(n679) );
  XOR2_X1 U741 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n669) );
  XNOR2_X1 U742 ( .A(G166), .B(KEYINPUT82), .ZN(n668) );
  XNOR2_X1 U743 ( .A(n669), .B(n668), .ZN(n671) );
  XOR2_X1 U744 ( .A(n671), .B(n670), .Z(n673) );
  XNOR2_X1 U745 ( .A(G290), .B(n771), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U747 ( .A(n674), .B(G305), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n675), .B(G288), .ZN(n903) );
  XOR2_X1 U749 ( .A(n903), .B(n676), .Z(n677) );
  NAND2_X1 U750 ( .A1(G868), .A2(n677), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2084), .A2(G2078), .ZN(n680) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n681), .ZN(n683) );
  XOR2_X1 U755 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n682) );
  XNOR2_X1 U756 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U757 ( .A1(G2072), .A2(n684), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U759 ( .A1(G132), .A2(G82), .ZN(n685) );
  XNOR2_X1 U760 ( .A(n685), .B(KEYINPUT22), .ZN(n686) );
  XNOR2_X1 U761 ( .A(n686), .B(KEYINPUT86), .ZN(n687) );
  NOR2_X1 U762 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U763 ( .A1(G96), .A2(n688), .ZN(n838) );
  NAND2_X1 U764 ( .A1(n838), .A2(G2106), .ZN(n692) );
  NAND2_X1 U765 ( .A1(G108), .A2(G120), .ZN(n689) );
  NOR2_X1 U766 ( .A1(G237), .A2(n689), .ZN(n690) );
  NAND2_X1 U767 ( .A1(G69), .A2(n690), .ZN(n839) );
  NAND2_X1 U768 ( .A1(n839), .A2(G567), .ZN(n691) );
  NAND2_X1 U769 ( .A1(n692), .A2(n691), .ZN(n840) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n693) );
  NOR2_X1 U771 ( .A1(n840), .A2(n693), .ZN(n837) );
  NAND2_X1 U772 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U773 ( .A1(G117), .A2(n883), .ZN(n695) );
  NAND2_X1 U774 ( .A1(G129), .A2(n884), .ZN(n694) );
  NAND2_X1 U775 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U776 ( .A1(n887), .A2(G105), .ZN(n696) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n696), .Z(n697) );
  NOR2_X1 U778 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U779 ( .A1(n888), .A2(G141), .ZN(n699) );
  NAND2_X1 U780 ( .A1(n700), .A2(n699), .ZN(n899) );
  NOR2_X1 U781 ( .A1(G1996), .A2(n899), .ZN(n1000) );
  NAND2_X1 U782 ( .A1(G107), .A2(n883), .ZN(n702) );
  NAND2_X1 U783 ( .A1(G131), .A2(n888), .ZN(n701) );
  NAND2_X1 U784 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U785 ( .A1(G95), .A2(n887), .ZN(n704) );
  NAND2_X1 U786 ( .A1(G119), .A2(n884), .ZN(n703) );
  NAND2_X1 U787 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U788 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U789 ( .A(n707), .B(KEYINPUT91), .ZN(n877) );
  NOR2_X1 U790 ( .A1(G1991), .A2(n877), .ZN(n1002) );
  NOR2_X1 U791 ( .A1(G290), .A2(G1986), .ZN(n708) );
  XNOR2_X1 U792 ( .A(KEYINPUT104), .B(n708), .ZN(n709) );
  NOR2_X1 U793 ( .A1(n1002), .A2(n709), .ZN(n712) );
  NAND2_X1 U794 ( .A1(G1991), .A2(n877), .ZN(n711) );
  NAND2_X1 U795 ( .A1(G1996), .A2(n899), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n711), .A2(n710), .ZN(n730) );
  NOR2_X1 U797 ( .A1(n712), .A2(n730), .ZN(n713) );
  NOR2_X1 U798 ( .A1(n1000), .A2(n713), .ZN(n714) );
  XNOR2_X1 U799 ( .A(KEYINPUT39), .B(n714), .ZN(n725) );
  NAND2_X1 U800 ( .A1(G116), .A2(n883), .ZN(n716) );
  NAND2_X1 U801 ( .A1(G128), .A2(n884), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U803 ( .A(n717), .B(KEYINPUT35), .ZN(n722) );
  NAND2_X1 U804 ( .A1(G104), .A2(n887), .ZN(n719) );
  NAND2_X1 U805 ( .A1(G140), .A2(n888), .ZN(n718) );
  NAND2_X1 U806 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U807 ( .A(KEYINPUT34), .B(n720), .Z(n721) );
  NAND2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U809 ( .A(n723), .B(KEYINPUT36), .Z(n878) );
  XOR2_X1 U810 ( .A(G2067), .B(KEYINPUT37), .Z(n724) );
  XOR2_X1 U811 ( .A(KEYINPUT90), .B(n724), .Z(n726) );
  OR2_X1 U812 ( .A1(n878), .A2(n726), .ZN(n731) );
  NAND2_X1 U813 ( .A1(n725), .A2(n731), .ZN(n727) );
  NAND2_X1 U814 ( .A1(n726), .A2(n878), .ZN(n1011) );
  NAND2_X1 U815 ( .A1(n727), .A2(n1011), .ZN(n729) );
  NAND2_X1 U816 ( .A1(G160), .A2(G40), .ZN(n728) );
  NOR2_X1 U817 ( .A1(n734), .A2(n728), .ZN(n825) );
  NAND2_X1 U818 ( .A1(n729), .A2(n825), .ZN(n832) );
  INV_X1 U819 ( .A(n730), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n1013) );
  NAND2_X1 U821 ( .A1(n825), .A2(n1013), .ZN(n733) );
  XNOR2_X1 U822 ( .A(KEYINPUT92), .B(n733), .ZN(n830) );
  NAND2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n789) );
  NAND2_X1 U824 ( .A1(n789), .A2(G8), .ZN(n736) );
  XNOR2_X1 U825 ( .A(n736), .B(KEYINPUT93), .ZN(n737) );
  BUF_X1 U826 ( .A(n737), .Z(n819) );
  NOR2_X1 U827 ( .A1(G2084), .A2(n789), .ZN(n738) );
  NAND2_X1 U828 ( .A1(G8), .A2(n738), .ZN(n788) );
  INV_X1 U829 ( .A(n737), .ZN(n809) );
  NOR2_X1 U830 ( .A1(G1966), .A2(n809), .ZN(n785) );
  NOR2_X1 U831 ( .A1(n738), .A2(n785), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n739), .A2(G8), .ZN(n742) );
  INV_X1 U833 ( .A(KEYINPUT30), .ZN(n740) );
  NOR2_X1 U834 ( .A1(n743), .A2(G168), .ZN(n745) );
  INV_X1 U835 ( .A(KEYINPUT100), .ZN(n744) );
  XNOR2_X1 U836 ( .A(n745), .B(n744), .ZN(n749) );
  XOR2_X1 U837 ( .A(G2078), .B(KEYINPUT25), .Z(n924) );
  NOR2_X1 U838 ( .A1(n924), .A2(n789), .ZN(n747) );
  INV_X1 U839 ( .A(n789), .ZN(n754) );
  NOR2_X1 U840 ( .A1(n754), .A2(G1961), .ZN(n746) );
  NOR2_X1 U841 ( .A1(n747), .A2(n746), .ZN(n779) );
  NAND2_X1 U842 ( .A1(n779), .A2(G301), .ZN(n748) );
  NAND2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U844 ( .A(n750), .B(KEYINPUT31), .ZN(n783) );
  NAND2_X1 U845 ( .A1(n754), .A2(G2067), .ZN(n752) );
  NAND2_X1 U846 ( .A1(G1348), .A2(n789), .ZN(n751) );
  NAND2_X1 U847 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U848 ( .A(n753), .B(KEYINPUT97), .Z(n761) );
  NAND2_X1 U849 ( .A1(n948), .A2(n761), .ZN(n765) );
  AND2_X1 U850 ( .A1(n754), .A2(G1996), .ZN(n755) );
  XOR2_X1 U851 ( .A(n755), .B(KEYINPUT26), .Z(n757) );
  NAND2_X1 U852 ( .A1(n789), .A2(G1341), .ZN(n756) );
  NAND2_X1 U853 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U854 ( .A1(n949), .A2(n758), .ZN(n760) );
  XNOR2_X1 U855 ( .A(n760), .B(n759), .ZN(n763) );
  OR2_X1 U856 ( .A1(n948), .A2(n761), .ZN(n762) );
  NAND2_X1 U857 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n754), .A2(G2072), .ZN(n766) );
  XNOR2_X1 U860 ( .A(n766), .B(KEYINPUT27), .ZN(n768) );
  XNOR2_X1 U861 ( .A(G1956), .B(KEYINPUT95), .ZN(n961) );
  NOR2_X1 U862 ( .A1(n961), .A2(n754), .ZN(n767) );
  NOR2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n769) );
  NAND2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n776) );
  NOR2_X1 U866 ( .A1(n772), .A2(n771), .ZN(n774) );
  XOR2_X1 U867 ( .A(KEYINPUT96), .B(KEYINPUT28), .Z(n773) );
  XNOR2_X1 U868 ( .A(n774), .B(n773), .ZN(n775) );
  NAND2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n778) );
  XOR2_X1 U870 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n777) );
  XNOR2_X1 U871 ( .A(n778), .B(n777), .ZN(n781) );
  OR2_X1 U872 ( .A1(n779), .A2(G301), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n793) );
  INV_X1 U875 ( .A(n793), .ZN(n784) );
  NOR2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U877 ( .A(KEYINPUT101), .B(n786), .Z(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n799) );
  NOR2_X1 U879 ( .A1(G1971), .A2(n809), .ZN(n791) );
  NOR2_X1 U880 ( .A1(G2090), .A2(n789), .ZN(n790) );
  NOR2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n792), .A2(G303), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G286), .A2(n793), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G8), .A2(n796), .ZN(n797) );
  XNOR2_X1 U886 ( .A(KEYINPUT32), .B(n797), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n807) );
  NOR2_X1 U888 ( .A1(G2090), .A2(G303), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G8), .A2(n800), .ZN(n801) );
  AND2_X1 U890 ( .A1(n807), .A2(n801), .ZN(n802) );
  XNOR2_X1 U891 ( .A(n802), .B(KEYINPUT102), .ZN(n803) );
  NOR2_X1 U892 ( .A1(n819), .A2(n803), .ZN(n824) );
  NOR2_X1 U893 ( .A1(G1976), .A2(G288), .ZN(n812) );
  NOR2_X1 U894 ( .A1(G1971), .A2(G303), .ZN(n804) );
  NOR2_X1 U895 ( .A1(n812), .A2(n804), .ZN(n942) );
  INV_X1 U896 ( .A(KEYINPUT33), .ZN(n805) );
  AND2_X1 U897 ( .A1(n942), .A2(n805), .ZN(n806) );
  NAND2_X1 U898 ( .A1(n807), .A2(n806), .ZN(n811) );
  NAND2_X1 U899 ( .A1(G1976), .A2(G288), .ZN(n946) );
  INV_X1 U900 ( .A(n946), .ZN(n808) );
  OR2_X1 U901 ( .A1(KEYINPUT33), .A2(n521), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n816) );
  AND2_X1 U903 ( .A1(n812), .A2(KEYINPUT33), .ZN(n813) );
  AND2_X1 U904 ( .A1(n813), .A2(n819), .ZN(n814) );
  XNOR2_X1 U905 ( .A(G1981), .B(G305), .ZN(n936) );
  OR2_X1 U906 ( .A1(n814), .A2(n936), .ZN(n815) );
  OR2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n822) );
  NOR2_X1 U908 ( .A1(G1981), .A2(G305), .ZN(n817) );
  XNOR2_X1 U909 ( .A(n817), .B(KEYINPUT24), .ZN(n818) );
  XNOR2_X1 U910 ( .A(n818), .B(KEYINPUT94), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U912 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U913 ( .A1(n824), .A2(n823), .ZN(n828) );
  XNOR2_X1 U914 ( .A(G290), .B(G1986), .ZN(n944) );
  NAND2_X1 U915 ( .A1(n825), .A2(n944), .ZN(n826) );
  XNOR2_X1 U916 ( .A(n826), .B(KEYINPUT89), .ZN(n827) );
  NOR2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U918 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U919 ( .A1(n832), .A2(n520), .ZN(n833) );
  XNOR2_X1 U920 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U923 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U925 ( .A1(n837), .A2(n836), .ZN(G188) );
  XNOR2_X1 U926 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G108), .ZN(G238) );
  INV_X1 U930 ( .A(G82), .ZN(G220) );
  NOR2_X1 U931 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n840), .ZN(G319) );
  XOR2_X1 U934 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n842) );
  XNOR2_X1 U935 ( .A(G2678), .B(KEYINPUT43), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U937 ( .A(KEYINPUT42), .B(G2090), .Z(n844) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U940 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U941 ( .A(G2096), .B(G2100), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n848), .B(n847), .ZN(n850) );
  XOR2_X1 U943 ( .A(G2084), .B(G2078), .Z(n849) );
  XNOR2_X1 U944 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1976), .B(G1971), .Z(n852) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1956), .ZN(n851) );
  XNOR2_X1 U947 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U948 ( .A(n853), .B(G2474), .Z(n855) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1981), .Z(n857) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1961), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U955 ( .A1(n884), .A2(G124), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U957 ( .A1(G136), .A2(n888), .ZN(n861) );
  NAND2_X1 U958 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U959 ( .A(KEYINPUT108), .B(n863), .ZN(n867) );
  NAND2_X1 U960 ( .A1(G100), .A2(n887), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G112), .A2(n883), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U963 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U964 ( .A1(G103), .A2(n887), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G139), .A2(n888), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n874) );
  NAND2_X1 U967 ( .A1(G115), .A2(n883), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G127), .A2(n884), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U972 ( .A(KEYINPUT110), .B(n875), .ZN(n994) );
  XOR2_X1 U973 ( .A(G164), .B(n1003), .Z(n876) );
  XNOR2_X1 U974 ( .A(n994), .B(n876), .ZN(n882) );
  XNOR2_X1 U975 ( .A(n877), .B(G162), .ZN(n880) );
  XOR2_X1 U976 ( .A(G160), .B(n878), .Z(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n882), .B(n881), .ZN(n901) );
  XOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n897) );
  NAND2_X1 U980 ( .A1(G118), .A2(n883), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G130), .A2(n884), .ZN(n885) );
  NAND2_X1 U982 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U983 ( .A1(G106), .A2(n887), .ZN(n890) );
  NAND2_X1 U984 ( .A1(G142), .A2(n888), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U986 ( .A(KEYINPUT109), .B(n891), .ZN(n892) );
  XNOR2_X1 U987 ( .A(KEYINPUT45), .B(n892), .ZN(n893) );
  NOR2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U989 ( .A(KEYINPUT111), .B(n895), .ZN(n896) );
  XNOR2_X1 U990 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U991 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U992 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U993 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U994 ( .A(n903), .B(KEYINPUT112), .ZN(n905) );
  XNOR2_X1 U995 ( .A(n949), .B(G286), .ZN(n904) );
  XNOR2_X1 U996 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U997 ( .A(n948), .B(G171), .Z(n906) );
  XNOR2_X1 U998 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U999 ( .A1(G37), .A2(n908), .ZN(G397) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1001 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n910), .B(n909), .ZN(n913) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(n911), .B(KEYINPUT114), .ZN(n912) );
  NAND2_X1 U1005 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n914), .ZN(n915) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n915), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G96), .ZN(G221) );
  INV_X1 U1010 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1011 ( .A(G1996), .B(G32), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(G1991), .B(G25), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n923) );
  XOR2_X1 U1014 ( .A(G2072), .B(G33), .Z(n918) );
  NAND2_X1 U1015 ( .A1(n918), .A2(G28), .ZN(n921) );
  XOR2_X1 U1016 ( .A(KEYINPUT119), .B(G2067), .Z(n919) );
  XNOR2_X1 U1017 ( .A(G26), .B(n919), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(G27), .B(n924), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1022 ( .A(KEYINPUT53), .B(n927), .Z(n930) );
  XOR2_X1 U1023 ( .A(G34), .B(KEYINPUT54), .Z(n928) );
  XNOR2_X1 U1024 ( .A(G2084), .B(n928), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(G35), .B(G2090), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1028 ( .A(KEYINPUT55), .B(n933), .Z(n934) );
  NOR2_X1 U1029 ( .A1(G29), .A2(n934), .ZN(n991) );
  XNOR2_X1 U1030 ( .A(G16), .B(KEYINPUT56), .ZN(n959) );
  XOR2_X1 U1031 ( .A(G168), .B(G1966), .Z(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1033 ( .A(KEYINPUT57), .B(n937), .Z(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT120), .B(n938), .ZN(n957) );
  XNOR2_X1 U1035 ( .A(G299), .B(G1956), .ZN(n940) );
  AND2_X1 U1036 ( .A1(G1971), .A2(G303), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(n947), .B(KEYINPUT121), .ZN(n953) );
  XNOR2_X1 U1042 ( .A(n948), .B(G1348), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(n949), .B(G1341), .ZN(n950) );
  NOR2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(G1961), .B(G301), .ZN(n954) );
  NOR2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1049 ( .A1(n959), .A2(n958), .ZN(n988) );
  INV_X1 U1050 ( .A(G16), .ZN(n986) );
  XOR2_X1 U1051 ( .A(G1348), .B(KEYINPUT59), .Z(n960) );
  XNOR2_X1 U1052 ( .A(G4), .B(n960), .ZN(n969) );
  XNOR2_X1 U1053 ( .A(G20), .B(n961), .ZN(n964) );
  XOR2_X1 U1054 ( .A(G1981), .B(KEYINPUT122), .Z(n962) );
  XNOR2_X1 U1055 ( .A(G6), .B(n962), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(G19), .B(G1341), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(n967), .B(KEYINPUT123), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(KEYINPUT124), .B(n970), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n971), .B(KEYINPUT60), .ZN(n975) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G21), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(G5), .B(G1961), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n982) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G23), .B(G1976), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n979) );
  XOR2_X1 U1070 ( .A(G1986), .B(G24), .Z(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(KEYINPUT58), .B(n980), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1074 ( .A(n983), .B(KEYINPUT61), .Z(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(n984), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n989), .B(KEYINPUT126), .ZN(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(G11), .A2(n992), .ZN(n993) );
  XOR2_X1 U1081 ( .A(KEYINPUT127), .B(n993), .Z(n1023) );
  XNOR2_X1 U1082 ( .A(G164), .B(G2078), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(G2072), .B(KEYINPUT116), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(n998), .B(KEYINPUT50), .ZN(n1010) );
  XOR2_X1 U1087 ( .A(G2090), .B(G162), .Z(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(KEYINPUT51), .B(n1001), .Z(n1008) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(n1004), .B(KEYINPUT115), .ZN(n1006) );
  XOR2_X1 U1092 ( .A(G160), .B(G2084), .Z(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1015) );
  INV_X1 U1096 ( .A(n1011), .ZN(n1012) );
  NOR2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1098 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(KEYINPUT52), .B(n1016), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(KEYINPUT117), .B(n1017), .ZN(n1019) );
  INV_X1 U1101 ( .A(KEYINPUT55), .ZN(n1018) );
  NAND2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1103 ( .A1(n1020), .A2(G29), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(KEYINPUT118), .B(n1021), .Z(n1022) );
  NOR2_X1 U1105 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1024), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

