//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n187), .A2(new_n188), .A3(G953), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT89), .B1(new_n191), .B2(G143), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT89), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(G128), .B2(new_n194), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G134), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n196), .B(new_n199), .C1(G128), .C2(new_n194), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G116), .B(G122), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT92), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(KEYINPUT92), .A3(new_n203), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT14), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n210), .A2(G122), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n203), .B1(new_n211), .B2(KEYINPUT14), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n206), .A2(new_n207), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n201), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT93), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n201), .A2(new_n213), .A3(KEYINPUT93), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n202), .A2(new_n203), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n204), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT88), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(KEYINPUT88), .A3(new_n204), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n200), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT13), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n196), .A2(new_n225), .B1(new_n191), .B2(G143), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT90), .B1(new_n196), .B2(new_n225), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n192), .A2(new_n195), .A3(new_n228), .A4(KEYINPUT13), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G134), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT91), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT91), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n233), .A3(G134), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n224), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n190), .B1(new_n218), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n216), .A2(new_n217), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n232), .A2(new_n234), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n237), .B(new_n189), .C1(new_n238), .C2(new_n224), .ZN(new_n239));
  AOI21_X1  g053(.A(G902), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G478), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(KEYINPUT15), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n240), .B(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G952), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G953), .ZN(new_n245));
  NAND2_X1  g059(.A1(G234), .A2(G237), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n246), .A2(G902), .A3(G953), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT21), .B(G898), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G113), .B(G122), .ZN(new_n253));
  INV_X1    g067(.A(G104), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G237), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(G214), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n194), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT83), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n262), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G131), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT17), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT83), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n259), .A2(new_n268), .A3(new_n260), .A4(new_n262), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n264), .A2(new_n266), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT16), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G125), .ZN(new_n274));
  INV_X1    g088(.A(G125), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(KEYINPUT71), .ZN(new_n276));
  OAI21_X1  g090(.A(G140), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(G125), .A2(G140), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n272), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT16), .A2(G140), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n275), .A2(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n273), .A2(G125), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n271), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G140), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n283), .B2(new_n284), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT16), .B1(new_n288), .B2(new_n278), .ZN(new_n289));
  INV_X1    g103(.A(new_n285), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(G146), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n265), .A2(KEYINPUT17), .A3(G131), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n270), .A2(new_n286), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT18), .A2(G131), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n265), .B(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(G125), .B(G140), .Z(new_n296));
  OR2_X1    g110(.A1(new_n296), .A2(G146), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT71), .B(G125), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n279), .B1(new_n298), .B2(new_n287), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n299), .B2(new_n271), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n255), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n255), .B(KEYINPUT85), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n293), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n293), .A2(new_n301), .A3(KEYINPUT86), .A4(new_n303), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n302), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G475), .B1(new_n308), .B2(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n307), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n264), .A2(new_n266), .A3(new_n269), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT19), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n313));
  OAI22_X1  g127(.A1(new_n299), .A2(new_n312), .B1(new_n296), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n311), .B(new_n291), .C1(G146), .C2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n255), .B1(new_n315), .B2(new_n301), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT20), .ZN(new_n319));
  NOR2_X1   g133(.A1(G475), .A2(G902), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n318), .A2(KEYINPUT87), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n316), .B1(new_n306), .B2(new_n307), .ZN(new_n322));
  INV_X1    g136(.A(new_n320), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT20), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n322), .A2(new_n323), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT87), .B1(new_n326), .B2(new_n319), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n309), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n252), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G469), .ZN(new_n332));
  INV_X1    g146(.A(G902), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n194), .A2(KEYINPUT1), .A3(G146), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n271), .A2(G143), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n194), .A2(G146), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n335), .B1(new_n338), .B2(new_n191), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n336), .A3(new_n337), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G143), .B(G146), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(KEYINPUT76), .A3(new_n340), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(new_n254), .B2(G107), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n203), .A3(G104), .ZN(new_n349));
  INV_X1    g163(.A(G101), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n254), .A2(G107), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n347), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n254), .A2(G107), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n203), .A2(G104), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n346), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT11), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n199), .B2(G137), .ZN(new_n361));
  INV_X1    g175(.A(G137), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT11), .A3(G134), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n199), .A2(G137), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(KEYINPUT66), .A2(G131), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n361), .A2(new_n363), .A3(new_n366), .A4(new_n364), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT0), .A2(G128), .ZN(new_n372));
  NOR3_X1   g186(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n344), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n338), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G101), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n379), .A2(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n378), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n358), .B1(new_n339), .B2(new_n341), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n356), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n359), .A2(new_n371), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n357), .A2(new_n358), .B1(new_n356), .B2(new_n385), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n371), .A4(new_n384), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n338), .A2(new_n191), .ZN(new_n393));
  INV_X1    g207(.A(new_n335), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n393), .A2(new_n394), .A3(new_n341), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n352), .A2(new_n355), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n357), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n370), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT12), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(KEYINPUT12), .A3(new_n370), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n392), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n257), .A2(G227), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT75), .ZN(new_n406));
  XNOR2_X1  g220(.A(G110), .B(G140), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n388), .B2(new_n391), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n389), .A2(new_n384), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n370), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n404), .A2(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n334), .B1(new_n412), .B2(G469), .ZN(new_n413));
  INV_X1    g227(.A(new_n408), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n392), .A2(new_n414), .A3(new_n403), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n388), .A2(new_n391), .B1(new_n370), .B2(new_n410), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n415), .B1(new_n416), .B2(new_n414), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n332), .A3(new_n333), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n331), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n298), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n378), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n394), .B(new_n341), .C1(G128), .C2(new_n344), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n298), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n257), .A2(G224), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n424), .B(KEYINPUT79), .Z(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT7), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT80), .ZN(new_n428));
  INV_X1    g242(.A(new_n426), .ZN(new_n429));
  INV_X1    g243(.A(new_n423), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n298), .B1(new_n374), .B2(new_n377), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT80), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n421), .A2(new_n433), .A3(new_n423), .A4(new_n426), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n428), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(G110), .B(G122), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT8), .ZN(new_n437));
  OR2_X1    g251(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n438));
  INV_X1    g252(.A(G119), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n438), .A2(G116), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(G116), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n210), .A2(G119), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT5), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n441), .A2(G113), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n443), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT2), .B(G113), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n445), .A2(new_n396), .A3(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n438), .A2(new_n440), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n441), .B(G113), .C1(new_n450), .C2(new_n446), .ZN(new_n451));
  INV_X1    g265(.A(new_n448), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n451), .A2(new_n452), .B1(new_n352), .B2(new_n355), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n437), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n356), .A2(new_n451), .A3(new_n452), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n446), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n447), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n447), .B1(new_n456), .B2(new_n446), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n381), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n382), .A2(new_n383), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n436), .B(new_n455), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n454), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n435), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G210), .B1(G237), .B2(G902), .ZN(new_n466));
  XOR2_X1   g280(.A(new_n466), .B(KEYINPUT81), .Z(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n455), .B1(new_n461), .B2(new_n462), .ZN(new_n469));
  INV_X1    g283(.A(new_n436), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n463), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n473), .A3(new_n470), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n421), .A2(new_n425), .A3(new_n423), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n425), .B1(new_n421), .B2(new_n423), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n465), .A2(new_n468), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n468), .B1(new_n465), .B2(new_n478), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT82), .ZN(new_n482));
  OAI21_X1  g296(.A(G214), .B1(G237), .B2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n465), .A2(new_n478), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n467), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n465), .A2(new_n478), .A3(new_n468), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT82), .B1(new_n489), .B2(new_n483), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n419), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n329), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n459), .A2(new_n460), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n370), .A2(new_n378), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n361), .A2(new_n363), .A3(new_n260), .A4(new_n364), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n199), .A2(G137), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n362), .A2(G134), .ZN(new_n498));
  OAI21_X1  g312(.A(G131), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n422), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT64), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT30), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n504));
  AOI211_X1 g318(.A(KEYINPUT64), .B(new_n504), .C1(new_n495), .C2(new_n500), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n494), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n496), .A2(new_n499), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n370), .A2(new_n378), .B1(new_n507), .B2(new_n422), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n493), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n261), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT27), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G101), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n506), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n501), .A2(new_n494), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n504), .B1(new_n508), .B2(KEYINPUT64), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT30), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n520), .B2(new_n494), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT68), .A3(new_n513), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n522), .A3(KEYINPUT31), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n493), .B1(new_n518), .B2(new_n519), .ZN(new_n524));
  INV_X1    g338(.A(new_n513), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n524), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n501), .A2(new_n494), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n509), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT28), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(KEYINPUT28), .B2(new_n517), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n526), .A2(new_n527), .B1(new_n531), .B2(new_n525), .ZN(new_n532));
  AOI211_X1 g346(.A(G472), .B(G902), .C1(new_n523), .C2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT28), .B1(new_n508), .B2(new_n493), .ZN(new_n534));
  AOI211_X1 g348(.A(new_n525), .B(new_n534), .C1(new_n529), .C2(KEYINPUT28), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n535), .B2(KEYINPUT29), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n506), .A2(new_n509), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n525), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n535), .B1(new_n538), .B2(KEYINPUT70), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(KEYINPUT70), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT29), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n536), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n533), .A2(KEYINPUT32), .B1(G472), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n533), .B2(KEYINPUT32), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n523), .B2(new_n532), .ZN(new_n547));
  INV_X1    g361(.A(G472), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT32), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT69), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT23), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n439), .B2(G128), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n554), .B(new_n555), .C1(G119), .C2(new_n191), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G110), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT24), .B(G110), .Z(new_n558));
  XNOR2_X1  g372(.A(G119), .B(G128), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n286), .B2(new_n291), .ZN(new_n562));
  OAI22_X1  g376(.A1(new_n556), .A2(G110), .B1(new_n559), .B2(new_n558), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n291), .A2(new_n297), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT72), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n561), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n280), .A2(new_n271), .A3(new_n285), .ZN(new_n567));
  AOI21_X1  g381(.A(G146), .B1(new_n289), .B2(new_n290), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT72), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n291), .A2(new_n297), .A3(new_n563), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n575), .B(KEYINPUT73), .Z(new_n576));
  NAND3_X1  g390(.A1(new_n565), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n569), .A2(new_n571), .A3(new_n575), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n333), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT74), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT25), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n577), .A2(new_n578), .A3(new_n333), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n188), .B1(G234), .B2(new_n333), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(G902), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n577), .A2(new_n578), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n492), .A2(new_n552), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  AOI21_X1  g407(.A(KEYINPUT68), .B1(new_n521), .B2(new_n513), .ZN(new_n594));
  NOR4_X1   g408(.A1(new_n524), .A2(new_n515), .A3(new_n517), .A4(new_n525), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n594), .A2(new_n595), .A3(new_n527), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n531), .A2(new_n525), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(KEYINPUT31), .B2(new_n514), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n333), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G472), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n549), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n590), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n236), .A2(new_n239), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT33), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n236), .A2(new_n239), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(G478), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n241), .A2(new_n333), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n240), .B2(new_n241), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n328), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n483), .B1(new_n488), .B2(KEYINPUT94), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n481), .B2(KEYINPUT94), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n251), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n602), .A2(new_n419), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT95), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  XOR2_X1   g433(.A(new_n240), .B(new_n242), .Z(new_n620));
  NAND3_X1  g434(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT96), .B1(new_n621), .B2(new_n324), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n621), .A2(KEYINPUT96), .A3(new_n324), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n620), .B(new_n309), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n614), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n602), .A2(new_n625), .A3(new_n419), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NAND2_X1  g442(.A1(new_n565), .A2(new_n572), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n629), .A2(KEYINPUT36), .A3(new_n576), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n576), .A2(KEYINPUT36), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n565), .B2(new_n572), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n588), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n587), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n492), .A2(new_n549), .A3(new_n600), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT97), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n247), .B1(new_n248), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n624), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n635), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n392), .A2(new_n411), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n644), .A2(new_n408), .B1(new_n409), .B2(new_n403), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n645), .A2(G469), .A3(G902), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n392), .A2(new_n411), .A3(new_n414), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n388), .A2(new_n391), .B1(new_n401), .B2(new_n402), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n647), .B(G469), .C1(new_n414), .C2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n334), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n330), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n643), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n552), .A2(new_n642), .A3(new_n613), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  NOR2_X1   g469(.A1(new_n594), .A2(new_n595), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n529), .A2(new_n525), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT99), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n548), .B1(new_n659), .B2(new_n333), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(KEYINPUT32), .B2(new_n533), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n546), .A3(new_n551), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n489), .B(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n664), .A2(new_n484), .A3(new_n243), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n662), .A2(new_n328), .A3(new_n643), .A4(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT100), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT100), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n641), .B(KEYINPUT39), .Z(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n652), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT40), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n667), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  INV_X1    g488(.A(new_n641), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n328), .A2(new_n610), .A3(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n552), .A2(new_n613), .A3(new_n653), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT101), .B(G146), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G48));
  OAI21_X1  g493(.A(G469), .B1(new_n645), .B2(G902), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n330), .A3(new_n418), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n552), .A2(new_n591), .A3(new_n615), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NAND4_X1  g499(.A1(new_n552), .A2(new_n625), .A3(new_n591), .A4(new_n682), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  AOI21_X1  g501(.A(new_n332), .B1(new_n417), .B2(new_n333), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n646), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n613), .A3(new_n635), .A4(new_n330), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n329), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n552), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT102), .B(G119), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G21));
  AOI21_X1  g508(.A(KEYINPUT103), .B1(new_n599), .B2(G472), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n601), .B2(KEYINPUT103), .ZN(new_n696));
  INV_X1    g510(.A(new_n328), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT94), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n484), .B1(new_n479), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n489), .B2(new_n698), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n697), .A2(new_n243), .A3(new_n700), .A4(new_n250), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n696), .A2(new_n701), .A3(new_n591), .A4(new_n682), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n681), .A2(new_n700), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n607), .A2(new_n609), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT87), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n621), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n321), .A3(new_n324), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n706), .B1(new_n709), .B2(new_n309), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n705), .A2(new_n710), .A3(new_n635), .A4(new_n675), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n523), .A2(new_n532), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n548), .B1(new_n712), .B2(new_n333), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT103), .B1(new_n713), .B2(new_n533), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n547), .B2(new_n548), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n704), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n328), .A2(new_n610), .A3(new_n675), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n690), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n696), .A2(new_n720), .A3(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  NAND2_X1  g537(.A1(new_n481), .A2(new_n483), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n725), .B1(new_n419), .B2(new_n726), .ZN(new_n727));
  AOI211_X1 g541(.A(KEYINPUT105), .B(new_n331), .C1(new_n413), .C2(new_n418), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n552), .A3(new_n591), .A4(new_n676), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n727), .A2(new_n719), .A3(new_n728), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n549), .A2(new_n550), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n590), .B1(new_n544), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(KEYINPUT42), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  AND4_X1   g552(.A1(new_n552), .A2(new_n729), .A3(new_n591), .A4(new_n642), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n199), .ZN(G36));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT43), .B1(new_n697), .B2(new_n610), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n328), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n709), .A2(KEYINPUT108), .A3(new_n309), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n607), .A2(KEYINPUT43), .A3(new_n609), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT109), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n744), .A2(new_n745), .A3(new_n749), .A4(new_n746), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n742), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n601), .A2(new_n635), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n741), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n748), .A2(new_n750), .ZN(new_n757));
  INV_X1    g571(.A(new_n742), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(KEYINPUT44), .A3(new_n601), .A4(new_n635), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n334), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n392), .A2(new_n411), .A3(new_n414), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n414), .B1(new_n392), .B2(new_n403), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n647), .B(KEYINPUT45), .C1(new_n414), .C2(new_n648), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(G469), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT106), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n647), .B1(new_n414), .B2(new_n648), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n332), .B1(new_n772), .B2(new_n765), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n769), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n764), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n761), .B1(new_n776), .B2(new_n646), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n774), .B1(new_n773), .B2(new_n769), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n774), .A2(new_n768), .A3(G469), .A4(new_n769), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n763), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(KEYINPUT107), .A3(new_n418), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n778), .A2(new_n779), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n762), .B1(new_n782), .B2(new_n334), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n777), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n330), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n670), .A3(new_n724), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n755), .A2(new_n756), .A3(new_n760), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  XNOR2_X1  g602(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(KEYINPUT111), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n784), .A2(new_n330), .A3(new_n794), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n552), .A2(new_n591), .A3(new_n719), .A4(new_n724), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NAND2_X1  g612(.A1(new_n664), .A2(new_n484), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n717), .A2(new_n799), .A3(new_n590), .A4(new_n681), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n759), .A2(new_n247), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n247), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n681), .A2(new_n724), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n751), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n714), .A2(new_n635), .A3(new_n716), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n751), .A2(new_n804), .ZN(new_n811));
  NOR2_X1   g625(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n800), .A3(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n661), .A2(new_n546), .A3(new_n551), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n591), .A3(new_n247), .A4(new_n805), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n697), .A2(new_n706), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n803), .A2(new_n810), .A3(new_n813), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n807), .B2(new_n809), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n822), .A3(new_n803), .A4(new_n813), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n680), .A2(new_n418), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n330), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n784), .A2(new_n330), .A3(new_n794), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n789), .B1(new_n784), .B2(new_n330), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n717), .A2(new_n590), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n247), .A2(new_n759), .A3(new_n831), .A4(new_n725), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n824), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n820), .A2(new_n823), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n811), .A2(new_n705), .A3(new_n831), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n835), .B(new_n245), .C1(new_n611), .C2(new_n815), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n807), .A2(new_n735), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(KEYINPUT48), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(KEYINPUT48), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n826), .B1(new_n791), .B2(new_n795), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n811), .A2(new_n831), .A3(new_n725), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n841), .A2(KEYINPUT115), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n830), .B2(new_n832), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n843), .A2(new_n845), .A3(new_n819), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n834), .B(new_n840), .C1(new_n846), .C2(KEYINPUT51), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT118), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n243), .A2(new_n309), .A3(new_n675), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n623), .A2(new_n622), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n850), .A2(new_n851), .A3(new_n724), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n552), .A2(new_n653), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n809), .B2(new_n733), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n724), .B1(new_n652), .B2(KEYINPUT105), .ZN(new_n856));
  INV_X1    g670(.A(new_n728), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n676), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n858), .A2(new_n808), .A3(KEYINPUT112), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n853), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n702), .A2(new_n686), .A3(new_n683), .A4(new_n692), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n491), .A2(new_n250), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n611), .B1(new_n328), .B2(new_n243), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n602), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n636), .A2(new_n592), .A3(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n860), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n552), .A2(new_n613), .A3(new_n653), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n642), .A2(new_n867), .B1(new_n718), .B2(new_n721), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n700), .A2(new_n243), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n328), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n652), .A2(new_n641), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n662), .A2(new_n872), .A3(new_n643), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n868), .A2(new_n869), .A3(new_n677), .A4(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n722), .A2(new_n654), .A3(new_n677), .A4(new_n874), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT52), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n739), .B1(new_n732), .B2(new_n736), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n866), .A2(new_n875), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n876), .A2(new_n868), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n849), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n861), .ZN(new_n882));
  INV_X1    g696(.A(new_n865), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n809), .A2(new_n733), .A3(new_n854), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT112), .B1(new_n858), .B2(new_n808), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n552), .A2(new_n653), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n884), .A2(new_n885), .B1(new_n886), .B2(new_n852), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n878), .A2(new_n882), .A3(new_n883), .A4(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n876), .A2(KEYINPUT52), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n875), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n881), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT54), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT115), .B1(new_n841), .B2(new_n842), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n803), .A2(new_n813), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n821), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n824), .B1(new_n898), .B2(new_n843), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n834), .A4(new_n840), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n879), .A2(new_n891), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT114), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n905));
  INV_X1    g719(.A(new_n880), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n890), .A2(KEYINPUT53), .A3(new_n875), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n879), .A2(KEYINPUT114), .A3(new_n891), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n904), .A2(new_n905), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n848), .A2(new_n895), .A3(new_n901), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT119), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n895), .A2(new_n909), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n848), .A4(new_n901), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n244), .A2(new_n257), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n689), .B(KEYINPUT49), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n706), .A2(new_n331), .A3(new_n484), .ZN(new_n918));
  AND4_X1   g732(.A1(new_n591), .A2(new_n917), .A3(new_n664), .A4(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n919), .A2(new_n814), .A3(new_n744), .A4(new_n745), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n920), .ZN(G75));
  NAND3_X1  g735(.A1(new_n904), .A2(new_n907), .A3(new_n908), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(G902), .A3(new_n467), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n472), .A2(new_n474), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n477), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n923), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n928), .B1(new_n923), .B2(new_n924), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n257), .A2(G952), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(G51));
  NAND2_X1  g746(.A1(new_n907), .A2(new_n908), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT114), .B1(new_n879), .B2(new_n891), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT54), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(KEYINPUT121), .A3(new_n909), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n922), .A2(new_n937), .A3(KEYINPUT54), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n334), .B(KEYINPUT57), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n417), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n922), .A2(G902), .A3(new_n782), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n931), .B1(new_n941), .B2(new_n942), .ZN(G54));
  NAND2_X1  g757(.A1(new_n922), .A2(G902), .ZN(new_n944));
  NAND2_X1  g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n322), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n931), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n944), .A2(new_n322), .A3(new_n945), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(G60));
  NAND2_X1  g764(.A1(new_n604), .A2(new_n606), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT122), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n608), .B(KEYINPUT59), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n938), .A2(new_n936), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n895), .B2(new_n909), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n947), .B1(new_n956), .B2(new_n952), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(G63));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n922), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n577), .A2(new_n578), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n633), .B(KEYINPUT123), .Z(new_n965));
  NAND3_X1  g779(.A1(new_n922), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n947), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n964), .A2(KEYINPUT61), .A3(new_n947), .A4(new_n966), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(G66));
  INV_X1    g785(.A(G224), .ZN(new_n972));
  OAI21_X1  g786(.A(G953), .B1(new_n249), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n861), .A2(new_n865), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n925), .B1(G898), .B2(new_n257), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  XNOR2_X1  g791(.A(new_n520), .B(new_n314), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n868), .A2(new_n677), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n673), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(KEYINPUT62), .A3(new_n673), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n552), .A2(new_n591), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n863), .A2(new_n671), .A3(new_n725), .ZN(new_n987));
  AOI22_X1  g801(.A1(new_n983), .A2(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n988), .A2(new_n787), .A3(new_n797), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n978), .B1(new_n989), .B2(G953), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n640), .A2(G953), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT124), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n787), .A2(new_n797), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n878), .A2(KEYINPUT125), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n878), .A2(KEYINPUT125), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n735), .A2(new_n872), .ZN(new_n996));
  OR3_X1    g810(.A1(new_n785), .A2(new_n670), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n994), .A2(new_n980), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n992), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  INV_X1    g814(.A(new_n978), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n990), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G72));
  XOR2_X1   g819(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1006));
  NOR2_X1   g820(.A1(new_n548), .A2(new_n333), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n656), .A2(new_n538), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n894), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1008), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(new_n989), .B2(new_n974), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n537), .A2(new_n513), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n999), .A2(new_n974), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1015), .A2(new_n1008), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n521), .A2(new_n525), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n947), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g834(.A(KEYINPUT127), .B(new_n947), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1014), .B1(new_n1020), .B2(new_n1021), .ZN(G57));
endmodule


