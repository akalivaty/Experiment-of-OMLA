//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G116), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n194), .B(new_n196), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n196), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT2), .B(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n203), .A3(KEYINPUT67), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G101), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n206), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(G101), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT76), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n208), .A2(new_n211), .A3(new_n219), .A4(new_n212), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT4), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n213), .A2(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(KEYINPUT4), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT76), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n216), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT5), .ZN(new_n226));
  OAI21_X1  g040(.A(G113), .B1(new_n194), .B2(KEYINPUT5), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n200), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n207), .A2(G107), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n210), .A2(G104), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n220), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n190), .B(new_n192), .C1(new_n225), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n224), .A2(new_n221), .ZN(new_n235));
  INV_X1    g049(.A(new_n216), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n191), .B1(new_n237), .B2(new_n189), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n189), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n234), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n241), .A2(KEYINPUT64), .A3(G143), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G146), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n244), .A2(new_n246), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n242), .A2(new_n249), .ZN(new_n251));
  OR2_X1    g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n245), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G125), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n248), .A2(G146), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n258));
  OAI21_X1  g072(.A(G128), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n251), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n244), .A2(new_n247), .A3(new_n249), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G125), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G224), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n266), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n240), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT81), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n240), .A2(new_n274), .A3(new_n271), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n264), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n255), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n278), .A2(KEYINPUT83), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n256), .B1(new_n278), .B2(KEYINPUT83), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n279), .A2(new_n280), .B1(KEYINPUT7), .B2(new_n268), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n189), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n233), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n228), .A2(new_n232), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n268), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n281), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n190), .B(new_n233), .C1(new_n235), .C2(new_n236), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n188), .B1(new_n276), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n190), .B1(new_n225), .B2(new_n233), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n293), .B1(new_n289), .B2(new_n191), .ZN(new_n294));
  AOI211_X1 g108(.A(KEYINPUT81), .B(new_n270), .C1(new_n294), .C2(new_n234), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n274), .B1(new_n240), .B2(new_n271), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n188), .B(new_n291), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n187), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G478), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(KEYINPUT15), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(KEYINPUT15), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G128), .B(G143), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G122), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT86), .B1(new_n310), .B2(G116), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT86), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n195), .A3(G122), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n310), .A2(G116), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G107), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n210), .A3(new_n315), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT13), .B1(new_n248), .B2(G128), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT87), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n248), .A2(KEYINPUT13), .A3(G128), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n321), .B(new_n322), .C1(G128), .C2(new_n248), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G134), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(KEYINPUT88), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(new_n323), .B2(G134), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n309), .B(new_n319), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n314), .A2(KEYINPUT14), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n314), .A2(KEYINPUT14), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n315), .A3(new_n330), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n307), .A2(new_n308), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n331), .A2(G107), .B1(new_n309), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n318), .B(KEYINPUT89), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT90), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n335), .B1(new_n333), .B2(new_n334), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n328), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT9), .B(G234), .Z(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT75), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(G217), .A3(new_n267), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n342), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n328), .B(new_n344), .C1(new_n337), .C2(new_n338), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT69), .B(G902), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n306), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n347), .ZN(new_n349));
  AOI211_X1 g163(.A(new_n349), .B(new_n305), .C1(new_n343), .C2(new_n345), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G131), .ZN(new_n352));
  NOR2_X1   g166(.A1(G237), .A2(G953), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(new_n248), .ZN(new_n355));
  NOR2_X1   g169(.A1(KEYINPUT84), .A2(G143), .ZN(new_n356));
  OAI211_X1 g170(.A(G214), .B(new_n353), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(G214), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n354), .B2(new_n248), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n352), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT17), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n357), .A2(new_n359), .A3(new_n352), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n363), .B1(new_n366), .B2(new_n362), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n255), .A2(KEYINPUT16), .A3(G140), .ZN(new_n368));
  XNOR2_X1  g182(.A(G125), .B(G140), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(KEYINPUT16), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n241), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT72), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(G146), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(KEYINPUT72), .A3(new_n241), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n360), .A2(KEYINPUT18), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n369), .B(new_n241), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT18), .A2(G131), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n357), .A2(new_n359), .A3(new_n380), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n367), .A2(new_n377), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n207), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n374), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n369), .B(KEYINPUT19), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n387), .B1(new_n241), .B2(new_n388), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n389), .A2(new_n365), .B1(new_n378), .B2(new_n382), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n385), .B1(new_n390), .B2(KEYINPUT85), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(KEYINPUT85), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n386), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NOR2_X1   g209(.A1(G475), .A2(G902), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n393), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n398), .A2(new_n391), .B1(new_n383), .B2(new_n385), .ZN(new_n399));
  INV_X1    g213(.A(new_n396), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT20), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G902), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n383), .A2(new_n385), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n383), .A2(new_n385), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n397), .A2(new_n401), .B1(G475), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(G234), .A2(G237), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(G952), .A3(new_n267), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT92), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n349), .A2(G953), .A3(new_n407), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT21), .B(G898), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n351), .A2(new_n406), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT93), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n351), .A2(new_n406), .A3(KEYINPUT93), .A4(new_n414), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n299), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n204), .A2(new_n206), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT11), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n308), .B2(G137), .ZN(new_n423));
  INV_X1    g237(.A(G137), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT11), .A3(G134), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n308), .A2(G137), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G131), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT66), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n423), .A2(new_n425), .A3(new_n352), .A4(new_n426), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n427), .A2(KEYINPUT66), .A3(G131), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n254), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n426), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n308), .A2(G137), .ZN(new_n435));
  OAI21_X1  g249(.A(G131), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n264), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n250), .A2(new_n253), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT65), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT65), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n250), .A2(new_n253), .A3(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n440), .A2(new_n431), .A3(new_n432), .A4(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n443), .A2(new_n437), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n421), .B(new_n438), .C1(new_n444), .C2(KEYINPUT30), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n433), .A2(new_n437), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n420), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n353), .A2(G210), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n450), .B(KEYINPUT27), .Z(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT26), .B(G101), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT28), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n443), .A2(new_n437), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n421), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n448), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n447), .A2(KEYINPUT68), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n421), .B1(new_n446), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT28), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n459), .A2(new_n463), .A3(new_n453), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n455), .A2(new_n464), .A3(KEYINPUT29), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n446), .B(new_n421), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n460), .A2(new_n462), .ZN(new_n467));
  MUX2_X1   g281(.A(new_n466), .B(new_n467), .S(new_n456), .Z(new_n468));
  INV_X1    g282(.A(new_n453), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT29), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n347), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G472), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT31), .B1(new_n449), .B2(new_n453), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n453), .B1(new_n459), .B2(new_n463), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT31), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n445), .A2(new_n475), .A3(new_n448), .A4(new_n469), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT32), .ZN(new_n478));
  NOR2_X1   g292(.A1(G472), .A2(G902), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n472), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G217), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n347), .B2(G234), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n261), .A2(KEYINPUT23), .A3(G119), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n261), .A2(G119), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT71), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n261), .A2(KEYINPUT71), .A3(G119), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n193), .A2(G128), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT23), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT23), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n486), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n487), .A2(new_n492), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT24), .B(G110), .Z(new_n500));
  AOI22_X1  g314(.A1(new_n498), .A2(G110), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n375), .A2(new_n501), .A3(new_n376), .ZN(new_n502));
  INV_X1    g316(.A(G110), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n486), .C1(new_n491), .C2(new_n497), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n499), .A2(new_n500), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n369), .A2(new_n241), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n370), .B2(G146), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n506), .A2(KEYINPUT73), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT73), .B1(new_n506), .B2(new_n508), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT74), .B(new_n502), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT22), .B(G137), .ZN(new_n515));
  INV_X1    g329(.A(G221), .ZN(new_n516));
  INV_X1    g330(.A(G234), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n516), .A2(new_n517), .A3(G953), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n515), .B(new_n518), .Z(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n511), .A2(new_n512), .A3(new_n519), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT25), .B1(new_n523), .B2(new_n347), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n525), .B(new_n349), .C1(new_n521), .C2(new_n522), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n485), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n485), .A2(G902), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n483), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n516), .B1(new_n341), .B2(new_n402), .ZN(new_n534));
  XNOR2_X1  g348(.A(G110), .B(G140), .ZN(new_n535));
  INV_X1    g349(.A(G227), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(G953), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n535), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n254), .A2(new_n215), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n221), .B2(new_n224), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n220), .A2(new_n231), .A3(KEYINPUT10), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n264), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n244), .A2(new_n247), .A3(new_n249), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n259), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n232), .B1(new_n544), .B2(new_n263), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT77), .B(KEYINPUT10), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n431), .A2(new_n432), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n538), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n545), .B1(new_n277), .B2(new_n232), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n552), .B2(new_n549), .ZN(new_n553));
  INV_X1    g367(.A(new_n549), .ZN(new_n554));
  INV_X1    g368(.A(new_n232), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n264), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n554), .B(KEYINPUT12), .C1(new_n545), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n538), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n235), .A2(new_n254), .A3(new_n215), .ZN(new_n561));
  INV_X1    g375(.A(new_n547), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n549), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n554), .B1(new_n540), .B2(new_n547), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n559), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n566), .A2(new_n347), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT79), .B(G469), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n560), .B1(new_n558), .B2(new_n563), .ZN(new_n570));
  INV_X1    g384(.A(new_n564), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n550), .B2(KEYINPUT78), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n563), .A2(new_n560), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n570), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G469), .B1(new_n576), .B2(G902), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n534), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n419), .A2(new_n533), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(G101), .ZN(G3));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n299), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n187), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n291), .B1(new_n295), .B2(new_n296), .ZN(new_n584));
  INV_X1    g398(.A(new_n188), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n583), .B1(new_n586), .B2(new_n297), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT94), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n413), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n477), .A2(new_n347), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n592), .A2(G472), .B1(new_n479), .B2(new_n477), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n531), .A2(new_n578), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n339), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT33), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n346), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n343), .A2(new_n596), .A3(new_n345), .A4(KEYINPUT33), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n349), .A2(new_n300), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n346), .A2(new_n347), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n300), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n405), .A2(G475), .ZN(new_n605));
  INV_X1    g419(.A(new_n397), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n395), .B1(new_n394), .B2(new_n396), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n591), .A2(new_n594), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NAND3_X1  g427(.A1(new_n397), .A2(new_n401), .A3(KEYINPUT96), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n616), .A3(new_n605), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n351), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n591), .A2(new_n594), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  INV_X1    g435(.A(new_n485), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n514), .A2(new_n520), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n506), .A2(new_n508), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT73), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n506), .A2(KEYINPUT73), .A3(new_n508), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT74), .B1(new_n628), .B2(new_n502), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n522), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n347), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n525), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n523), .A2(KEYINPUT25), .A3(new_n347), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n622), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n511), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n528), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT97), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n527), .A2(new_n641), .A3(new_n638), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n419), .A2(new_n643), .A3(new_n578), .A4(new_n593), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  XOR2_X1   g460(.A(KEYINPUT98), .B(G900), .Z(new_n647));
  AOI21_X1  g461(.A(new_n410), .B1(new_n411), .B2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n617), .A2(new_n351), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n586), .A2(new_n297), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT94), .B1(new_n650), .B2(new_n187), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n581), .B(new_n583), .C1(new_n586), .C2(new_n297), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n483), .A2(new_n640), .A3(new_n578), .A4(new_n642), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT99), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AND4_X1   g469(.A1(new_n483), .A2(new_n640), .A3(new_n578), .A4(new_n642), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n656), .A2(new_n589), .A3(new_n657), .A4(new_n649), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XOR2_X1   g474(.A(new_n648), .B(KEYINPUT39), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n578), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT40), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n650), .B(KEYINPUT38), .ZN(new_n664));
  INV_X1    g478(.A(G472), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n466), .A2(new_n469), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(G902), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n449), .A2(new_n469), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n477), .A2(new_n479), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT32), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n669), .B1(new_n671), .B2(new_n480), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n608), .B1(new_n348), .B2(new_n350), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n527), .A2(new_n638), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n672), .A2(new_n673), .A3(new_n583), .A4(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n663), .A2(new_n664), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT100), .B(G143), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G45));
  INV_X1    g492(.A(new_n648), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n604), .A2(new_n608), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n582), .B2(new_n588), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n656), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  INV_X1    g497(.A(new_n534), .ZN(new_n684));
  INV_X1    g498(.A(G469), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n569), .B(new_n684), .C1(new_n685), .C2(new_n567), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n532), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n589), .A3(new_n414), .A4(new_n610), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n687), .A2(new_n589), .A3(new_n414), .A4(new_n618), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NAND2_X1  g506(.A1(new_n417), .A2(new_n418), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n643), .A3(new_n483), .ZN(new_n694));
  INV_X1    g508(.A(new_n686), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(new_n651), .B2(new_n652), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT101), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n589), .A2(KEYINPUT101), .A3(new_n695), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n694), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT102), .B(G119), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G21));
  NAND2_X1  g516(.A1(new_n468), .A2(new_n453), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n473), .A3(new_n476), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n479), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT103), .B1(new_n592), .B2(G472), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n707), .B(new_n665), .C1(new_n477), .C2(new_n347), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n530), .ZN(new_n710));
  INV_X1    g524(.A(new_n673), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n686), .A2(new_n413), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n710), .A2(new_n589), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  INV_X1    g528(.A(new_n674), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n709), .A2(new_n680), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT101), .B1(new_n589), .B2(new_n695), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n697), .B(new_n686), .C1(new_n582), .C2(new_n588), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NOR2_X1   g534(.A1(new_n650), .A2(new_n583), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n570), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n724), .A2(new_n685), .A3(G902), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n564), .B1(new_n573), .B2(new_n574), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n550), .A2(KEYINPUT78), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n723), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n577), .B2(new_n724), .ZN(new_n730));
  INV_X1    g544(.A(new_n569), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n684), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n722), .A2(new_n532), .A3(new_n732), .A4(new_n680), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT42), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G131), .ZN(G33));
  NOR2_X1   g549(.A1(new_n722), .A2(new_n732), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n533), .A3(new_n649), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT105), .B(G134), .Z(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G36));
  OAI21_X1  g553(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n685), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n741), .B2(new_n740), .ZN(new_n743));
  NAND2_X1  g557(.A1(G469), .A2(G902), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n569), .B1(new_n745), .B2(KEYINPUT46), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n684), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n661), .ZN(new_n751));
  INV_X1    g565(.A(new_n604), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n752), .A2(KEYINPUT43), .A3(new_n608), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n406), .B(KEYINPUT106), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n604), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n753), .B1(new_n755), .B2(KEYINPUT43), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n715), .A2(new_n593), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT44), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n756), .A2(KEYINPUT44), .A3(new_n757), .ZN(new_n759));
  OR4_X1    g573(.A1(new_n722), .A2(new_n751), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  OAI21_X1  g575(.A(new_n749), .B1(KEYINPUT107), .B2(KEYINPUT47), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n722), .A2(new_n531), .A3(new_n680), .A4(new_n483), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n764));
  OAI211_X1 g578(.A(new_n762), .B(new_n763), .C1(new_n749), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n698), .A2(new_n699), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n769), .A2(new_n716), .B1(new_n655), .B2(new_n658), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n672), .B(new_n673), .C1(new_n582), .C2(new_n588), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n527), .A2(new_n638), .A3(new_n679), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT112), .B1(new_n732), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n685), .B1(new_n740), .B2(new_n402), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n728), .B1(new_n774), .B2(KEYINPUT104), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n534), .B1(new_n775), .B2(new_n569), .ZN(new_n776));
  INV_X1    g590(.A(new_n772), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n771), .A2(new_n780), .B1(new_n656), .B2(new_n681), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n768), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n768), .A2(new_n719), .A3(new_n781), .A4(new_n659), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT113), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n719), .A2(new_n781), .A3(new_n659), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT52), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n770), .A2(new_n768), .A3(new_n781), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n609), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n299), .A2(new_n413), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n594), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n608), .A2(new_n351), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(KEYINPUT110), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n414), .A3(new_n587), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n798), .A3(new_n594), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n793), .A2(new_n799), .A3(new_n644), .A4(new_n579), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n351), .A2(new_n679), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n617), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n802), .A2(new_n617), .A3(new_n801), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n656), .A2(new_n721), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n716), .A2(new_n736), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n737), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n800), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n688), .A2(new_n691), .A3(new_n713), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n700), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n808), .A2(new_n810), .A3(new_n734), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n784), .A2(new_n789), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT53), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n786), .A2(new_n787), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n808), .A2(new_n810), .A3(new_n734), .A4(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT54), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n812), .A2(new_n816), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n810), .A2(new_n734), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(new_n824));
  AND4_X1   g638(.A1(KEYINPUT53), .A2(new_n786), .A3(new_n787), .A4(new_n808), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n820), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n818), .B1(new_n812), .B2(KEYINPUT53), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n814), .B1(new_n830), .B2(KEYINPUT54), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n767), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n762), .B1(new_n749), .B2(new_n764), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n569), .B1(new_n685), .B2(new_n567), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n684), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n756), .A2(new_n410), .A3(new_n710), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n721), .A3(new_n837), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n836), .A2(new_n187), .A3(new_n664), .A4(new_n686), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT50), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n756), .A2(new_n410), .A3(new_n695), .A4(new_n721), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT117), .Z(new_n842));
  NOR2_X1   g656(.A1(new_n709), .A2(new_n715), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n672), .A2(new_n531), .A3(new_n410), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n844), .A2(new_n722), .A3(new_n686), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n604), .A2(new_n608), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n842), .A2(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n838), .A2(new_n840), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n842), .A2(new_n533), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n851), .A2(KEYINPUT119), .A3(KEYINPUT48), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n845), .A2(new_n610), .ZN(new_n853));
  XNOR2_X1  g667(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n836), .B1(new_n698), .B2(new_n699), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n848), .A2(new_n849), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n850), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n813), .A2(KEYINPUT54), .A3(new_n819), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT116), .A3(new_n828), .A4(new_n820), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n832), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(G952), .B(new_n267), .C1(new_n863), .C2(KEYINPUT118), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n865));
  OAI21_X1  g679(.A(G953), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n530), .A2(new_n583), .A3(new_n534), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT108), .ZN(new_n868));
  INV_X1    g682(.A(new_n664), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n834), .B(KEYINPUT49), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n755), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n868), .A2(new_n869), .A3(new_n871), .A4(new_n672), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n864), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT120), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(G75));
  NOR2_X1   g691(.A1(new_n267), .A2(G952), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n347), .B1(new_n821), .B2(new_n826), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n880), .B2(new_n585), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n240), .B(new_n270), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT55), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n879), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n881), .B2(new_n883), .ZN(G51));
  NAND2_X1  g699(.A1(new_n821), .A2(new_n826), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n828), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n744), .B(KEYINPUT57), .Z(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n566), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n880), .B(new_n742), .C1(new_n741), .C2(new_n740), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n878), .B1(new_n891), .B2(new_n892), .ZN(G54));
  NAND3_X1  g707(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n894), .A2(KEYINPUT121), .A3(new_n399), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n879), .B1(new_n894), .B2(new_n399), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT121), .B1(new_n894), .B2(new_n399), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G60));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT59), .Z(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n832), .B2(new_n862), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n598), .A2(new_n599), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT122), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n900), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n878), .B1(new_n888), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n901), .A2(KEYINPUT122), .A3(new_n902), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT123), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n901), .A2(KEYINPUT122), .A3(new_n902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n903), .A4(new_n906), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n909), .A2(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT60), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n886), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT124), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n878), .B1(new_n917), .B2(new_n637), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n523), .B(KEYINPUT125), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G66));
  INV_X1    g736(.A(new_n412), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n267), .B1(new_n923), .B2(G224), .ZN(new_n924));
  OR3_X1    g738(.A1(new_n800), .A2(new_n809), .A3(new_n700), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n267), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n294), .B(new_n234), .C1(G898), .C2(new_n267), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n926), .B(new_n927), .Z(G69));
  MUX2_X1   g742(.A(new_n444), .B(new_n446), .S(KEYINPUT30), .Z(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n388), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(G900), .B(G953), .C1(new_n931), .C2(new_n536), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n536), .B2(new_n931), .ZN(new_n933));
  INV_X1    g747(.A(new_n737), .ZN(new_n934));
  INV_X1    g748(.A(new_n751), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n590), .A2(new_n532), .A3(new_n673), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n760), .A2(new_n937), .A3(new_n734), .A4(new_n765), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n770), .A2(new_n682), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(G953), .B1(new_n940), .B2(new_n930), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n770), .A2(new_n676), .A3(new_n682), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n722), .A2(new_n662), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n944), .B(new_n533), .C1(new_n791), .C2(new_n794), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n760), .A2(new_n765), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n931), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n933), .B1(new_n941), .B2(new_n950), .ZN(G72));
  XNOR2_X1  g765(.A(new_n449), .B(new_n469), .ZN(new_n952));
  NAND2_X1  g766(.A1(G472), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT63), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n878), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n946), .A2(new_n949), .A3(new_n668), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n449), .A2(new_n469), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n940), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n956), .B1(new_n959), .B2(new_n925), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n952), .A2(new_n955), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n830), .B2(new_n961), .ZN(G57));
endmodule


