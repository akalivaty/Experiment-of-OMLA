

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589;

  XOR2_X1 U320 ( .A(n455), .B(n454), .Z(n541) );
  XNOR2_X1 U321 ( .A(n333), .B(n332), .ZN(n334) );
  NOR2_X1 U322 ( .A1(n579), .A2(n342), .ZN(n343) );
  INV_X1 U323 ( .A(KEYINPUT70), .ZN(n288) );
  XNOR2_X1 U324 ( .A(n289), .B(n288), .ZN(n291) );
  XNOR2_X1 U325 ( .A(n291), .B(n290), .ZN(n424) );
  XOR2_X1 U326 ( .A(n325), .B(KEYINPUT10), .Z(n327) );
  XNOR2_X1 U327 ( .A(n297), .B(n296), .ZN(n325) );
  NOR2_X1 U328 ( .A1(n573), .A2(n477), .ZN(n431) );
  NAND2_X1 U329 ( .A1(n418), .A2(n528), .ZN(n573) );
  XNOR2_X1 U330 ( .A(n298), .B(n325), .ZN(n299) );
  XNOR2_X1 U331 ( .A(n300), .B(n299), .ZN(n305) );
  XNOR2_X1 U332 ( .A(n335), .B(n334), .ZN(n339) );
  XNOR2_X1 U333 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U334 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XNOR2_X1 U335 ( .A(G204GAT), .B(G78GAT), .ZN(n289) );
  XOR2_X1 U336 ( .A(G148GAT), .B(G106GAT), .Z(n290) );
  XNOR2_X1 U337 ( .A(n424), .B(KEYINPUT73), .ZN(n293) );
  XOR2_X1 U338 ( .A(G71GAT), .B(KEYINPUT13), .Z(n308) );
  XOR2_X1 U339 ( .A(n308), .B(KEYINPUT32), .Z(n292) );
  OR2_X1 U340 ( .A1(n293), .A2(n292), .ZN(n295) );
  NAND2_X1 U341 ( .A1(n293), .A2(n292), .ZN(n294) );
  NAND2_X1 U342 ( .A1(n295), .A2(n294), .ZN(n300) );
  XOR2_X1 U343 ( .A(G120GAT), .B(G57GAT), .Z(n404) );
  XOR2_X1 U344 ( .A(G176GAT), .B(G64GAT), .Z(n378) );
  XOR2_X1 U345 ( .A(n404), .B(n378), .Z(n298) );
  XOR2_X1 U346 ( .A(KEYINPUT71), .B(G92GAT), .Z(n297) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .ZN(n296) );
  XOR2_X1 U348 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n302) );
  NAND2_X1 U349 ( .A1(G230GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(KEYINPUT31), .B(n303), .Z(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n579) );
  XOR2_X1 U353 ( .A(n579), .B(KEYINPUT41), .Z(n558) );
  INV_X1 U354 ( .A(n558), .ZN(n515) );
  XOR2_X1 U355 ( .A(G57GAT), .B(G211GAT), .Z(n307) );
  XNOR2_X1 U356 ( .A(G183GAT), .B(G127GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n322) );
  XOR2_X1 U358 ( .A(n308), .B(G155GAT), .Z(n311) );
  XNOR2_X1 U359 ( .A(G22GAT), .B(G15GAT), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n309), .B(G8GAT), .ZN(n350) );
  XNOR2_X1 U361 ( .A(n350), .B(G78GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U363 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n313) );
  NAND2_X1 U364 ( .A1(G231GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U367 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n317) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(G64GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n318), .B(KEYINPUT15), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n583) );
  INV_X1 U373 ( .A(n583), .ZN(n569) );
  INV_X1 U374 ( .A(KEYINPUT36), .ZN(n340) );
  XOR2_X1 U375 ( .A(G36GAT), .B(G190GAT), .Z(n381) );
  XOR2_X1 U376 ( .A(KEYINPUT76), .B(n381), .Z(n324) );
  XOR2_X1 U377 ( .A(G29GAT), .B(G134GAT), .Z(n405) );
  XNOR2_X1 U378 ( .A(G218GAT), .B(n405), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n329) );
  NAND2_X1 U380 ( .A1(G232GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U382 ( .A(n329), .B(n328), .Z(n335) );
  XOR2_X1 U383 ( .A(KEYINPUT75), .B(KEYINPUT9), .Z(n331) );
  XNOR2_X1 U384 ( .A(KEYINPUT65), .B(KEYINPUT11), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n333) );
  XNOR2_X1 U386 ( .A(G106GAT), .B(G162GAT), .ZN(n332) );
  XOR2_X1 U387 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n337) );
  XNOR2_X1 U388 ( .A(G50GAT), .B(G43GAT), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U390 ( .A(KEYINPUT69), .B(n338), .ZN(n357) );
  XNOR2_X1 U391 ( .A(n339), .B(n357), .ZN(n565) );
  XNOR2_X1 U392 ( .A(n340), .B(n565), .ZN(n498) );
  NOR2_X1 U393 ( .A1(n569), .A2(n498), .ZN(n341) );
  XOR2_X1 U394 ( .A(KEYINPUT45), .B(n341), .Z(n342) );
  NAND2_X1 U395 ( .A1(KEYINPUT114), .A2(n343), .ZN(n347) );
  INV_X1 U396 ( .A(KEYINPUT114), .ZN(n345) );
  INV_X1 U397 ( .A(n343), .ZN(n344) );
  NAND2_X1 U398 ( .A1(n345), .A2(n344), .ZN(n346) );
  NAND2_X1 U399 ( .A1(n347), .A2(n346), .ZN(n362) );
  XOR2_X1 U400 ( .A(KEYINPUT67), .B(G197GAT), .Z(n349) );
  XNOR2_X1 U401 ( .A(G169GAT), .B(G141GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n361) );
  XOR2_X1 U403 ( .A(G113GAT), .B(G1GAT), .Z(n401) );
  XOR2_X1 U404 ( .A(n350), .B(n401), .Z(n352) );
  XNOR2_X1 U405 ( .A(G36GAT), .B(G29GAT), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U407 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n354) );
  NAND2_X1 U408 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U410 ( .A(n356), .B(n355), .Z(n359) );
  XOR2_X1 U411 ( .A(n357), .B(KEYINPUT29), .Z(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n361), .B(n360), .ZN(n576) );
  INV_X1 U414 ( .A(n576), .ZN(n567) );
  NAND2_X1 U415 ( .A1(n362), .A2(n567), .ZN(n371) );
  NAND2_X1 U416 ( .A1(n558), .A2(n576), .ZN(n364) );
  XNOR2_X1 U417 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n365) );
  NAND2_X1 U419 ( .A1(n365), .A2(n569), .ZN(n367) );
  INV_X1 U420 ( .A(KEYINPUT113), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n368) );
  NOR2_X1 U422 ( .A1(n368), .A2(n565), .ZN(n369) );
  XNOR2_X1 U423 ( .A(KEYINPUT47), .B(n369), .ZN(n370) );
  NAND2_X1 U424 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n372), .B(KEYINPUT48), .ZN(n539) );
  XOR2_X1 U426 ( .A(KEYINPUT18), .B(KEYINPUT81), .Z(n374) );
  XNOR2_X1 U427 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U429 ( .A(n375), .B(KEYINPUT82), .Z(n377) );
  XNOR2_X1 U430 ( .A(G169GAT), .B(G183GAT), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n377), .B(n376), .ZN(n455) );
  XOR2_X1 U432 ( .A(KEYINPUT95), .B(n378), .Z(n380) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U435 ( .A(n382), .B(n381), .Z(n391) );
  XNOR2_X1 U436 ( .A(G211GAT), .B(KEYINPUT88), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n383), .B(KEYINPUT87), .ZN(n384) );
  XOR2_X1 U438 ( .A(n384), .B(KEYINPUT21), .Z(n386) );
  XNOR2_X1 U439 ( .A(G197GAT), .B(G218GAT), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n386), .B(n385), .ZN(n425) );
  XOR2_X1 U441 ( .A(KEYINPUT96), .B(G92GAT), .Z(n388) );
  XNOR2_X1 U442 ( .A(G8GAT), .B(G204GAT), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n425), .B(n389), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n455), .B(n392), .ZN(n530) );
  INV_X1 U447 ( .A(n530), .ZN(n393) );
  NAND2_X1 U448 ( .A1(n539), .A2(n393), .ZN(n395) );
  XOR2_X1 U449 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n418) );
  XOR2_X1 U451 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n397) );
  XNOR2_X1 U452 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n417) );
  XOR2_X1 U454 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n399) );
  XNOR2_X1 U455 ( .A(KEYINPUT5), .B(KEYINPUT93), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U457 ( .A(n400), .B(G85GAT), .Z(n403) );
  XNOR2_X1 U458 ( .A(n401), .B(G148GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n409) );
  XOR2_X1 U460 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U461 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U463 ( .A(n409), .B(n408), .Z(n415) );
  XOR2_X1 U464 ( .A(KEYINPUT0), .B(G127GAT), .Z(n445) );
  XNOR2_X1 U465 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n410), .B(KEYINPUT89), .ZN(n411) );
  XOR2_X1 U467 ( .A(n411), .B(KEYINPUT3), .Z(n413) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(G162GAT), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n423) );
  XNOR2_X1 U470 ( .A(n445), .B(n423), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n483) );
  XNOR2_X1 U473 ( .A(KEYINPUT94), .B(n483), .ZN(n528) );
  XOR2_X1 U474 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n420) );
  XNOR2_X1 U475 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U477 ( .A(G50GAT), .B(G22GAT), .Z(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n428) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n430) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n477) );
  XNOR2_X1 U484 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n432) );
  NAND2_X1 U485 ( .A1(n431), .A2(n432), .ZN(n436) );
  INV_X1 U486 ( .A(n431), .ZN(n434) );
  INV_X1 U487 ( .A(n432), .ZN(n433) );
  NAND2_X1 U488 ( .A1(n434), .A2(n433), .ZN(n435) );
  NAND2_X1 U489 ( .A1(n436), .A2(n435), .ZN(n456) );
  XOR2_X1 U490 ( .A(KEYINPUT80), .B(KEYINPUT84), .Z(n438) );
  XNOR2_X1 U491 ( .A(KEYINPUT85), .B(G176GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U493 ( .A(G120GAT), .B(KEYINPUT20), .Z(n440) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G134GAT), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n453) );
  XOR2_X1 U497 ( .A(G71GAT), .B(KEYINPUT64), .Z(n444) );
  XNOR2_X1 U498 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n449) );
  XOR2_X1 U500 ( .A(G190GAT), .B(G99GAT), .Z(n447) );
  XNOR2_X1 U501 ( .A(G15GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n451) );
  NAND2_X1 U504 ( .A1(G227GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n454) );
  INV_X1 U507 ( .A(n541), .ZN(n470) );
  NAND2_X1 U508 ( .A1(n456), .A2(n470), .ZN(n460) );
  NOR2_X1 U509 ( .A1(n515), .A2(n460), .ZN(n459) );
  XNOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(G176GAT), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  INV_X1 U513 ( .A(n565), .ZN(n465) );
  NOR2_X1 U514 ( .A1(n465), .A2(n460), .ZN(n464) );
  XNOR2_X1 U515 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n462) );
  INV_X1 U516 ( .A(G190GAT), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n583), .A2(n465), .ZN(n466) );
  XNOR2_X1 U518 ( .A(n466), .B(KEYINPUT79), .ZN(n467) );
  XNOR2_X1 U519 ( .A(KEYINPUT16), .B(n467), .ZN(n488) );
  XNOR2_X1 U520 ( .A(n530), .B(KEYINPUT27), .ZN(n474) );
  NOR2_X1 U521 ( .A1(n528), .A2(n474), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT97), .B(n468), .Z(n540) );
  XNOR2_X1 U523 ( .A(n477), .B(KEYINPUT66), .ZN(n469) );
  XOR2_X2 U524 ( .A(n469), .B(KEYINPUT28), .Z(n536) );
  INV_X1 U525 ( .A(n536), .ZN(n544) );
  NOR2_X1 U526 ( .A1(n544), .A2(n470), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n540), .A2(n471), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT98), .ZN(n486) );
  NAND2_X1 U529 ( .A1(n477), .A2(n541), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT26), .ZN(n574) );
  NOR2_X1 U531 ( .A1(n574), .A2(n474), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n475), .B(KEYINPUT99), .ZN(n482) );
  XOR2_X1 U533 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n480) );
  NOR2_X1 U534 ( .A1(n541), .A2(n530), .ZN(n476) );
  NOR2_X1 U535 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT100), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U538 ( .A1(n482), .A2(n481), .ZN(n484) );
  NAND2_X1 U539 ( .A1(n484), .A2(n483), .ZN(n485) );
  NAND2_X1 U540 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U541 ( .A(KEYINPUT102), .B(n487), .ZN(n500) );
  AND2_X1 U542 ( .A1(n488), .A2(n500), .ZN(n516) );
  NOR2_X1 U543 ( .A1(n579), .A2(n567), .ZN(n489) );
  XNOR2_X1 U544 ( .A(n489), .B(KEYINPUT74), .ZN(n502) );
  NAND2_X1 U545 ( .A1(n516), .A2(n502), .ZN(n496) );
  NOR2_X1 U546 ( .A1(n528), .A2(n496), .ZN(n490) );
  XOR2_X1 U547 ( .A(G1GAT), .B(n490), .Z(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(n491), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n530), .A2(n496), .ZN(n493) );
  XNOR2_X1 U550 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(G1325GAT) );
  NOR2_X1 U552 ( .A1(n541), .A2(n496), .ZN(n495) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NOR2_X1 U555 ( .A1(n536), .A2(n496), .ZN(n497) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n497), .Z(G1327GAT) );
  NOR2_X1 U557 ( .A1(n498), .A2(n583), .ZN(n499) );
  NAND2_X1 U558 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U559 ( .A(KEYINPUT37), .B(n501), .ZN(n527) );
  NAND2_X1 U560 ( .A1(n502), .A2(n527), .ZN(n503) );
  XNOR2_X1 U561 ( .A(n503), .B(KEYINPUT38), .ZN(n504) );
  XNOR2_X1 U562 ( .A(KEYINPUT104), .B(n504), .ZN(n512) );
  NOR2_X1 U563 ( .A1(n528), .A2(n512), .ZN(n506) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U566 ( .A1(n530), .A2(n512), .ZN(n508) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n508), .B(n507), .ZN(G1329GAT) );
  NOR2_X1 U569 ( .A1(n541), .A2(n512), .ZN(n510) );
  XNOR2_X1 U570 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U572 ( .A(G43GAT), .B(n511), .Z(G1330GAT) );
  NOR2_X1 U573 ( .A1(n536), .A2(n512), .ZN(n514) );
  XNOR2_X1 U574 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n514), .B(n513), .ZN(G1331GAT) );
  NOR2_X1 U576 ( .A1(n515), .A2(n576), .ZN(n526) );
  NAND2_X1 U577 ( .A1(n526), .A2(n516), .ZN(n522) );
  NOR2_X1 U578 ( .A1(n528), .A2(n522), .ZN(n518) );
  XNOR2_X1 U579 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n519), .Z(G1332GAT) );
  NOR2_X1 U582 ( .A1(n530), .A2(n522), .ZN(n520) );
  XOR2_X1 U583 ( .A(G64GAT), .B(n520), .Z(G1333GAT) );
  NOR2_X1 U584 ( .A1(n541), .A2(n522), .ZN(n521) );
  XOR2_X1 U585 ( .A(G71GAT), .B(n521), .Z(G1334GAT) );
  NOR2_X1 U586 ( .A1(n536), .A2(n522), .ZN(n524) );
  XNOR2_X1 U587 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U589 ( .A(G78GAT), .B(n525), .Z(G1335GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n535) );
  NOR2_X1 U591 ( .A1(n528), .A2(n535), .ZN(n529) );
  XOR2_X1 U592 ( .A(G85GAT), .B(n529), .Z(G1336GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n535), .ZN(n531) );
  XOR2_X1 U594 ( .A(G92GAT), .B(n531), .Z(G1337GAT) );
  NOR2_X1 U595 ( .A1(n541), .A2(n535), .ZN(n532) );
  XOR2_X1 U596 ( .A(G99GAT), .B(n532), .Z(G1338GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n534) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n538) );
  NOR2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U601 ( .A(n538), .B(n537), .Z(G1339GAT) );
  NAND2_X1 U602 ( .A1(n539), .A2(n540), .ZN(n556) );
  NOR2_X1 U603 ( .A1(n541), .A2(n556), .ZN(n542) );
  XNOR2_X1 U604 ( .A(n542), .B(KEYINPUT115), .ZN(n543) );
  NOR2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n576), .A2(n552), .ZN(n545) );
  XNOR2_X1 U607 ( .A(n545), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n547) );
  NAND2_X1 U609 ( .A1(n552), .A2(n558), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n550) );
  NAND2_X1 U613 ( .A1(n552), .A2(n583), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n554) );
  NAND2_X1 U617 ( .A1(n552), .A2(n565), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(n555), .ZN(G1343GAT) );
  NOR2_X1 U620 ( .A1(n574), .A2(n556), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n564), .A2(n576), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n560) );
  NAND2_X1 U624 ( .A1(n564), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT53), .Z(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n583), .A2(n564), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n460), .ZN(n568) );
  XOR2_X1 U633 ( .A(G169GAT), .B(n568), .Z(G1348GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n460), .ZN(n570) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n570), .Z(G1350GAT) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT59), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(n572), .Z(n578) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT123), .B(n575), .ZN(n587) );
  INV_X1 U641 ( .A(n587), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n582), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT125), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n589) );
  NOR2_X1 U652 ( .A1(n498), .A2(n587), .ZN(n588) );
  XOR2_X1 U653 ( .A(n589), .B(n588), .Z(G1355GAT) );
endmodule

