

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792;

  XNOR2_X1 U378 ( .A(n488), .B(n465), .ZN(n572) );
  XNOR2_X1 U379 ( .A(n590), .B(KEYINPUT42), .ZN(n792) );
  NOR2_X1 U380 ( .A1(n587), .A2(n586), .ZN(n709) );
  NOR2_X2 U381 ( .A1(n435), .A2(n441), .ZN(n584) );
  XNOR2_X2 U382 ( .A(n513), .B(n449), .ZN(n502) );
  XNOR2_X2 U383 ( .A(n572), .B(n571), .ZN(n618) );
  NOR2_X2 U384 ( .A1(n499), .A2(n566), .ZN(n389) );
  XNOR2_X2 U385 ( .A(n588), .B(KEYINPUT41), .ZN(n706) );
  AND2_X1 U386 ( .A1(n375), .A2(n788), .ZN(n374) );
  NAND2_X1 U387 ( .A1(n425), .A2(n423), .ZN(n634) );
  INV_X1 U388 ( .A(KEYINPUT83), .ZN(n598) );
  AND2_X1 U389 ( .A1(n685), .A2(n684), .ZN(n687) );
  NAND2_X1 U390 ( .A1(n453), .A2(n452), .ZN(n664) );
  XNOR2_X1 U391 ( .A(n417), .B(KEYINPUT35), .ZN(n729) );
  XNOR2_X1 U392 ( .A(n624), .B(n419), .ZN(n418) );
  NAND2_X1 U393 ( .A1(n359), .A2(n432), .ZN(n423) );
  BUF_X1 U394 ( .A(n558), .Z(n611) );
  XNOR2_X1 U395 ( .A(n496), .B(n495), .ZN(n558) );
  BUF_X1 U396 ( .A(n567), .Z(n595) );
  XNOR2_X1 U397 ( .A(n385), .B(n774), .ZN(n659) );
  XNOR2_X1 U398 ( .A(n502), .B(n486), .ZN(n736) );
  XNOR2_X1 U399 ( .A(n387), .B(n386), .ZN(n385) );
  XNOR2_X1 U400 ( .A(n471), .B(KEYINPUT24), .ZN(n386) );
  XNOR2_X1 U401 ( .A(n478), .B(n477), .ZN(n771) );
  XNOR2_X1 U402 ( .A(n433), .B(G134), .ZN(n478) );
  XNOR2_X1 U403 ( .A(G128), .B(G137), .ZN(n474) );
  XNOR2_X1 U404 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n472) );
  XNOR2_X1 U405 ( .A(G902), .B(KEYINPUT15), .ZN(n655) );
  INV_X2 U406 ( .A(G953), .ZN(n480) );
  NAND2_X1 U407 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U408 ( .A(n476), .B(n357), .ZN(n387) );
  XNOR2_X1 U409 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U410 ( .A(n607), .B(n399), .ZN(n398) );
  XNOR2_X1 U411 ( .A(n413), .B(G146), .ZN(n510) );
  INV_X1 U412 ( .A(G125), .ZN(n413) );
  AND2_X1 U413 ( .A1(n618), .A2(n617), .ZN(n635) );
  AND2_X1 U414 ( .A1(n428), .A2(n426), .ZN(n425) );
  NOR2_X1 U415 ( .A1(G902), .A2(n736), .ZN(n488) );
  XNOR2_X1 U416 ( .A(n591), .B(KEYINPUT46), .ZN(n380) );
  AND2_X1 U417 ( .A1(n410), .A2(n751), .ZN(n580) );
  XNOR2_X1 U418 ( .A(n412), .B(n411), .ZN(n410) );
  INV_X1 U419 ( .A(KEYINPUT47), .ZN(n411) );
  XNOR2_X1 U420 ( .A(n615), .B(KEYINPUT86), .ZN(n630) );
  NAND2_X1 U421 ( .A1(n664), .A2(n663), .ZN(n615) );
  INV_X1 U422 ( .A(KEYINPUT71), .ZN(n433) );
  INV_X1 U423 ( .A(KEYINPUT4), .ZN(n479) );
  XNOR2_X1 U424 ( .A(G122), .B(G113), .ZN(n550) );
  NAND2_X1 U425 ( .A1(n462), .A2(n367), .ZN(n429) );
  NAND2_X1 U426 ( .A1(n395), .A2(n394), .ZN(n393) );
  AND2_X1 U427 ( .A1(n423), .A2(n425), .ZN(n395) );
  INV_X1 U428 ( .A(n608), .ZN(n397) );
  NOR2_X1 U429 ( .A1(n396), .A2(n398), .ZN(n391) );
  INV_X1 U430 ( .A(n423), .ZN(n396) );
  INV_X1 U431 ( .A(n606), .ZN(n402) );
  INV_X1 U432 ( .A(G902), .ZN(n554) );
  XNOR2_X1 U433 ( .A(n502), .B(n448), .ZN(n666) );
  XNOR2_X1 U434 ( .A(n506), .B(n501), .ZN(n448) );
  XNOR2_X1 U435 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n509) );
  NAND2_X1 U436 ( .A1(n360), .A2(G953), .ZN(n400) );
  NAND2_X1 U437 ( .A1(n440), .A2(n439), .ZN(n438) );
  AND2_X1 U438 ( .A1(n445), .A2(n443), .ZN(n439) );
  INV_X1 U439 ( .A(n565), .ZN(n440) );
  NAND2_X1 U440 ( .A1(n444), .A2(n442), .ZN(n441) );
  OR2_X1 U441 ( .A1(n445), .A2(n443), .ZN(n442) );
  NAND2_X1 U442 ( .A1(n565), .A2(n582), .ZN(n444) );
  INV_X1 U443 ( .A(KEYINPUT32), .ZN(n457) );
  OR2_X1 U444 ( .A1(n610), .A2(n457), .ZN(n456) );
  AND2_X1 U445 ( .A1(n414), .A2(n559), .ZN(n589) );
  XNOR2_X1 U446 ( .A(n416), .B(n415), .ZN(n414) );
  INV_X1 U447 ( .A(KEYINPUT28), .ZN(n415) );
  NAND2_X1 U448 ( .A1(n614), .A2(n619), .ZN(n632) );
  INV_X1 U449 ( .A(n630), .ZN(n405) );
  NAND2_X1 U450 ( .A1(n580), .A2(n579), .ZN(n381) );
  NAND2_X1 U451 ( .A1(n380), .A2(KEYINPUT48), .ZN(n377) );
  NOR2_X1 U452 ( .A1(n616), .A2(KEYINPUT85), .ZN(n627) );
  XNOR2_X1 U453 ( .A(G116), .B(G113), .ZN(n500) );
  XNOR2_X1 U454 ( .A(n510), .B(n467), .ZN(n546) );
  INV_X1 U455 ( .A(KEYINPUT10), .ZN(n467) );
  XNOR2_X1 U456 ( .A(KEYINPUT3), .B(G119), .ZN(n517) );
  XNOR2_X1 U457 ( .A(G116), .B(G107), .ZN(n533) );
  XNOR2_X1 U458 ( .A(n403), .B(n365), .ZN(n489) );
  XNOR2_X1 U459 ( .A(KEYINPUT75), .B(KEYINPUT14), .ZN(n403) );
  OR2_X1 U460 ( .A1(G902), .A2(G237), .ZN(n523) );
  NOR2_X1 U461 ( .A1(n708), .A2(n707), .ZN(n712) );
  AND2_X1 U462 ( .A1(n585), .A2(n446), .ZN(n445) );
  INV_X1 U463 ( .A(n566), .ZN(n446) );
  XNOR2_X1 U464 ( .A(n494), .B(KEYINPUT25), .ZN(n495) );
  NAND2_X1 U465 ( .A1(n659), .A2(n554), .ZN(n496) );
  XNOR2_X1 U466 ( .A(n546), .B(n468), .ZN(n774) );
  INV_X1 U467 ( .A(n483), .ZN(n468) );
  XNOR2_X1 U468 ( .A(G110), .B(G119), .ZN(n469) );
  XNOR2_X1 U469 ( .A(G122), .B(G134), .ZN(n529) );
  NOR2_X1 U470 ( .A1(G237), .A2(G953), .ZN(n503) );
  XNOR2_X1 U471 ( .A(G143), .B(G104), .ZN(n548) );
  INV_X1 U472 ( .A(n546), .ZN(n409) );
  XNOR2_X1 U473 ( .A(G131), .B(KEYINPUT12), .ZN(n542) );
  XOR2_X1 U474 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n543) );
  XNOR2_X1 U475 ( .A(n771), .B(n450), .ZN(n449) );
  INV_X1 U476 ( .A(G146), .ZN(n450) );
  INV_X1 U477 ( .A(G107), .ZN(n481) );
  XNOR2_X1 U478 ( .A(G110), .B(G104), .ZN(n515) );
  XNOR2_X1 U479 ( .A(n623), .B(n622), .ZN(n716) );
  NAND2_X1 U480 ( .A1(n716), .A2(n639), .ZN(n624) );
  INV_X1 U481 ( .A(KEYINPUT34), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n540), .B(n539), .ZN(n568) );
  XNOR2_X1 U483 ( .A(n556), .B(n555), .ZN(n587) );
  NAND2_X1 U484 ( .A1(n392), .A2(n390), .ZN(n614) );
  NAND2_X1 U485 ( .A1(n391), .A2(n364), .ZN(n390) );
  AND2_X2 U486 ( .A1(n657), .A2(n466), .ZN(n733) );
  XNOR2_X1 U487 ( .A(n407), .B(n765), .ZN(n679) );
  XNOR2_X1 U488 ( .A(n513), .B(n514), .ZN(n407) );
  NOR2_X1 U489 ( .A1(n480), .A2(G952), .ZN(n739) );
  NAND2_X1 U490 ( .A1(n384), .A2(n368), .ZN(n383) );
  INV_X1 U491 ( .A(KEYINPUT120), .ZN(n401) );
  NAND2_X1 U492 ( .A1(n436), .A2(n438), .ZN(n600) );
  INV_X1 U493 ( .A(n441), .ZN(n436) );
  NAND2_X1 U494 ( .A1(n438), .A2(n437), .ZN(n435) );
  NAND2_X1 U495 ( .A1(n455), .A2(n454), .ZN(n452) );
  AND2_X1 U496 ( .A1(n458), .A2(n456), .ZN(n453) );
  AND2_X1 U497 ( .A1(n610), .A2(n457), .ZN(n454) );
  NAND2_X1 U498 ( .A1(n589), .A2(n358), .ZN(n388) );
  AND2_X1 U499 ( .A1(n580), .A2(n366), .ZN(n356) );
  XOR2_X1 U500 ( .A(n475), .B(n474), .Z(n357) );
  AND2_X1 U501 ( .A1(n432), .A2(n431), .ZN(n358) );
  AND2_X1 U502 ( .A1(n431), .A2(n424), .ZN(n359) );
  OR2_X1 U503 ( .A1(n723), .A2(n721), .ZN(n360) );
  AND2_X1 U504 ( .A1(n573), .A2(n463), .ZN(n361) );
  AND2_X1 U505 ( .A1(n383), .A2(n382), .ZN(n362) );
  INV_X1 U506 ( .A(n707), .ZN(n463) );
  XNOR2_X1 U507 ( .A(n561), .B(n560), .ZN(n638) );
  XOR2_X1 U508 ( .A(KEYINPUT90), .B(n490), .Z(n363) );
  AND2_X1 U509 ( .A1(n425), .A2(n608), .ZN(n364) );
  AND2_X1 U510 ( .A1(G234), .A2(G237), .ZN(n365) );
  AND2_X1 U511 ( .A1(n579), .A2(n373), .ZN(n366) );
  OR2_X1 U512 ( .A1(n463), .A2(n461), .ZN(n367) );
  AND2_X1 U513 ( .A1(n400), .A2(n401), .ZN(n368) );
  AND2_X1 U514 ( .A1(n727), .A2(n726), .ZN(n369) );
  INV_X1 U515 ( .A(n741), .ZN(n437) );
  OR2_X1 U516 ( .A1(KEYINPUT85), .A2(KEYINPUT44), .ZN(n370) );
  NAND2_X1 U517 ( .A1(n371), .A2(n618), .ZN(n578) );
  XNOR2_X1 U518 ( .A(n577), .B(n576), .ZN(n371) );
  AND2_X1 U519 ( .A1(n629), .A2(KEYINPUT44), .ZN(n406) );
  NAND2_X1 U520 ( .A1(n393), .A2(n397), .ZN(n392) );
  AND2_X1 U521 ( .A1(n372), .A2(n656), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n688), .A2(n372), .ZN(n690) );
  NAND2_X1 U523 ( .A1(n654), .A2(n451), .ZN(n372) );
  INV_X1 U524 ( .A(KEYINPUT48), .ZN(n373) );
  NAND2_X2 U525 ( .A1(n376), .A2(n374), .ZN(n434) );
  NAND2_X1 U526 ( .A1(n381), .A2(KEYINPUT48), .ZN(n375) );
  AND2_X2 U527 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U528 ( .A1(n356), .A2(n379), .ZN(n378) );
  INV_X1 U529 ( .A(n380), .ZN(n379) );
  NAND2_X1 U530 ( .A1(n722), .A2(n369), .ZN(n382) );
  NAND2_X1 U531 ( .A1(n722), .A2(n360), .ZN(n384) );
  NAND2_X1 U532 ( .A1(n753), .A2(n711), .ZN(n412) );
  XNOR2_X2 U533 ( .A(n388), .B(KEYINPUT79), .ZN(n753) );
  NAND2_X1 U534 ( .A1(n389), .A2(n573), .ZN(n416) );
  NAND2_X1 U535 ( .A1(n574), .A2(n389), .ZN(n592) );
  INV_X1 U536 ( .A(n398), .ZN(n394) );
  INV_X1 U537 ( .A(KEYINPUT105), .ZN(n399) );
  NOR2_X1 U538 ( .A1(n421), .A2(n430), .ZN(n420) );
  INV_X1 U539 ( .A(n429), .ZN(n432) );
  NOR2_X2 U540 ( .A1(n558), .A2(n402), .ZN(n617) );
  NAND2_X1 U541 ( .A1(n559), .A2(n617), .ZN(n561) );
  NOR2_X1 U542 ( .A1(n459), .A2(n604), .ZN(n421) );
  INV_X1 U543 ( .A(n604), .ZN(n427) );
  NAND2_X1 U544 ( .A1(n418), .A2(n626), .ZN(n417) );
  NAND2_X1 U545 ( .A1(n404), .A2(n370), .ZN(n645) );
  NAND2_X1 U546 ( .A1(n406), .A2(n405), .ZN(n404) );
  NAND2_X1 U547 ( .A1(n429), .A2(n605), .ZN(n428) );
  INV_X1 U548 ( .A(n617), .ZN(n693) );
  NAND2_X1 U549 ( .A1(n567), .A2(n527), .ZN(n462) );
  XNOR2_X2 U550 ( .A(n464), .B(n522), .ZN(n567) );
  XNOR2_X1 U551 ( .A(n408), .B(n547), .ZN(n672) );
  XNOR2_X1 U552 ( .A(n553), .B(n409), .ZN(n408) );
  NAND2_X1 U553 ( .A1(n567), .A2(n427), .ZN(n422) );
  NAND2_X1 U554 ( .A1(n460), .A2(n459), .ZN(n431) );
  NAND2_X1 U555 ( .A1(n422), .A2(n420), .ZN(n426) );
  NOR2_X1 U556 ( .A1(n604), .A2(n605), .ZN(n424) );
  INV_X1 U557 ( .A(n605), .ZN(n430) );
  XNOR2_X2 U558 ( .A(n434), .B(n598), .ZN(n653) );
  INV_X1 U559 ( .A(n582), .ZN(n443) );
  NOR2_X1 U560 ( .A1(n565), .A2(n566), .ZN(n581) );
  NAND2_X1 U561 ( .A1(n447), .A2(n611), .ZN(n612) );
  INV_X1 U562 ( .A(n573), .ZN(n447) );
  XNOR2_X2 U563 ( .A(n772), .B(G101), .ZN(n513) );
  NAND2_X1 U564 ( .A1(n451), .A2(n480), .ZN(n763) );
  INV_X1 U565 ( .A(n685), .ZN(n451) );
  INV_X1 U566 ( .A(n632), .ZN(n455) );
  NAND2_X1 U567 ( .A1(n632), .A2(KEYINPUT32), .ZN(n458) );
  NAND2_X1 U568 ( .A1(n460), .A2(n463), .ZN(n575) );
  NOR2_X1 U569 ( .A1(n707), .A2(n527), .ZN(n459) );
  INV_X1 U570 ( .A(n567), .ZN(n460) );
  INV_X1 U571 ( .A(n527), .ZN(n461) );
  NAND2_X1 U572 ( .A1(n679), .A2(n655), .ZN(n464) );
  XOR2_X1 U573 ( .A(n487), .B(KEYINPUT72), .Z(n465) );
  INV_X1 U574 ( .A(KEYINPUT82), .ZN(n686) );
  INV_X1 U575 ( .A(n572), .ZN(n559) );
  XNOR2_X1 U576 ( .A(n517), .B(n500), .ZN(n501) );
  XNOR2_X1 U577 ( .A(n482), .B(n481), .ZN(n484) );
  INV_X1 U578 ( .A(KEYINPUT95), .ZN(n560) );
  XNOR2_X1 U579 ( .A(n505), .B(n504), .ZN(n506) );
  INV_X1 U580 ( .A(KEYINPUT110), .ZN(n562) );
  XNOR2_X1 U581 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U582 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U583 ( .A(G140), .B(KEYINPUT70), .Z(n483) );
  XOR2_X1 U584 ( .A(KEYINPUT74), .B(KEYINPUT92), .Z(n470) );
  XNOR2_X1 U585 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U586 ( .A1(n480), .A2(G234), .ZN(n473) );
  XNOR2_X1 U587 ( .A(n473), .B(n472), .ZN(n532) );
  AND2_X1 U588 ( .A1(n532), .A2(G221), .ZN(n476) );
  XOR2_X1 U589 ( .A(KEYINPUT23), .B(KEYINPUT93), .Z(n475) );
  XNOR2_X1 U590 ( .A(G137), .B(G131), .ZN(n477) );
  XOR2_X2 U591 ( .A(G143), .B(G128), .Z(n528) );
  XNOR2_X2 U592 ( .A(n528), .B(n479), .ZN(n772) );
  NAND2_X1 U593 ( .A1(G227), .A2(n480), .ZN(n482) );
  XNOR2_X1 U594 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U595 ( .A(n485), .B(n515), .ZN(n486) );
  XNOR2_X1 U596 ( .A(G469), .B(KEYINPUT73), .ZN(n487) );
  AND2_X1 U597 ( .A1(n489), .A2(G952), .ZN(n724) );
  AND2_X1 U598 ( .A1(n724), .A2(n480), .ZN(n720) );
  NAND2_X1 U599 ( .A1(G902), .A2(n489), .ZN(n490) );
  NAND2_X1 U600 ( .A1(G953), .A2(n363), .ZN(n602) );
  XNOR2_X1 U601 ( .A(KEYINPUT108), .B(n602), .ZN(n491) );
  NOR2_X1 U602 ( .A1(G900), .A2(n491), .ZN(n492) );
  NOR2_X1 U603 ( .A1(n720), .A2(n492), .ZN(n566) );
  NAND2_X1 U604 ( .A1(G234), .A2(n655), .ZN(n493) );
  XNOR2_X1 U605 ( .A(KEYINPUT20), .B(n493), .ZN(n497) );
  NAND2_X1 U606 ( .A1(G217), .A2(n497), .ZN(n494) );
  NAND2_X1 U607 ( .A1(n497), .A2(G221), .ZN(n498) );
  XOR2_X1 U608 ( .A(KEYINPUT21), .B(n498), .Z(n697) );
  NAND2_X1 U609 ( .A1(n611), .A2(n697), .ZN(n499) );
  XNOR2_X1 U610 ( .A(n503), .B(KEYINPUT76), .ZN(n541) );
  AND2_X1 U611 ( .A1(n541), .A2(G210), .ZN(n505) );
  XOR2_X1 U612 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n504) );
  NAND2_X1 U613 ( .A1(n666), .A2(n554), .ZN(n507) );
  XNOR2_X2 U614 ( .A(n507), .B(G472), .ZN(n573) );
  NAND2_X1 U615 ( .A1(n480), .A2(G224), .ZN(n508) );
  XNOR2_X1 U616 ( .A(n508), .B(KEYINPUT78), .ZN(n512) );
  XNOR2_X1 U617 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U618 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X1 U619 ( .A(n533), .B(KEYINPUT16), .ZN(n516) );
  XNOR2_X1 U620 ( .A(n516), .B(n515), .ZN(n519) );
  XNOR2_X1 U621 ( .A(n517), .B(n550), .ZN(n518) );
  XNOR2_X1 U622 ( .A(n519), .B(n518), .ZN(n765) );
  NAND2_X1 U623 ( .A1(n523), .A2(G210), .ZN(n521) );
  XNOR2_X1 U624 ( .A(KEYINPUT80), .B(KEYINPUT88), .ZN(n520) );
  NAND2_X1 U625 ( .A1(n523), .A2(G214), .ZN(n524) );
  XNOR2_X1 U626 ( .A(n524), .B(KEYINPUT89), .ZN(n707) );
  XNOR2_X1 U627 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n526) );
  INV_X1 U628 ( .A(KEYINPUT67), .ZN(n525) );
  XNOR2_X1 U629 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U630 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n530) );
  XNOR2_X1 U631 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U632 ( .A(n528), .B(n531), .ZN(n538) );
  AND2_X1 U633 ( .A1(n532), .A2(G217), .ZN(n536) );
  XOR2_X1 U634 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n534) );
  XNOR2_X1 U635 ( .A(n538), .B(n537), .ZN(n731) );
  NAND2_X1 U636 ( .A1(n731), .A2(n554), .ZN(n540) );
  INV_X1 U637 ( .A(G478), .ZN(n539) );
  NAND2_X1 U638 ( .A1(n541), .A2(G214), .ZN(n545) );
  XNOR2_X1 U639 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U640 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n549) );
  XNOR2_X1 U642 ( .A(n549), .B(n548), .ZN(n552) );
  XNOR2_X1 U643 ( .A(n550), .B(G140), .ZN(n551) );
  XNOR2_X1 U644 ( .A(n552), .B(n551), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n672), .A2(n554), .ZN(n556) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(G475), .Z(n555) );
  NOR2_X1 U647 ( .A1(n568), .A2(n587), .ZN(n557) );
  XOR2_X1 U648 ( .A(n557), .B(KEYINPUT103), .Z(n756) );
  XOR2_X1 U649 ( .A(KEYINPUT104), .B(n756), .Z(n599) );
  NAND2_X1 U650 ( .A1(n587), .A2(n568), .ZN(n741) );
  NAND2_X1 U651 ( .A1(n599), .A2(n741), .ZN(n711) );
  XNOR2_X1 U652 ( .A(KEYINPUT94), .B(n697), .ZN(n606) );
  XNOR2_X1 U653 ( .A(n638), .B(n562), .ZN(n564) );
  XNOR2_X1 U654 ( .A(KEYINPUT30), .B(n361), .ZN(n563) );
  INV_X1 U655 ( .A(n568), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n625) );
  NOR2_X1 U657 ( .A1(n595), .A2(n625), .ZN(n569) );
  NAND2_X1 U658 ( .A1(n581), .A2(n569), .ZN(n751) );
  INV_X1 U659 ( .A(KEYINPUT66), .ZN(n570) );
  XNOR2_X1 U660 ( .A(n570), .B(KEYINPUT1), .ZN(n571) );
  XNOR2_X1 U661 ( .A(n573), .B(KEYINPUT6), .ZN(n619) );
  NOR2_X1 U662 ( .A1(n741), .A2(n619), .ZN(n574) );
  NOR2_X1 U663 ( .A1(n592), .A2(n575), .ZN(n577) );
  XNOR2_X1 U664 ( .A(KEYINPUT112), .B(KEYINPUT36), .ZN(n576) );
  XNOR2_X1 U665 ( .A(n578), .B(KEYINPUT113), .ZN(n784) );
  INV_X1 U666 ( .A(n784), .ZN(n579) );
  XNOR2_X1 U667 ( .A(n595), .B(KEYINPUT38), .ZN(n585) );
  XOR2_X1 U668 ( .A(KEYINPUT84), .B(KEYINPUT39), .Z(n582) );
  XNOR2_X1 U669 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n584), .B(n583), .ZN(n789) );
  INV_X1 U671 ( .A(n585), .ZN(n708) );
  NAND2_X1 U672 ( .A1(n712), .A2(n709), .ZN(n588) );
  NAND2_X1 U673 ( .A1(n589), .A2(n706), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n789), .A2(n792), .ZN(n591) );
  OR2_X1 U675 ( .A1(n618), .A2(n592), .ZN(n593) );
  NOR2_X1 U676 ( .A1(n707), .A2(n593), .ZN(n594) );
  XNOR2_X1 U677 ( .A(n594), .B(KEYINPUT43), .ZN(n596) );
  NOR2_X1 U678 ( .A1(n596), .A2(n460), .ZN(n597) );
  XNOR2_X1 U679 ( .A(n597), .B(KEYINPUT109), .ZN(n788) );
  INV_X1 U680 ( .A(n653), .ZN(n601) );
  OR2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n759) );
  NAND2_X2 U682 ( .A1(n601), .A2(n759), .ZN(n778) );
  NOR2_X1 U683 ( .A1(n602), .A2(G898), .ZN(n603) );
  NOR2_X1 U684 ( .A1(n603), .A2(n720), .ZN(n604) );
  XNOR2_X1 U685 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n709), .A2(n606), .ZN(n607) );
  XOR2_X1 U687 ( .A(KEYINPUT65), .B(KEYINPUT22), .Z(n608) );
  INV_X1 U688 ( .A(n618), .ZN(n694) );
  INV_X1 U689 ( .A(KEYINPUT106), .ZN(n609) );
  XNOR2_X1 U690 ( .A(n611), .B(n609), .ZN(n696) );
  NOR2_X1 U691 ( .A1(n694), .A2(n696), .ZN(n610) );
  NOR2_X1 U692 ( .A1(n618), .A2(n612), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n663) );
  NOR2_X1 U694 ( .A1(n630), .A2(KEYINPUT44), .ZN(n616) );
  INV_X1 U695 ( .A(n619), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n635), .A2(n620), .ZN(n623) );
  INV_X1 U697 ( .A(KEYINPUT87), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n621), .B(KEYINPUT33), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n634), .B(KEYINPUT91), .ZN(n639) );
  INV_X1 U700 ( .A(n625), .ZN(n626) );
  NOR2_X1 U701 ( .A1(n627), .A2(n729), .ZN(n647) );
  INV_X1 U702 ( .A(KEYINPUT85), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n729), .A2(n628), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n694), .A2(n696), .ZN(n631) );
  NOR2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U706 ( .A(KEYINPUT107), .B(n633), .Z(n787) );
  XOR2_X1 U707 ( .A(KEYINPUT31), .B(KEYINPUT97), .Z(n637) );
  NAND2_X1 U708 ( .A1(n635), .A2(n573), .ZN(n702) );
  NOR2_X1 U709 ( .A1(n634), .A2(n702), .ZN(n636) );
  XOR2_X1 U710 ( .A(n637), .B(n636), .Z(n757) );
  NOR2_X1 U711 ( .A1(n638), .A2(n573), .ZN(n640) );
  AND2_X1 U712 ( .A1(n640), .A2(n639), .ZN(n743) );
  NOR2_X1 U713 ( .A1(n757), .A2(n743), .ZN(n642) );
  INV_X1 U714 ( .A(n711), .ZN(n641) );
  NOR2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U716 ( .A1(n787), .A2(n643), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n649) );
  XNOR2_X1 U719 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n685) );
  NOR2_X1 U721 ( .A1(n778), .A2(n685), .ZN(n650) );
  OR2_X1 U722 ( .A1(n650), .A2(KEYINPUT2), .ZN(n657) );
  NAND2_X1 U723 ( .A1(n759), .A2(KEYINPUT2), .ZN(n651) );
  XOR2_X1 U724 ( .A(KEYINPUT81), .B(n651), .Z(n652) );
  NOR2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  INV_X1 U726 ( .A(n655), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n733), .A2(G217), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n661) );
  INV_X1 U729 ( .A(n739), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT123), .ZN(G66) );
  XNOR2_X1 U732 ( .A(n663), .B(G110), .ZN(G12) );
  XNOR2_X1 U733 ( .A(n664), .B(G119), .ZN(G21) );
  NAND2_X1 U734 ( .A1(n733), .A2(G472), .ZN(n668) );
  XOR2_X1 U735 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n665) );
  XNOR2_X1 U736 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X2 U738 ( .A1(n669), .A2(n739), .ZN(n671) );
  XNOR2_X1 U739 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(G57) );
  NAND2_X1 U741 ( .A1(n733), .A2(G475), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n672), .B(KEYINPUT59), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X2 U744 ( .A1(n675), .A2(n739), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n676), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U746 ( .A1(n733), .A2(G210), .ZN(n681) );
  XOR2_X1 U747 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n677) );
  XNOR2_X1 U748 ( .A(n677), .B(KEYINPUT55), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X2 U751 ( .A1(n682), .A2(n739), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n683), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U753 ( .A(KEYINPUT53), .ZN(n728) );
  INV_X1 U754 ( .A(KEYINPUT2), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n687), .B(n686), .ZN(n688) );
  AND2_X1 U756 ( .A1(n778), .A2(n684), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n692) );
  AND2_X1 U758 ( .A1(n716), .A2(n706), .ZN(n691) );
  NOR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n722) );
  NAND2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U761 ( .A(n695), .B(KEYINPUT50), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U763 ( .A(KEYINPUT49), .B(n698), .Z(n699) );
  NOR2_X1 U764 ( .A1(n573), .A2(n699), .ZN(n700) );
  NAND2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U767 ( .A(KEYINPUT51), .B(n704), .Z(n705) );
  NAND2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n718) );
  NAND2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U772 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U774 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U775 ( .A(KEYINPUT52), .B(n719), .Z(n723) );
  INV_X1 U776 ( .A(n720), .ZN(n721) );
  INV_X1 U777 ( .A(n723), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n725), .A2(n724), .ZN(n727) );
  AND2_X1 U779 ( .A1(n480), .A2(KEYINPUT120), .ZN(n726) );
  XNOR2_X1 U780 ( .A(n728), .B(n362), .ZN(G75) );
  XOR2_X1 U781 ( .A(G122), .B(n729), .Z(G24) );
  NAND2_X1 U782 ( .A1(n733), .A2(G478), .ZN(n730) );
  XOR2_X1 U783 ( .A(n731), .B(n730), .Z(n732) );
  NOR2_X1 U784 ( .A1(n732), .A2(n739), .ZN(G63) );
  NAND2_X1 U785 ( .A1(n733), .A2(G469), .ZN(n738) );
  XOR2_X1 U786 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n734) );
  XNOR2_X1 U787 ( .A(n734), .B(KEYINPUT58), .ZN(n735) );
  XNOR2_X1 U788 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U789 ( .A(n738), .B(n737), .ZN(n740) );
  NOR2_X1 U790 ( .A1(n740), .A2(n739), .ZN(G54) );
  NAND2_X1 U791 ( .A1(n437), .A2(n743), .ZN(n742) );
  XNOR2_X1 U792 ( .A(G104), .B(n742), .ZN(G6) );
  NAND2_X1 U793 ( .A1(n743), .A2(n756), .ZN(n744) );
  XNOR2_X1 U794 ( .A(n744), .B(KEYINPUT27), .ZN(n745) );
  XOR2_X1 U795 ( .A(n745), .B(KEYINPUT116), .Z(n747) );
  XNOR2_X1 U796 ( .A(G107), .B(KEYINPUT26), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n747), .B(n746), .ZN(G9) );
  XOR2_X1 U798 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n749) );
  NAND2_X1 U799 ( .A1(n753), .A2(n756), .ZN(n748) );
  XNOR2_X1 U800 ( .A(n749), .B(n748), .ZN(n750) );
  XOR2_X1 U801 ( .A(G128), .B(n750), .Z(G30) );
  XNOR2_X1 U802 ( .A(G143), .B(KEYINPUT118), .ZN(n752) );
  XNOR2_X1 U803 ( .A(n752), .B(n751), .ZN(G45) );
  NAND2_X1 U804 ( .A1(n753), .A2(n437), .ZN(n754) );
  XNOR2_X1 U805 ( .A(n754), .B(G146), .ZN(G48) );
  NAND2_X1 U806 ( .A1(n757), .A2(n437), .ZN(n755) );
  XNOR2_X1 U807 ( .A(n755), .B(G113), .ZN(G15) );
  NAND2_X1 U808 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U809 ( .A(n758), .B(G116), .ZN(G18) );
  XNOR2_X1 U810 ( .A(G134), .B(n759), .ZN(G36) );
  NAND2_X1 U811 ( .A1(G953), .A2(G224), .ZN(n760) );
  XNOR2_X1 U812 ( .A(KEYINPUT61), .B(n760), .ZN(n761) );
  NAND2_X1 U813 ( .A1(n761), .A2(G898), .ZN(n762) );
  NAND2_X1 U814 ( .A1(n763), .A2(n762), .ZN(n769) );
  XNOR2_X1 U815 ( .A(G101), .B(KEYINPUT124), .ZN(n764) );
  XNOR2_X1 U816 ( .A(n765), .B(n764), .ZN(n767) );
  NOR2_X1 U817 ( .A1(G898), .A2(n480), .ZN(n766) );
  NOR2_X1 U818 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n769), .B(n768), .ZN(n770) );
  XOR2_X1 U820 ( .A(KEYINPUT125), .B(n770), .Z(G69) );
  XOR2_X1 U821 ( .A(n772), .B(n771), .Z(n773) );
  XOR2_X1 U822 ( .A(n774), .B(n773), .Z(n780) );
  XOR2_X1 U823 ( .A(G227), .B(n780), .Z(n775) );
  NAND2_X1 U824 ( .A1(n775), .A2(G900), .ZN(n776) );
  NAND2_X1 U825 ( .A1(G953), .A2(n776), .ZN(n777) );
  XNOR2_X1 U826 ( .A(n777), .B(KEYINPUT126), .ZN(n783) );
  INV_X1 U827 ( .A(n778), .ZN(n779) );
  XNOR2_X1 U828 ( .A(n780), .B(n779), .ZN(n781) );
  NAND2_X1 U829 ( .A1(n781), .A2(n480), .ZN(n782) );
  NAND2_X1 U830 ( .A1(n783), .A2(n782), .ZN(G72) );
  XOR2_X1 U831 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n786) );
  XNOR2_X1 U832 ( .A(G125), .B(n784), .ZN(n785) );
  XNOR2_X1 U833 ( .A(n786), .B(n785), .ZN(G27) );
  XOR2_X1 U834 ( .A(G101), .B(n787), .Z(G3) );
  XNOR2_X1 U835 ( .A(G140), .B(n788), .ZN(G42) );
  BUF_X1 U836 ( .A(n789), .Z(n790) );
  XOR2_X1 U837 ( .A(n790), .B(G131), .Z(n791) );
  XNOR2_X1 U838 ( .A(KEYINPUT127), .B(n791), .ZN(G33) );
  XNOR2_X1 U839 ( .A(n792), .B(G137), .ZN(G39) );
endmodule

