//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT64), .A2(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n195), .B1(G143), .B2(new_n187), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n191), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n195), .A3(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G137), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n203), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n202), .A2(G137), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n204), .A2(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(G131), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n208), .A2(new_n211), .A3(KEYINPUT67), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT67), .B1(new_n208), .B2(new_n211), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n200), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n188), .A2(new_n190), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT0), .B(G128), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n198), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n217), .A2(new_n218), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n218), .B1(new_n217), .B2(new_n223), .ZN(new_n225));
  OAI211_X1 g039(.A(KEYINPUT30), .B(new_n214), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n217), .A2(new_n223), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT64), .B(G128), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n198), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AND4_X1   g045(.A1(new_n195), .A2(new_n188), .A3(new_n190), .A4(G128), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n208), .B(new_n211), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT30), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n227), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n217), .A2(new_n218), .A3(new_n223), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n240), .A2(new_n227), .A3(KEYINPUT30), .A4(new_n214), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G119), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT65), .B1(new_n243), .B2(G116), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n245));
  INV_X1    g059(.A(G116), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G119), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n244), .A2(new_n247), .B1(G116), .B2(new_n243), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT2), .B(G113), .Z(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n242), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n250), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n252), .B(new_n214), .C1(new_n224), .C2(new_n225), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n240), .A2(new_n255), .A3(new_n252), .A4(new_n214), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(G237), .A2(G953), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G210), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n259), .B(KEYINPUT27), .Z(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n251), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT31), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n242), .A2(new_n250), .B1(new_n256), .B2(new_n254), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT31), .A3(new_n263), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n252), .A2(new_n228), .ZN(new_n270));
  INV_X1    g084(.A(new_n214), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n254), .A2(new_n256), .B1(new_n250), .B2(new_n234), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n269), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n266), .A2(new_n268), .B1(new_n274), .B2(new_n262), .ZN(new_n275));
  NOR2_X1   g089(.A1(G472), .A2(G902), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT70), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n262), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n252), .B1(new_n237), .B2(new_n241), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n254), .A2(new_n256), .ZN(new_n282));
  NOR4_X1   g096(.A1(new_n281), .A2(new_n282), .A3(new_n265), .A4(new_n262), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT31), .B1(new_n267), .B2(new_n263), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n276), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n278), .A2(new_n279), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n266), .A2(new_n268), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n277), .B1(new_n289), .B2(new_n280), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT32), .ZN(new_n291));
  INV_X1    g105(.A(new_n272), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n240), .A2(new_n214), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n250), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n257), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n292), .B1(new_n295), .B2(KEYINPUT28), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT29), .A3(new_n263), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n272), .B(new_n263), .C1(new_n273), .C2(new_n269), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n262), .B1(new_n281), .B2(new_n282), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G472), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n288), .A2(new_n291), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G140), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(KEYINPUT71), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(G125), .A3(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(KEYINPUT16), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(G125), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT16), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n187), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n311), .A2(new_n187), .A3(new_n314), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n311), .A2(new_n314), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT72), .A3(new_n187), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n322));
  INV_X1    g136(.A(G128), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT23), .B1(new_n323), .B2(G119), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(G119), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n194), .B2(G119), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT24), .B(G110), .Z(new_n329));
  AOI22_X1  g143(.A1(new_n327), .A2(G110), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n321), .A2(new_n330), .ZN(new_n331));
  OAI22_X1  g145(.A1(new_n327), .A2(G110), .B1(new_n328), .B2(new_n329), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n307), .A2(G140), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n312), .A2(new_n333), .A3(new_n187), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n332), .B(new_n334), .C1(new_n187), .C2(new_n319), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G137), .ZN(new_n337));
  INV_X1    g151(.A(G953), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n338), .A2(G221), .A3(G234), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n337), .B(new_n339), .Z(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n331), .A2(new_n335), .A3(new_n340), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n298), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n342), .A2(KEYINPUT25), .A3(new_n298), .A4(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G217), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G234), .B2(new_n298), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n342), .A2(new_n343), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(G902), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n348), .A2(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G210), .B1(G237), .B2(G902), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT76), .ZN(new_n355));
  INV_X1    g169(.A(G104), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT3), .B1(new_n356), .B2(G107), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n358));
  INV_X1    g172(.A(G107), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(G104), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(G107), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G101), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT73), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n362), .A2(new_n366), .A3(new_n363), .A4(G101), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(G101), .ZN(new_n369));
  INV_X1    g183(.A(G101), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n357), .A2(new_n360), .A3(new_n370), .A4(new_n361), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(KEYINPUT4), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n250), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT5), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n243), .A3(G116), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G113), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n248), .B2(KEYINPUT5), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n248), .A2(new_n249), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n356), .A2(G107), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n359), .A2(G104), .ZN(new_n381));
  OAI21_X1  g195(.A(G101), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n371), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n378), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n373), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n373), .A2(new_n387), .A3(new_n385), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n222), .A2(G125), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n200), .B2(G125), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n338), .A2(G224), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n393), .B(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n386), .A2(new_n397), .A3(new_n388), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n391), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n393), .B1(new_n401), .B2(new_n395), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n395), .A2(new_n401), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n392), .B(new_n403), .C1(new_n200), .C2(G125), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n387), .B(KEYINPUT8), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n379), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n383), .B1(new_n408), .B2(new_n377), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n385), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n400), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n384), .B1(new_n378), .B2(new_n379), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n408), .A2(new_n377), .A3(new_n383), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n406), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n414), .A2(KEYINPUT75), .A3(new_n402), .A4(new_n404), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n415), .A3(new_n390), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n298), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n355), .B1(new_n399), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n391), .A2(new_n396), .A3(new_n398), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n419), .A2(new_n298), .A3(new_n354), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT9), .B(G234), .ZN(new_n422));
  OAI21_X1  g236(.A(G221), .B1(new_n422), .B2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n368), .A2(new_n223), .A3(new_n372), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n229), .A2(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n371), .B(new_n382), .C1(new_n426), .C2(new_n232), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(new_n197), .B2(new_n199), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n427), .A2(new_n428), .B1(new_n429), .B2(new_n384), .ZN(new_n430));
  INV_X1    g244(.A(new_n217), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n425), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G140), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n338), .A2(G227), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n425), .A2(new_n430), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n217), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n427), .B1(new_n200), .B2(new_n384), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n441), .A2(KEYINPUT12), .A3(new_n217), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT12), .B1(new_n441), .B2(new_n217), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n432), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n438), .A2(new_n440), .B1(new_n444), .B2(new_n435), .ZN(new_n445));
  OAI21_X1  g259(.A(G469), .B1(new_n445), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(G469), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n441), .A2(KEYINPUT12), .A3(new_n217), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n441), .A2(new_n217), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n437), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n436), .B1(new_n440), .B2(new_n432), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n447), .B(new_n298), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n424), .B1(new_n446), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G214), .B1(G237), .B2(G902), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT74), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n421), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n460));
  OAI21_X1  g274(.A(G478), .B1(KEYINPUT85), .B2(KEYINPUT15), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(KEYINPUT85), .B2(KEYINPUT15), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n323), .A2(G143), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n202), .B(new_n467), .C1(new_n230), .C2(new_n189), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT83), .B1(new_n246), .B2(G122), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n470));
  INV_X1    g284(.A(G122), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(G116), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n246), .A2(G122), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n473), .A2(new_n359), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n359), .B1(new_n473), .B2(new_n474), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT13), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n466), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G134), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n466), .B1(new_n194), .B2(G143), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n481), .B2(KEYINPUT13), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n465), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n469), .A2(new_n472), .B1(new_n246), .B2(G122), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(new_n359), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n467), .B1(new_n230), .B2(new_n189), .ZN(new_n486));
  OAI211_X1 g300(.A(G134), .B(new_n479), .C1(new_n486), .C2(new_n478), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n485), .A2(KEYINPUT84), .A3(new_n487), .A4(new_n468), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n359), .B1(new_n473), .B2(KEYINPUT14), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n484), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(G134), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n468), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n422), .A2(new_n349), .A3(G953), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n489), .A2(new_n494), .A3(new_n496), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n464), .B1(new_n500), .B2(new_n298), .ZN(new_n501));
  AOI221_X4 g315(.A(new_n497), .B1(new_n491), .B2(new_n493), .C1(new_n483), .C2(new_n488), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n496), .B1(new_n489), .B2(new_n494), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n464), .B(new_n298), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n463), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n462), .ZN(new_n507));
  INV_X1    g321(.A(G952), .ZN(new_n508));
  AOI211_X1 g322(.A(G953), .B(new_n508), .C1(G234), .C2(G237), .ZN(new_n509));
  AOI211_X1 g323(.A(new_n298), .B(new_n338), .C1(G234), .C2(G237), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT21), .B(G898), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n506), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G113), .B(G122), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(new_n356), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n516), .B(KEYINPUT80), .Z(new_n517));
  INV_X1    g331(.A(KEYINPUT78), .ZN(new_n518));
  INV_X1    g332(.A(G237), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n338), .A3(G214), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n189), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n258), .A2(G143), .A3(G214), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n206), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n206), .B1(new_n521), .B2(new_n522), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n518), .A2(new_n524), .B1(new_n525), .B2(KEYINPUT18), .ZN(new_n526));
  INV_X1    g340(.A(new_n524), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT78), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT77), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n308), .A2(new_n529), .A3(new_n310), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n529), .B1(new_n308), .B2(new_n310), .ZN(new_n531));
  OAI21_X1  g345(.A(G146), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n334), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n526), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n525), .A2(KEYINPUT17), .ZN(new_n535));
  INV_X1    g349(.A(new_n522), .ZN(new_n536));
  AOI21_X1  g350(.A(G143), .B1(new_n258), .B2(G214), .ZN(new_n537));
  OAI21_X1  g351(.A(G131), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n521), .A2(new_n206), .A3(new_n522), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n318), .A2(new_n320), .A3(new_n535), .A4(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n517), .A2(new_n534), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT82), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n542), .B2(new_n534), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(new_n516), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n542), .A2(new_n544), .A3(new_n534), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n543), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G475), .B1(new_n549), .B2(G902), .ZN(new_n550));
  AOI22_X1  g364(.A1(KEYINPUT78), .A2(new_n527), .B1(new_n532), .B2(new_n334), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT19), .B1(new_n530), .B2(new_n531), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT19), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n312), .A2(new_n333), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n187), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n315), .B1(new_n540), .B2(new_n538), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n551), .A2(new_n526), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT79), .B1(new_n557), .B2(new_n516), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n556), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n534), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT79), .ZN(new_n561));
  INV_X1    g375(.A(new_n516), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n543), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(G475), .A2(G902), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT81), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n564), .A2(KEYINPUT20), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT20), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n517), .A2(new_n534), .A3(new_n542), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n561), .B1(new_n560), .B2(new_n562), .ZN(new_n570));
  AOI211_X1 g384(.A(KEYINPUT79), .B(new_n516), .C1(new_n534), .C2(new_n559), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n566), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n550), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n460), .B1(new_n514), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n298), .B1(new_n502), .B2(new_n503), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT86), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n462), .B1(new_n578), .B2(new_n504), .ZN(new_n579));
  INV_X1    g393(.A(new_n507), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT20), .B1(new_n564), .B2(new_n566), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n572), .A2(new_n568), .A3(new_n573), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n547), .A2(new_n545), .A3(new_n516), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n298), .B1(new_n584), .B2(new_n543), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n582), .A2(new_n583), .B1(new_n585), .B2(G475), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n581), .A2(KEYINPUT87), .A3(new_n586), .A4(new_n513), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n459), .B1(new_n576), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n305), .A2(new_n353), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT88), .B(G101), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G3));
  OAI21_X1  g405(.A(G472), .B1(new_n275), .B2(G902), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n455), .A2(new_n353), .ZN(new_n593));
  AND4_X1   g407(.A1(new_n278), .A2(new_n592), .A3(new_n593), .A4(new_n287), .ZN(new_n594));
  INV_X1    g408(.A(new_n417), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n595), .A2(KEYINPUT89), .A3(new_n354), .A4(new_n419), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT89), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n420), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n354), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n399), .B2(new_n417), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G478), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G902), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT90), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT33), .B1(new_n500), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n604), .B(KEYINPUT33), .C1(new_n502), .C2(new_n503), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n603), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n577), .A2(new_n602), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n582), .A2(new_n583), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n608), .A2(new_n609), .B1(new_n610), .B2(new_n550), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n512), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n594), .A2(new_n456), .A3(new_n601), .A4(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT91), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT92), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(new_n594), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n601), .A2(new_n456), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n567), .A2(KEYINPUT93), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n610), .B2(KEYINPUT93), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n550), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n506), .B2(new_n507), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n513), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n619), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT35), .B(G107), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NAND3_X1  g443(.A1(new_n278), .A2(new_n592), .A3(new_n287), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n348), .A2(new_n350), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n341), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n336), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n352), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n631), .A2(new_n588), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT94), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n510), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n509), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n623), .A2(new_n625), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n601), .A2(new_n636), .A3(new_n456), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n305), .A2(new_n455), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  XNOR2_X1  g463(.A(KEYINPUT97), .B(KEYINPUT39), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n644), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n455), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT40), .Z(new_n653));
  XOR2_X1   g467(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n421), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n506), .A2(new_n507), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n575), .ZN(new_n657));
  INV_X1    g471(.A(new_n456), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n657), .A2(new_n658), .A3(new_n636), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n653), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n267), .A2(new_n262), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n298), .B1(new_n295), .B2(new_n263), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n288), .A2(new_n291), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT96), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(KEYINPUT96), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n660), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n189), .ZN(G45));
  INV_X1    g482(.A(KEYINPUT98), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n611), .B2(new_n644), .ZN(new_n670));
  INV_X1    g484(.A(new_n609), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n604), .B1(new_n502), .B2(new_n503), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT33), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n606), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n671), .B1(new_n675), .B2(new_n603), .ZN(new_n676));
  INV_X1    g490(.A(new_n644), .ZN(new_n677));
  NOR4_X1   g491(.A1(new_n676), .A2(new_n586), .A3(KEYINPUT98), .A4(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n670), .A2(new_n678), .A3(new_n646), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n305), .A3(new_n455), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  OR2_X1    g495(.A1(new_n452), .A2(new_n453), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n447), .B1(new_n682), .B2(new_n298), .ZN(new_n683));
  INV_X1    g497(.A(new_n454), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n423), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n620), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n353), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n612), .A2(new_n688), .A3(new_n512), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n305), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT99), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n690), .B(new_n692), .ZN(G15));
  NOR2_X1   g507(.A1(new_n626), .A2(new_n688), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n305), .A2(new_n687), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  INV_X1    g510(.A(new_n636), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n576), .B2(new_n587), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n305), .A2(new_n687), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT100), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT100), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n305), .A2(new_n701), .A3(new_n687), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  OAI22_X1  g518(.A1(new_n283), .A2(new_n284), .B1(new_n296), .B2(new_n263), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n276), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n592), .A2(new_n353), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT101), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n592), .A2(new_n709), .A3(new_n353), .A4(new_n706), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n683), .A2(new_n684), .A3(new_n512), .A4(new_n424), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n581), .A2(new_n586), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n456), .A4(new_n601), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT102), .B1(new_n711), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n717), .B(new_n714), .C1(new_n708), .C2(new_n710), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT103), .B(G122), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G24));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n670), .B2(new_n678), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n592), .A2(new_n636), .A3(new_n706), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n603), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n674), .B2(new_n606), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n575), .B(new_n644), .C1(new_n671), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT98), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n608), .A2(new_n609), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n669), .A3(new_n575), .A4(new_n644), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(KEYINPUT104), .A3(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n723), .A2(new_n725), .A3(new_n687), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n421), .A2(new_n658), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n455), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n305), .A2(new_n353), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n723), .A2(new_n732), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n735), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n729), .A2(KEYINPUT104), .A3(new_n731), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT104), .B1(new_n729), .B2(new_n731), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n291), .A2(KEYINPUT105), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n290), .A2(new_n747), .A3(KEYINPUT32), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n279), .B1(new_n275), .B2(new_n277), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n746), .A2(new_n304), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n737), .A2(new_n735), .A3(new_n738), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n745), .A2(new_n353), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n742), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  INV_X1    g568(.A(new_n645), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n305), .A2(new_n353), .A3(new_n755), .A4(new_n739), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n730), .A2(new_n758), .A3(new_n586), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n676), .B2(new_n575), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n759), .A2(new_n760), .A3(new_n636), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT44), .A3(new_n630), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT44), .B1(new_n761), .B2(new_n630), .ZN(new_n764));
  INV_X1    g578(.A(new_n651), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n451), .A2(new_n448), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n436), .B1(new_n767), .B2(new_n432), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n440), .A2(new_n432), .A3(new_n436), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n438), .A2(new_n440), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n444), .A2(new_n435), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT45), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(G469), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(G469), .A2(G902), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT46), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n684), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n775), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n424), .B(new_n765), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n736), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n763), .A2(new_n764), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n204), .ZN(G39));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n775), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n774), .B2(new_n775), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n785), .A2(new_n786), .A3(new_n684), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n784), .B1(new_n787), .B2(new_n424), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n778), .A2(new_n779), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(KEYINPUT47), .A3(new_n423), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n288), .A2(new_n291), .A3(new_n304), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n688), .A2(new_n729), .A3(new_n731), .A4(new_n736), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  NAND2_X1  g609(.A1(new_n665), .A2(new_n666), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n353), .A2(new_n458), .A3(new_n423), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT106), .ZN(new_n798));
  INV_X1    g612(.A(new_n685), .ZN(new_n799));
  AOI211_X1 g613(.A(new_n575), .B(new_n676), .C1(new_n799), .C2(KEYINPUT49), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(KEYINPUT49), .B2(new_n799), .ZN(new_n801));
  OR4_X1    g615(.A1(new_n796), .A2(new_n655), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n508), .A2(new_n338), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n759), .A2(new_n760), .A3(new_n509), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n711), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n655), .A2(new_n456), .A3(new_n686), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n806), .A2(new_n736), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n788), .B(new_n790), .C1(new_n423), .C2(new_n799), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n737), .A2(new_n686), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n725), .A2(new_n805), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n353), .A3(new_n509), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n796), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n676), .A2(new_n586), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n804), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n508), .B(G953), .C1(new_n806), .C2(new_n687), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n818), .B2(new_n612), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n750), .A2(new_n353), .A3(new_n815), .A4(new_n805), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(KEYINPUT48), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT113), .Z(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(KEYINPUT48), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT114), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n823), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n820), .A2(KEYINPUT111), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n812), .B(KEYINPUT112), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n811), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n810), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n820), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n821), .B(new_n829), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n711), .A2(new_n715), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n717), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n711), .A2(KEYINPUT102), .A3(new_n715), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n457), .B1(new_n418), .B2(new_n420), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n594), .A2(new_n840), .A3(new_n613), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n513), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT107), .B1(new_n581), .B2(new_n575), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT107), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n656), .A2(new_n844), .A3(new_n586), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n842), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n594), .A2(new_n846), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n589), .A2(new_n637), .A3(new_n841), .A4(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n305), .B(new_n687), .C1(new_n689), .C2(new_n694), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n839), .A2(new_n703), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n305), .A2(new_n353), .A3(new_n755), .A4(new_n739), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n723), .A2(new_n592), .A3(new_n706), .A4(new_n732), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n622), .A2(new_n656), .A3(new_n624), .A4(new_n677), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n305), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n737), .A2(new_n738), .A3(new_n697), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n753), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n697), .A2(new_n455), .A3(new_n644), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n620), .A3(new_n657), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n664), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n680), .A2(new_n648), .A3(new_n733), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT108), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n865), .A4(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n697), .B(new_n459), .C1(new_n576), .C2(new_n587), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n871), .A2(new_n631), .B1(new_n594), .B2(new_n846), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n849), .A3(new_n589), .A4(new_n841), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n719), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n703), .A3(new_n753), .A4(new_n857), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n863), .B(KEYINPUT52), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n870), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n869), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n870), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n876), .A2(new_n850), .A3(new_n858), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n700), .A2(new_n702), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n882), .A2(new_n719), .A3(new_n873), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n857), .A2(new_n753), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n865), .A4(new_n868), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n880), .A2(new_n881), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n879), .B(KEYINPUT110), .C1(new_n887), .C2(new_n878), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT110), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n885), .A2(new_n886), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n875), .A2(new_n870), .A3(new_n876), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n889), .B(KEYINPUT54), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n835), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n803), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g709(.A(KEYINPUT115), .B(new_n835), .C1(new_n888), .C2(new_n892), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n802), .B1(new_n895), .B2(new_n896), .ZN(G75));
  AOI21_X1  g711(.A(new_n298), .B1(new_n869), .B2(new_n877), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n898), .A2(KEYINPUT117), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(KEYINPUT117), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n355), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n391), .A2(new_n398), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n396), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n898), .A2(new_n907), .A3(G210), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n907), .B1(new_n898), .B2(G210), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n338), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n906), .A2(new_n912), .A3(new_n914), .ZN(G51));
  NAND2_X1  g729(.A1(new_n869), .A2(new_n877), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n878), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n775), .B(KEYINPUT57), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n682), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n774), .B(KEYINPUT118), .Z(new_n920));
  NAND3_X1  g734(.A1(new_n899), .A2(new_n900), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n913), .B1(new_n919), .B2(new_n921), .ZN(G54));
  AND2_X1   g736(.A1(KEYINPUT58), .A2(G475), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n899), .A2(new_n900), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n564), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n899), .A2(new_n572), .A3(new_n900), .A4(new_n923), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n925), .A2(new_n914), .A3(new_n926), .ZN(G60));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n675), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n914), .B1(new_n917), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n675), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n888), .A2(new_n892), .A3(new_n930), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT119), .Z(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT60), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n869), .B2(new_n877), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n351), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n913), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n940), .A2(new_n634), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT120), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n914), .B(new_n948), .C1(new_n940), .C2(new_n351), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n940), .A2(new_n950), .A3(new_n634), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n947), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n943), .A2(new_n946), .A3(new_n948), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n945), .A2(new_n952), .B1(new_n953), .B2(KEYINPUT61), .ZN(G66));
  INV_X1    g768(.A(new_n511), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n338), .B1(new_n955), .B2(G224), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n850), .B2(new_n338), .ZN(new_n957));
  INV_X1    g771(.A(G898), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n902), .B1(new_n958), .B2(G953), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  AND3_X1   g774(.A1(new_n680), .A2(new_n648), .A3(new_n733), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n764), .A2(new_n781), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n762), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n680), .A2(new_n648), .A3(new_n733), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT122), .B1(new_n782), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n620), .A2(new_n657), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n750), .A2(new_n353), .A3(new_n969), .A4(new_n780), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n794), .A2(new_n756), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n742), .B2(new_n752), .ZN(new_n972));
  AOI21_X1  g786(.A(G953), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n338), .A2(G900), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT123), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n976));
  INV_X1    g790(.A(new_n974), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n794), .A2(new_n756), .A3(new_n970), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n753), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n967), .B2(new_n965), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n976), .B(new_n977), .C1(new_n980), .C2(G953), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n552), .A2(new_n554), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n242), .B(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n975), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n843), .A2(new_n845), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n652), .B(new_n737), .C1(new_n987), .C2(new_n612), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n305), .A3(new_n353), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n963), .A2(new_n794), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n660), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n796), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(KEYINPUT62), .A3(new_n961), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n667), .B2(new_n966), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n990), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n983), .B1(new_n996), .B2(G953), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n338), .B1(G227), .B2(G900), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n985), .A2(new_n986), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n986), .B1(new_n985), .B2(new_n1000), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n973), .A2(new_n974), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n983), .B1(new_n1004), .B2(new_n976), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n1005), .B2(new_n975), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT125), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n975), .A2(new_n981), .A3(new_n1007), .A4(new_n984), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n998), .ZN(new_n1009));
  OAI22_X1  g823(.A1(new_n1001), .A2(new_n1002), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT126), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI221_X1 g826(.A(KEYINPUT126), .B1(new_n1006), .B2(new_n1009), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(G72));
  NAND2_X1  g828(.A1(new_n996), .A2(new_n883), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n661), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT127), .Z(new_n1020));
  NAND2_X1  g834(.A1(new_n301), .A2(new_n264), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n1017), .B(new_n1021), .C1(new_n890), .C2(new_n891), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n980), .A2(new_n883), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n1017), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n281), .A2(new_n282), .A3(new_n263), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n913), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n1020), .A2(new_n1022), .A3(new_n1026), .ZN(G57));
endmodule


