

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707;

  INV_X2 U368 ( .A(G953), .ZN(n384) );
  OR2_X1 U369 ( .A1(n588), .A2(n577), .ZN(n437) );
  AND2_X1 U370 ( .A1(n571), .A2(n672), .ZN(n560) );
  XNOR2_X1 U371 ( .A(n560), .B(n559), .ZN(n705) );
  NOR2_X2 U372 ( .A1(n584), .A2(n615), .ZN(n586) );
  NOR2_X2 U373 ( .A1(n591), .A2(n615), .ZN(n592) );
  NOR2_X2 U374 ( .A1(n596), .A2(n615), .ZN(n598) );
  XNOR2_X2 U375 ( .A(n694), .B(n389), .ZN(n411) );
  XNOR2_X2 U376 ( .A(n450), .B(n388), .ZN(n694) );
  NOR2_X1 U377 ( .A1(n496), .A2(n635), .ZN(n506) );
  AND2_X1 U378 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U379 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U380 ( .A(n349), .B(n348), .ZN(n599) );
  NOR2_X1 U381 ( .A1(n555), .A2(n621), .ZN(n557) );
  XNOR2_X1 U382 ( .A(n380), .B(KEYINPUT66), .ZN(n635) );
  NOR2_X1 U383 ( .A1(G902), .A2(n612), .ZN(n392) );
  XNOR2_X1 U384 ( .A(n390), .B(n411), .ZN(n612) );
  XNOR2_X1 U385 ( .A(n366), .B(n365), .ZN(n454) );
  XNOR2_X1 U386 ( .A(G143), .B(G128), .ZN(n422) );
  XNOR2_X1 U387 ( .A(G119), .B(G116), .ZN(n407) );
  XNOR2_X2 U388 ( .A(n524), .B(n523), .ZN(n680) );
  INV_X1 U389 ( .A(G137), .ZN(n387) );
  INV_X1 U390 ( .A(KEYINPUT8), .ZN(n365) );
  XNOR2_X1 U391 ( .A(G137), .B(G119), .ZN(n362) );
  INV_X1 U392 ( .A(G146), .ZN(n389) );
  XNOR2_X1 U393 ( .A(n359), .B(n383), .ZN(n419) );
  XNOR2_X1 U394 ( .A(n382), .B(n381), .ZN(n359) );
  XNOR2_X1 U395 ( .A(G107), .B(G104), .ZN(n382) );
  NAND2_X2 U396 ( .A1(n356), .A2(n353), .ZN(n600) );
  NAND2_X1 U397 ( .A1(n579), .A2(n354), .ZN(n353) );
  OR2_X2 U398 ( .A1(n617), .A2(n357), .ZN(n356) );
  XNOR2_X1 U399 ( .A(n352), .B(n500), .ZN(n351) );
  XNOR2_X1 U400 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U401 ( .A(n528), .B(KEYINPUT105), .ZN(n529) );
  BUF_X1 U402 ( .A(n600), .Z(n609) );
  NOR2_X1 U403 ( .A1(n384), .A2(G952), .ZN(n615) );
  INV_X1 U404 ( .A(KEYINPUT5), .ZN(n403) );
  XOR2_X1 U405 ( .A(G122), .B(G104), .Z(n444) );
  XNOR2_X1 U406 ( .A(G101), .B(KEYINPUT74), .ZN(n381) );
  NAND2_X1 U407 ( .A1(n577), .A2(n578), .ZN(n355) );
  NAND2_X1 U408 ( .A1(n577), .A2(KEYINPUT2), .ZN(n357) );
  INV_X1 U409 ( .A(KEYINPUT28), .ZN(n528) );
  XNOR2_X1 U410 ( .A(G116), .B(G107), .ZN(n451) );
  XNOR2_X1 U411 ( .A(n557), .B(n556), .ZN(n571) );
  XNOR2_X1 U412 ( .A(n467), .B(KEYINPUT0), .ZN(n512) );
  XNOR2_X1 U413 ( .A(n347), .B(n438), .ZN(n367) );
  XNOR2_X1 U414 ( .A(n419), .B(n358), .ZN(n390) );
  XNOR2_X1 U415 ( .A(n385), .B(n439), .ZN(n358) );
  NAND2_X1 U416 ( .A1(n351), .A2(n350), .ZN(n349) );
  INV_X1 U417 ( .A(n501), .ZN(n350) );
  NOR2_X1 U418 ( .A1(n561), .A2(n534), .ZN(n669) );
  INV_X1 U419 ( .A(n605), .ZN(n606) );
  AND2_X1 U420 ( .A1(n454), .A2(G221), .ZN(n347) );
  XOR2_X1 U421 ( .A(KEYINPUT76), .B(KEYINPUT35), .Z(n348) );
  NAND2_X1 U422 ( .A1(n650), .A2(n508), .ZN(n352) );
  NAND2_X1 U423 ( .A1(n600), .A2(G210), .ZN(n590) );
  NOR2_X1 U424 ( .A1(n680), .A2(n355), .ZN(n354) );
  XNOR2_X2 U425 ( .A(n525), .B(KEYINPUT1), .ZN(n496) );
  XOR2_X1 U426 ( .A(G140), .B(G110), .Z(n360) );
  INV_X1 U427 ( .A(n630), .ZN(n378) );
  XNOR2_X1 U428 ( .A(n404), .B(n403), .ZN(n405) );
  NAND2_X1 U429 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U430 ( .A(n406), .B(n405), .ZN(n410) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n472) );
  INV_X1 U432 ( .A(KEYINPUT39), .ZN(n556) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n601) );
  INV_X1 U434 ( .A(n601), .ZN(n602) );
  XNOR2_X1 U435 ( .A(n558), .B(KEYINPUT106), .ZN(n559) );
  XNOR2_X1 U436 ( .A(G128), .B(KEYINPUT24), .ZN(n361) );
  XNOR2_X1 U437 ( .A(n361), .B(KEYINPUT23), .ZN(n364) );
  XNOR2_X1 U438 ( .A(n360), .B(n362), .ZN(n363) );
  XOR2_X1 U439 ( .A(n364), .B(n363), .Z(n368) );
  NAND2_X1 U440 ( .A1(n384), .A2(G234), .ZN(n366) );
  XNOR2_X1 U441 ( .A(G146), .B(G125), .ZN(n425) );
  XNOR2_X1 U442 ( .A(n425), .B(KEYINPUT10), .ZN(n438) );
  INV_X1 U443 ( .A(G902), .ZN(n459) );
  NAND2_X1 U444 ( .A1(n601), .A2(n459), .ZN(n374) );
  XNOR2_X1 U445 ( .A(KEYINPUT84), .B(KEYINPUT15), .ZN(n369) );
  XNOR2_X1 U446 ( .A(n369), .B(G902), .ZN(n580) );
  NAND2_X1 U447 ( .A1(n580), .A2(G234), .ZN(n370) );
  XNOR2_X1 U448 ( .A(KEYINPUT20), .B(n370), .ZN(n375) );
  NAND2_X1 U449 ( .A1(n375), .A2(G217), .ZN(n372) );
  XOR2_X1 U450 ( .A(KEYINPUT25), .B(KEYINPUT90), .Z(n371) );
  XOR2_X1 U451 ( .A(n372), .B(n371), .Z(n373) );
  INV_X1 U452 ( .A(n472), .ZN(n379) );
  AND2_X1 U453 ( .A1(n375), .A2(G221), .ZN(n377) );
  XNOR2_X1 U454 ( .A(KEYINPUT91), .B(KEYINPUT21), .ZN(n376) );
  XNOR2_X1 U455 ( .A(n377), .B(n376), .ZN(n630) );
  XNOR2_X1 U456 ( .A(KEYINPUT85), .B(G110), .ZN(n383) );
  XOR2_X1 U457 ( .A(G131), .B(G140), .Z(n439) );
  NAND2_X1 U458 ( .A1(G227), .A2(n384), .ZN(n385) );
  XNOR2_X1 U459 ( .A(n422), .B(G134), .ZN(n450) );
  INV_X1 U460 ( .A(KEYINPUT68), .ZN(n386) );
  XNOR2_X1 U461 ( .A(n386), .B(KEYINPUT4), .ZN(n424) );
  XNOR2_X1 U462 ( .A(n424), .B(n387), .ZN(n388) );
  XNOR2_X1 U463 ( .A(KEYINPUT70), .B(G469), .ZN(n391) );
  XNOR2_X2 U464 ( .A(n392), .B(n391), .ZN(n525) );
  NOR2_X1 U465 ( .A1(n635), .A2(n525), .ZN(n511) );
  XNOR2_X1 U466 ( .A(n511), .B(KEYINPUT103), .ZN(n399) );
  XOR2_X1 U467 ( .A(KEYINPUT14), .B(KEYINPUT89), .Z(n394) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n393) );
  XNOR2_X1 U469 ( .A(n394), .B(n393), .ZN(n395) );
  NAND2_X1 U470 ( .A1(G952), .A2(n395), .ZN(n648) );
  NOR2_X1 U471 ( .A1(n648), .A2(G953), .ZN(n465) );
  NAND2_X1 U472 ( .A1(G902), .A2(n395), .ZN(n463) );
  NOR2_X1 U473 ( .A1(G900), .A2(n463), .ZN(n396) );
  NAND2_X1 U474 ( .A1(G953), .A2(n396), .ZN(n397) );
  XNOR2_X1 U475 ( .A(KEYINPUT101), .B(n397), .ZN(n398) );
  NOR2_X1 U476 ( .A1(n465), .A2(n398), .ZN(n477) );
  NOR2_X1 U477 ( .A1(n399), .A2(n477), .ZN(n416) );
  OR2_X1 U478 ( .A1(G237), .A2(G902), .ZN(n432) );
  NAND2_X1 U479 ( .A1(n432), .A2(G214), .ZN(n400) );
  XNOR2_X1 U480 ( .A(n400), .B(KEYINPUT88), .ZN(n482) );
  INV_X1 U481 ( .A(n482), .ZN(n620) );
  XOR2_X1 U482 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n402) );
  NOR2_X1 U483 ( .A1(G953), .A2(G237), .ZN(n440) );
  NAND2_X1 U484 ( .A1(n440), .A2(G210), .ZN(n401) );
  XNOR2_X1 U485 ( .A(n402), .B(n401), .ZN(n406) );
  XNOR2_X1 U486 ( .A(G101), .B(G131), .ZN(n404) );
  XNOR2_X1 U487 ( .A(n407), .B(KEYINPUT3), .ZN(n409) );
  XNOR2_X1 U488 ( .A(G113), .B(KEYINPUT71), .ZN(n408) );
  XNOR2_X1 U489 ( .A(n409), .B(n408), .ZN(n418) );
  XNOR2_X1 U490 ( .A(n410), .B(n418), .ZN(n412) );
  XNOR2_X1 U491 ( .A(n412), .B(n411), .ZN(n593) );
  NAND2_X1 U492 ( .A1(n593), .A2(n459), .ZN(n413) );
  XNOR2_X2 U493 ( .A(n413), .B(G472), .ZN(n633) );
  XNOR2_X1 U494 ( .A(n633), .B(KEYINPUT99), .ZN(n527) );
  NOR2_X1 U495 ( .A1(n620), .A2(n527), .ZN(n414) );
  XNOR2_X1 U496 ( .A(n414), .B(KEYINPUT30), .ZN(n415) );
  NAND2_X1 U497 ( .A1(n416), .A2(n415), .ZN(n555) );
  XNOR2_X1 U498 ( .A(KEYINPUT16), .B(G122), .ZN(n417) );
  XNOR2_X1 U499 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U500 ( .A(n420), .B(n419), .ZN(n687) );
  XNOR2_X1 U501 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n421) );
  XNOR2_X1 U502 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U503 ( .A(n424), .B(n423), .ZN(n430) );
  INV_X1 U504 ( .A(n425), .ZN(n428) );
  NAND2_X1 U505 ( .A1(n384), .A2(G224), .ZN(n426) );
  XNOR2_X1 U506 ( .A(n426), .B(KEYINPUT86), .ZN(n427) );
  XNOR2_X1 U507 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U508 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U509 ( .A(n687), .B(n431), .ZN(n588) );
  INV_X1 U510 ( .A(n580), .ZN(n577) );
  NAND2_X1 U511 ( .A1(n432), .A2(G210), .ZN(n435) );
  INV_X1 U512 ( .A(KEYINPUT78), .ZN(n433) );
  XNOR2_X1 U513 ( .A(n433), .B(KEYINPUT87), .ZN(n434) );
  XNOR2_X1 U514 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X2 U515 ( .A(n437), .B(n436), .ZN(n554) );
  XNOR2_X1 U516 ( .A(n439), .B(n438), .ZN(n693) );
  XOR2_X1 U517 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n442) );
  NAND2_X1 U518 ( .A1(G214), .A2(n440), .ZN(n441) );
  XNOR2_X1 U519 ( .A(n442), .B(n441), .ZN(n446) );
  XNOR2_X1 U520 ( .A(G143), .B(G113), .ZN(n443) );
  XNOR2_X1 U521 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U522 ( .A(n446), .B(n445), .Z(n447) );
  XNOR2_X1 U523 ( .A(n693), .B(n447), .ZN(n581) );
  NAND2_X1 U524 ( .A1(n581), .A2(n459), .ZN(n449) );
  XOR2_X1 U525 ( .A(KEYINPUT13), .B(G475), .Z(n448) );
  XNOR2_X1 U526 ( .A(n449), .B(n448), .ZN(n516) );
  XOR2_X1 U527 ( .A(KEYINPUT9), .B(G122), .Z(n452) );
  XNOR2_X1 U528 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U529 ( .A(n450), .B(n453), .ZN(n458) );
  NAND2_X1 U530 ( .A1(G217), .A2(n454), .ZN(n456) );
  XNOR2_X1 U531 ( .A(KEYINPUT7), .B(KEYINPUT96), .ZN(n455) );
  XNOR2_X1 U532 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U533 ( .A(n458), .B(n457), .ZN(n605) );
  NAND2_X1 U534 ( .A1(n605), .A2(n459), .ZN(n461) );
  INV_X1 U535 ( .A(G478), .ZN(n460) );
  XNOR2_X1 U536 ( .A(n461), .B(n460), .ZN(n515) );
  INV_X1 U537 ( .A(n515), .ZN(n468) );
  NAND2_X1 U538 ( .A1(n516), .A2(n468), .ZN(n501) );
  OR2_X1 U539 ( .A1(n554), .A2(n501), .ZN(n462) );
  NOR2_X1 U540 ( .A1(n555), .A2(n462), .ZN(n540) );
  XOR2_X1 U541 ( .A(G143), .B(n540), .Z(G45) );
  OR2_X2 U542 ( .A1(n554), .A2(n620), .ZN(n545) );
  XNOR2_X2 U543 ( .A(n545), .B(KEYINPUT19), .ZN(n533) );
  INV_X1 U544 ( .A(G898), .ZN(n684) );
  NAND2_X1 U545 ( .A1(G953), .A2(n684), .ZN(n688) );
  NOR2_X1 U546 ( .A1(n463), .A2(n688), .ZN(n464) );
  OR2_X1 U547 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U548 ( .A1(n533), .A2(n466), .ZN(n467) );
  NOR2_X1 U549 ( .A1(n468), .A2(n516), .ZN(n622) );
  NAND2_X1 U550 ( .A1(n622), .A2(n378), .ZN(n469) );
  OR2_X1 U551 ( .A1(n512), .A2(n469), .ZN(n471) );
  XNOR2_X1 U552 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n470) );
  XNOR2_X2 U553 ( .A(n471), .B(n470), .ZN(n493) );
  INV_X1 U554 ( .A(n527), .ZN(n474) );
  INV_X1 U555 ( .A(n496), .ZN(n490) );
  NAND2_X1 U556 ( .A1(n472), .A2(n496), .ZN(n473) );
  NOR2_X1 U557 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U558 ( .A1(n493), .A2(n475), .ZN(n502) );
  XNOR2_X1 U559 ( .A(n502), .B(G110), .ZN(G12) );
  NAND2_X1 U560 ( .A1(n515), .A2(n516), .ZN(n476) );
  XNOR2_X1 U561 ( .A(n476), .B(KEYINPUT97), .ZN(n672) );
  NOR2_X1 U562 ( .A1(n477), .A2(n630), .ZN(n478) );
  XOR2_X1 U563 ( .A(KEYINPUT69), .B(n478), .Z(n479) );
  NAND2_X1 U564 ( .A1(n479), .A2(n472), .ZN(n526) );
  XNOR2_X1 U565 ( .A(n633), .B(KEYINPUT6), .ZN(n486) );
  NOR2_X1 U566 ( .A1(n526), .A2(n486), .ZN(n480) );
  NAND2_X1 U567 ( .A1(n672), .A2(n480), .ZN(n481) );
  XNOR2_X1 U568 ( .A(KEYINPUT102), .B(n481), .ZN(n546) );
  NAND2_X1 U569 ( .A1(n482), .A2(n496), .ZN(n483) );
  NOR2_X1 U570 ( .A1(n546), .A2(n483), .ZN(n484) );
  XOR2_X1 U571 ( .A(n484), .B(KEYINPUT43), .Z(n485) );
  NAND2_X1 U572 ( .A1(n485), .A2(n554), .ZN(n574) );
  XNOR2_X1 U573 ( .A(n574), .B(G140), .ZN(G42) );
  INV_X1 U574 ( .A(n486), .ZN(n497) );
  NAND2_X1 U575 ( .A1(n379), .A2(n496), .ZN(n487) );
  NOR2_X1 U576 ( .A1(n497), .A2(n487), .ZN(n488) );
  NAND2_X1 U577 ( .A1(n493), .A2(n488), .ZN(n489) );
  XOR2_X1 U578 ( .A(KEYINPUT98), .B(n489), .Z(n518) );
  XOR2_X1 U579 ( .A(G101), .B(n518), .Z(G3) );
  XOR2_X1 U580 ( .A(KEYINPUT83), .B(n490), .Z(n548) );
  NOR2_X1 U581 ( .A1(n497), .A2(n379), .ZN(n491) );
  NAND2_X1 U582 ( .A1(n548), .A2(n491), .ZN(n492) );
  XNOR2_X1 U583 ( .A(n492), .B(KEYINPUT77), .ZN(n494) );
  NAND2_X1 U584 ( .A1(n494), .A2(n493), .ZN(n495) );
  XOR2_X1 U585 ( .A(KEYINPUT32), .B(n495), .Z(n503) );
  XOR2_X1 U586 ( .A(n503), .B(G119), .Z(G21) );
  XNOR2_X1 U587 ( .A(n506), .B(KEYINPUT100), .ZN(n498) );
  NAND2_X1 U588 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X2 U589 ( .A(n499), .B(KEYINPUT33), .ZN(n650) );
  INV_X1 U590 ( .A(n512), .ZN(n508) );
  XOR2_X1 U591 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n500) );
  NAND2_X1 U592 ( .A1(n599), .A2(n502), .ZN(n504) );
  XNOR2_X1 U593 ( .A(n505), .B(KEYINPUT44), .ZN(n521) );
  NAND2_X1 U594 ( .A1(n506), .A2(n633), .ZN(n507) );
  XNOR2_X1 U595 ( .A(n507), .B(KEYINPUT95), .ZN(n640) );
  NAND2_X1 U596 ( .A1(n640), .A2(n508), .ZN(n509) );
  XNOR2_X1 U597 ( .A(n509), .B(KEYINPUT31), .ZN(n675) );
  INV_X1 U598 ( .A(n633), .ZN(n510) );
  NAND2_X1 U599 ( .A1(n511), .A2(n510), .ZN(n513) );
  NOR2_X1 U600 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U601 ( .A(n514), .B(KEYINPUT94), .ZN(n661) );
  NOR2_X1 U602 ( .A1(n675), .A2(n661), .ZN(n517) );
  NOR2_X1 U603 ( .A1(n516), .A2(n515), .ZN(n674) );
  NOR2_X1 U604 ( .A1(n674), .A2(n672), .ZN(n541) );
  INV_X1 U605 ( .A(n541), .ZN(n624) );
  XNOR2_X1 U606 ( .A(KEYINPUT81), .B(n624), .ZN(n537) );
  NOR2_X1 U607 ( .A1(n517), .A2(n537), .ZN(n519) );
  NOR2_X1 U608 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U609 ( .A1(n521), .A2(n520), .ZN(n524) );
  XNOR2_X1 U610 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n522) );
  XNOR2_X1 U611 ( .A(n522), .B(KEYINPUT65), .ZN(n523) );
  XOR2_X1 U612 ( .A(n525), .B(KEYINPUT104), .Z(n532) );
  NOR2_X1 U613 ( .A1(n527), .A2(n526), .ZN(n530) );
  NAND2_X1 U614 ( .A1(n532), .A2(n531), .ZN(n561) );
  INV_X1 U615 ( .A(n533), .ZN(n534) );
  INV_X1 U616 ( .A(KEYINPUT67), .ZN(n535) );
  NAND2_X1 U617 ( .A1(n669), .A2(n535), .ZN(n536) );
  XNOR2_X1 U618 ( .A(n536), .B(KEYINPUT47), .ZN(n539) );
  NAND2_X1 U619 ( .A1(n669), .A2(n537), .ZN(n538) );
  AND2_X1 U620 ( .A1(n539), .A2(n538), .ZN(n552) );
  INV_X1 U621 ( .A(n540), .ZN(n543) );
  NAND2_X1 U622 ( .A1(KEYINPUT47), .A2(n541), .ZN(n542) );
  NAND2_X1 U623 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U624 ( .A(n544), .B(KEYINPUT79), .ZN(n550) );
  NOR2_X1 U625 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U626 ( .A(n547), .B(KEYINPUT36), .ZN(n549) );
  NAND2_X1 U627 ( .A1(n549), .A2(n548), .ZN(n678) );
  NAND2_X1 U628 ( .A1(n550), .A2(n678), .ZN(n551) );
  NOR2_X1 U629 ( .A1(n552), .A2(n551), .ZN(n569) );
  INV_X1 U630 ( .A(KEYINPUT38), .ZN(n553) );
  XNOR2_X1 U631 ( .A(n554), .B(n553), .ZN(n621) );
  XNOR2_X1 U632 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n558) );
  INV_X1 U633 ( .A(n561), .ZN(n564) );
  NOR2_X1 U634 ( .A1(n621), .A2(n620), .ZN(n562) );
  XNOR2_X1 U635 ( .A(n562), .B(KEYINPUT108), .ZN(n625) );
  NAND2_X1 U636 ( .A1(n625), .A2(n622), .ZN(n563) );
  XNOR2_X1 U637 ( .A(n563), .B(KEYINPUT41), .ZN(n651) );
  NAND2_X1 U638 ( .A1(n564), .A2(n651), .ZN(n565) );
  XNOR2_X1 U639 ( .A(n565), .B(KEYINPUT42), .ZN(n707) );
  NAND2_X1 U640 ( .A1(n705), .A2(n707), .ZN(n567) );
  XOR2_X1 U641 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n566) );
  XNOR2_X1 U642 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U643 ( .A(n570), .B(KEYINPUT48), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n571), .A2(n674), .ZN(n573) );
  INV_X1 U645 ( .A(KEYINPUT109), .ZN(n572) );
  XNOR2_X1 U646 ( .A(n573), .B(n572), .ZN(n706) );
  AND2_X1 U647 ( .A1(n706), .A2(n574), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n698) );
  NOR2_X1 U649 ( .A1(n680), .A2(n698), .ZN(n617) );
  INV_X1 U650 ( .A(KEYINPUT2), .ZN(n578) );
  XNOR2_X1 U651 ( .A(n698), .B(KEYINPUT75), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n600), .A2(G475), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n581), .B(KEYINPUT59), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U655 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n585) );
  XNOR2_X1 U656 ( .A(n586), .B(n585), .ZN(G60) );
  XOR2_X1 U657 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n587) );
  XNOR2_X1 U658 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U659 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n592), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U661 ( .A1(n600), .A2(G472), .ZN(n595) );
  XOR2_X1 U662 ( .A(n593), .B(KEYINPUT62), .Z(n594) );
  XNOR2_X1 U663 ( .A(n595), .B(n594), .ZN(n596) );
  XOR2_X1 U664 ( .A(KEYINPUT110), .B(KEYINPUT63), .Z(n597) );
  XNOR2_X1 U665 ( .A(n598), .B(n597), .ZN(G57) );
  XNOR2_X1 U666 ( .A(n599), .B(G122), .ZN(G24) );
  NAND2_X1 U667 ( .A1(n609), .A2(G217), .ZN(n603) );
  XNOR2_X1 U668 ( .A(n603), .B(n602), .ZN(n604) );
  NOR2_X1 U669 ( .A1(n604), .A2(n615), .ZN(G66) );
  NAND2_X1 U670 ( .A1(n609), .A2(G478), .ZN(n607) );
  XNOR2_X1 U671 ( .A(n607), .B(n606), .ZN(n608) );
  NOR2_X1 U672 ( .A1(n608), .A2(n615), .ZN(G63) );
  NAND2_X1 U673 ( .A1(n609), .A2(G469), .ZN(n614) );
  XNOR2_X1 U674 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n610) );
  XNOR2_X1 U675 ( .A(n610), .B(KEYINPUT58), .ZN(n611) );
  XNOR2_X1 U676 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U677 ( .A(n614), .B(n613), .ZN(n616) );
  NOR2_X1 U678 ( .A1(n616), .A2(n615), .ZN(G54) );
  INV_X1 U679 ( .A(n617), .ZN(n618) );
  NAND2_X1 U680 ( .A1(n618), .A2(KEYINPUT80), .ZN(n619) );
  XNOR2_X1 U681 ( .A(n619), .B(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U682 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U683 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U684 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U685 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U686 ( .A1(n650), .A2(n628), .ZN(n629) );
  XNOR2_X1 U687 ( .A(n629), .B(KEYINPUT118), .ZN(n644) );
  NAND2_X1 U688 ( .A1(n630), .A2(n472), .ZN(n631) );
  XNOR2_X1 U689 ( .A(KEYINPUT49), .B(n631), .ZN(n632) );
  NOR2_X1 U690 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U691 ( .A(KEYINPUT117), .B(n634), .ZN(n638) );
  NAND2_X1 U692 ( .A1(n635), .A2(n496), .ZN(n636) );
  XOR2_X1 U693 ( .A(KEYINPUT50), .B(n636), .Z(n637) );
  NOR2_X1 U694 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U695 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U696 ( .A(KEYINPUT51), .B(n641), .ZN(n642) );
  NAND2_X1 U697 ( .A1(n642), .A2(n651), .ZN(n643) );
  NAND2_X1 U698 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U699 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n645) );
  XNOR2_X1 U700 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X1 U701 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U702 ( .A(n649), .B(KEYINPUT120), .ZN(n654) );
  NAND2_X1 U703 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U704 ( .A1(n652), .A2(n384), .ZN(n653) );
  NOR2_X1 U705 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U706 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U707 ( .A(KEYINPUT53), .B(n657), .Z(G75) );
  NAND2_X1 U708 ( .A1(n661), .A2(n672), .ZN(n658) );
  XNOR2_X1 U709 ( .A(n658), .B(G104), .ZN(G6) );
  XOR2_X1 U710 ( .A(KEYINPUT113), .B(KEYINPUT27), .Z(n660) );
  XNOR2_X1 U711 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n659) );
  XNOR2_X1 U712 ( .A(n660), .B(n659), .ZN(n665) );
  XNOR2_X1 U713 ( .A(G107), .B(KEYINPUT26), .ZN(n663) );
  NAND2_X1 U714 ( .A1(n674), .A2(n661), .ZN(n662) );
  XNOR2_X1 U715 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U716 ( .A(n665), .B(n664), .ZN(G9) );
  XOR2_X1 U717 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n667) );
  NAND2_X1 U718 ( .A1(n669), .A2(n674), .ZN(n666) );
  XNOR2_X1 U719 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U720 ( .A(G128), .B(n668), .ZN(G30) );
  XOR2_X1 U721 ( .A(G146), .B(KEYINPUT115), .Z(n671) );
  NAND2_X1 U722 ( .A1(n669), .A2(n672), .ZN(n670) );
  XNOR2_X1 U723 ( .A(n671), .B(n670), .ZN(G48) );
  NAND2_X1 U724 ( .A1(n675), .A2(n672), .ZN(n673) );
  XNOR2_X1 U725 ( .A(n673), .B(G113), .ZN(G15) );
  NAND2_X1 U726 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U727 ( .A(n676), .B(G116), .ZN(G18) );
  XOR2_X1 U728 ( .A(KEYINPUT116), .B(KEYINPUT37), .Z(n677) );
  XNOR2_X1 U729 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U730 ( .A(G125), .B(n679), .ZN(G27) );
  NOR2_X1 U731 ( .A1(n680), .A2(G953), .ZN(n686) );
  NAND2_X1 U732 ( .A1(G224), .A2(G953), .ZN(n681) );
  XNOR2_X1 U733 ( .A(n681), .B(KEYINPUT123), .ZN(n682) );
  XNOR2_X1 U734 ( .A(n682), .B(KEYINPUT61), .ZN(n683) );
  NOR2_X1 U735 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U736 ( .A1(n686), .A2(n685), .ZN(n691) );
  INV_X1 U737 ( .A(n687), .ZN(n689) );
  NAND2_X1 U738 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U739 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U740 ( .A(KEYINPUT124), .B(n692), .ZN(G69) );
  XOR2_X1 U741 ( .A(n694), .B(n693), .Z(n699) );
  XOR2_X1 U742 ( .A(G227), .B(n699), .Z(n695) );
  NAND2_X1 U743 ( .A1(n695), .A2(G900), .ZN(n696) );
  NAND2_X1 U744 ( .A1(G953), .A2(n696), .ZN(n697) );
  XOR2_X1 U745 ( .A(KEYINPUT126), .B(n697), .Z(n703) );
  XNOR2_X1 U746 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U747 ( .A1(G953), .A2(n700), .ZN(n701) );
  XOR2_X1 U748 ( .A(KEYINPUT125), .B(n701), .Z(n702) );
  NOR2_X1 U749 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U750 ( .A(KEYINPUT127), .B(n704), .ZN(G72) );
  XNOR2_X1 U751 ( .A(n705), .B(G131), .ZN(G33) );
  XNOR2_X1 U752 ( .A(G134), .B(n706), .ZN(G36) );
  XNOR2_X1 U753 ( .A(G137), .B(n707), .ZN(G39) );
endmodule

