//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G116), .A2(G270), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G87), .A2(G250), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G50), .B2(G226), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G107), .A2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n218), .B(new_n219), .C1(new_n202), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n203), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n210), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT64), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n225), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n208), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n202), .A2(new_n203), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n213), .B(new_n229), .C1(new_n231), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AOI21_X1  g0050(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n220), .A2(G1698), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n253), .B(new_n254), .C1(G226), .C2(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n252), .A2(G238), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  XOR2_X1   g0062(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR4_X1   g0065(.A1(new_n257), .A2(new_n259), .A3(new_n261), .A4(new_n263), .ZN(new_n266));
  OAI21_X1  g0066(.A(G200), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT69), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n230), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G77), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G50), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(new_n208), .B2(G68), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n271), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  XOR2_X1   g0080(.A(new_n280), .B(KEYINPUT11), .Z(new_n281));
  AOI21_X1  g0081(.A(new_n271), .B1(new_n207), .B2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n203), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n203), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT12), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n281), .A2(new_n284), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT70), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT13), .ZN(new_n292));
  OR3_X1    g0092(.A1(new_n262), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n291), .B1(new_n262), .B2(new_n292), .ZN(new_n294));
  INV_X1    g0094(.A(new_n266), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n293), .A2(new_n294), .A3(G190), .A4(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n296), .A2(new_n297), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n269), .B(new_n290), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(G169), .B1(new_n265), .B2(new_n266), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(KEYINPUT72), .B2(KEYINPUT14), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n293), .A2(new_n294), .A3(G179), .A4(new_n295), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n305));
  OAI211_X1 g0105(.A(G169), .B(new_n305), .C1(new_n265), .C2(new_n266), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n290), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT73), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n252), .A2(new_n258), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n312), .A2(G244), .ZN(new_n313));
  INV_X1    g0113(.A(G1698), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n253), .A2(G232), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n253), .A2(G238), .A3(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G107), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(new_n253), .ZN(new_n318));
  AOI211_X1 g0118(.A(new_n261), .B(new_n313), .C1(new_n318), .C2(new_n251), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(KEYINPUT8), .A2(G58), .ZN(new_n322));
  NAND2_X1  g0122(.A1(KEYINPUT8), .A2(G58), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n277), .B1(G20), .B2(G77), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n274), .B2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n271), .B1(new_n275), .B2(new_n286), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n275), .B2(new_n283), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n321), .B(new_n329), .C1(G169), .C2(new_n319), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n312), .A2(G226), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G222), .A2(G1698), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n314), .A2(G223), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n253), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(new_n251), .C1(G77), .C2(new_n253), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n332), .B(new_n336), .C1(new_n260), .C2(new_n258), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G200), .ZN(new_n338));
  INV_X1    g0138(.A(G190), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR3_X1   g0141(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT66), .B1(new_n342), .B2(new_n208), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT66), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n204), .A2(new_n344), .A3(G20), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n273), .A2(new_n322), .A3(new_n323), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n277), .A2(G150), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n343), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n271), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n286), .A2(new_n201), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n282), .A2(G50), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(KEYINPUT67), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT67), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n348), .A2(new_n271), .B1(new_n201), .B2(new_n286), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(new_n351), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT9), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n352), .A2(KEYINPUT67), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(new_n354), .A3(new_n351), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT9), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n338), .B(new_n341), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT10), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n357), .B1(new_n353), .B2(new_n356), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n359), .A2(KEYINPUT9), .A3(new_n360), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n340), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT10), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n338), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n331), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n311), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n271), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT3), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G33), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT7), .B1(new_n375), .B2(new_n208), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n377), .B(G20), .C1(new_n372), .C2(new_n374), .ZN(new_n378));
  OAI21_X1  g0178(.A(G68), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(KEYINPUT75), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(KEYINPUT75), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n232), .A3(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(G20), .B1(G159), .B2(new_n277), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n371), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n372), .A2(new_n374), .A3(KEYINPUT74), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT74), .B1(new_n372), .B2(new_n374), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n208), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n378), .B1(new_n390), .B2(new_n377), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT16), .B(new_n384), .C1(new_n391), .C2(new_n203), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n207), .A2(G20), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n324), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n286), .A2(new_n271), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n324), .A2(KEYINPUT76), .A3(new_n394), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n324), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n286), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n393), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G169), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n253), .B1(G223), .B2(G1698), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n314), .A2(G226), .ZN(new_n408));
  INV_X1    g0208(.A(G87), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n407), .A2(new_n408), .B1(new_n272), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n251), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n261), .B1(new_n312), .B2(G232), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n411), .A2(new_n412), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n320), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n405), .A2(new_n416), .A3(KEYINPUT18), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n411), .A2(new_n412), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n413), .B1(G179), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n403), .B1(new_n387), .B2(new_n392), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n415), .A2(G200), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n393), .A2(new_n404), .A3(new_n424), .ZN(new_n425));
  OR2_X1    g0225(.A1(KEYINPUT77), .A2(G190), .ZN(new_n426));
  NAND2_X1  g0226(.A1(KEYINPUT77), .A2(G190), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n415), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n425), .A2(KEYINPUT78), .A3(KEYINPUT17), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n421), .A2(new_n429), .A3(new_n424), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n423), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n337), .A2(G179), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n337), .A2(new_n406), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n352), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT73), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n300), .A2(new_n309), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n319), .A2(G190), .ZN(new_n443));
  INV_X1    g0243(.A(new_n329), .ZN(new_n444));
  INV_X1    g0244(.A(G200), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n443), .B(new_n444), .C1(new_n445), .C2(new_n319), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n370), .A2(KEYINPUT79), .A3(new_n440), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT79), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n311), .A2(new_n369), .A3(new_n442), .A4(new_n446), .ZN(new_n450));
  INV_X1    g0250(.A(new_n440), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n372), .A2(new_n374), .A3(new_n208), .A4(G87), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT22), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n253), .A2(new_n456), .A3(new_n208), .A4(G87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n273), .A2(G116), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n208), .A2(G107), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n460), .B(KEYINPUT23), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT85), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT85), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n458), .A2(new_n464), .A3(new_n459), .A4(new_n461), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(KEYINPUT24), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(KEYINPUT85), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n271), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n207), .A2(G33), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n285), .A2(new_n470), .A3(new_n230), .A4(new_n270), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G107), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n285), .A2(G107), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT25), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n469), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G45), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G1), .ZN(new_n478));
  INV_X1    g0278(.A(G41), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT5), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G41), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n252), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G264), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n483), .A2(new_n260), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n253), .A2(G250), .A3(new_n314), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n253), .A2(G257), .A3(G1698), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G294), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n485), .B(new_n486), .C1(new_n490), .C2(new_n252), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G179), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n406), .B2(new_n491), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n476), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT86), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT86), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n476), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n491), .A2(G200), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n476), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n339), .B2(new_n491), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n286), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n472), .A2(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  INV_X1    g0306(.A(G97), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n208), .C1(G33), .C2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n508), .B(new_n271), .C1(new_n208), .C2(G116), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT20), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n509), .A2(new_n510), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n504), .B(new_n505), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n253), .A2(G264), .A3(G1698), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n253), .A2(G257), .A3(new_n314), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n375), .A2(G303), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n251), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n484), .A2(G270), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n486), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n513), .A2(new_n520), .A3(G169), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(G200), .ZN(new_n524));
  INV_X1    g0324(.A(new_n513), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n525), .C1(new_n428), .C2(new_n520), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n513), .A2(new_n520), .A3(KEYINPUT21), .A4(G169), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n520), .A2(new_n320), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n513), .ZN(new_n529));
  AND4_X1   g0329(.A1(new_n523), .A2(new_n526), .A3(new_n527), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n253), .A2(new_n208), .A3(G68), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n274), .B2(new_n507), .ZN(new_n533));
  AND4_X1   g0333(.A1(KEYINPUT82), .A2(new_n409), .A3(new_n507), .A4(new_n317), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G97), .A2(G107), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT82), .B1(new_n535), .B2(new_n409), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n256), .A2(new_n532), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G20), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n531), .B(new_n533), .C1(new_n537), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n271), .ZN(new_n541));
  INV_X1    g0341(.A(new_n326), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n472), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n326), .A2(new_n286), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n222), .A2(new_n314), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n314), .A2(G244), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n253), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n251), .A2(new_n478), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n550), .A2(new_n251), .B1(new_n551), .B2(G250), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n478), .A2(G274), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n552), .A2(new_n320), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(G169), .B1(new_n552), .B2(new_n553), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n545), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n553), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n339), .ZN(new_n558));
  OR3_X1    g0358(.A1(new_n471), .A2(KEYINPUT83), .A3(new_n409), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT83), .B1(new_n471), .B2(new_n409), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n541), .A2(new_n561), .A3(new_n544), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n445), .B1(new_n552), .B2(new_n553), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n558), .B1(new_n564), .B2(KEYINPUT84), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT84), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n562), .B2(new_n563), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n556), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n506), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n253), .A2(G244), .A3(new_n314), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n253), .A2(KEYINPUT4), .A3(G244), .A4(new_n314), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT81), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT81), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n253), .A2(new_n576), .A3(G250), .A4(G1698), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n572), .A2(new_n573), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n251), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n484), .A2(G257), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n486), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n578), .A2(new_n251), .B1(G257), .B2(new_n484), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(G190), .A3(new_n486), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n285), .A2(G97), .ZN(new_n585));
  OAI21_X1  g0385(.A(G107), .B1(new_n376), .B2(new_n378), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n317), .A2(KEYINPUT6), .A3(G97), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n507), .A2(new_n317), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(new_n535), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n587), .B1(new_n589), .B2(KEYINPUT6), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G20), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n277), .A2(G77), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n585), .B1(new_n593), .B2(new_n271), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n472), .A2(G97), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n594), .A2(KEYINPUT80), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT80), .B1(new_n594), .B2(new_n595), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n582), .B(new_n584), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n595), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n583), .A2(G179), .A3(new_n486), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n406), .B1(new_n583), .B2(new_n486), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND4_X1   g0403(.A1(new_n530), .A2(new_n568), .A3(new_n598), .A4(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n453), .A2(new_n502), .A3(new_n604), .ZN(G372));
  NAND2_X1  g0405(.A1(new_n598), .A2(new_n603), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT87), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n562), .B1(new_n608), .B2(new_n563), .ZN(new_n609));
  OAI221_X1 g0409(.A(new_n609), .B1(new_n608), .B2(new_n563), .C1(new_n339), .C2(new_n557), .ZN(new_n610));
  INV_X1    g0410(.A(new_n556), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n523), .A2(new_n527), .A3(new_n529), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n494), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n607), .A2(new_n501), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT88), .B1(new_n601), .B2(new_n602), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n596), .A2(new_n597), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n581), .A2(G169), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(new_n600), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n612), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n603), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n568), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n556), .B1(new_n625), .B2(KEYINPUT26), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n615), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n453), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n300), .A2(new_n331), .B1(new_n308), .B2(new_n307), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n430), .A2(new_n434), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n423), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT89), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n362), .A2(KEYINPUT10), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n367), .B1(new_n366), .B2(new_n338), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n363), .A2(new_n368), .A3(KEYINPUT89), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n439), .B1(new_n631), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n628), .A2(new_n638), .ZN(G369));
  INV_X1    g0439(.A(G13), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G20), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n207), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n476), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n502), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n476), .A2(new_n493), .A3(new_n647), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n513), .A2(new_n647), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT90), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n613), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n530), .B2(new_n653), .ZN(new_n655));
  INV_X1    g0455(.A(G330), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n613), .A2(new_n647), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n498), .A2(new_n501), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n647), .B(KEYINPUT91), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n494), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n658), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n211), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G1), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n537), .A2(new_n503), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n668), .A2(new_n669), .B1(new_n233), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT92), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT28), .ZN(new_n672));
  INV_X1    g0472(.A(new_n661), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n627), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT95), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n498), .A2(new_n613), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(new_n501), .A3(new_n607), .A4(new_n610), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT96), .B1(new_n625), .B2(new_n622), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n621), .A2(new_n612), .A3(KEYINPUT26), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n621), .A2(new_n612), .A3(KEYINPUT96), .A4(KEYINPUT26), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n679), .A2(new_n611), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n647), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(KEYINPUT29), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT95), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n674), .A2(new_n687), .A3(new_n675), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n677), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n604), .A2(new_n498), .A3(new_n501), .A4(new_n673), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT94), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n491), .A2(new_n557), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n528), .A3(new_n583), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n692), .A2(new_n528), .A3(new_n583), .A4(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n581), .A2(new_n491), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n520), .A2(new_n557), .A3(new_n320), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT93), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n520), .A2(new_n557), .A3(KEYINPUT93), .A4(new_n320), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n698), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n691), .B1(new_n697), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n581), .A2(new_n491), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(KEYINPUT94), .A3(new_n695), .A4(new_n696), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n704), .A2(new_n708), .A3(new_n647), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT31), .B(new_n661), .C1(new_n697), .C2(new_n703), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n690), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n689), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n672), .B1(new_n716), .B2(G1), .ZN(G364));
  INV_X1    g0517(.A(new_n657), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n668), .B1(G45), .B2(new_n641), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n655), .A2(new_n656), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT97), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n208), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT98), .Z(new_n726));
  NAND2_X1  g0526(.A1(new_n655), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n388), .A2(new_n389), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n665), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n234), .A2(new_n477), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n729), .B(new_n730), .C1(new_n477), .C2(new_n249), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n211), .A2(G355), .A3(new_n253), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n731), .B(new_n732), .C1(G116), .C2(new_n211), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n230), .B1(G20), .B2(new_n406), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n208), .A2(new_n320), .A3(G200), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n428), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G20), .A3(new_n339), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G159), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n739), .A2(G58), .B1(new_n743), .B2(KEYINPUT32), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n208), .A2(new_n320), .A3(new_n445), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n428), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n744), .B1(KEYINPUT32), .B2(new_n743), .C1(new_n201), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n746), .A2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n738), .A2(G190), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G68), .A2(new_n750), .B1(new_n751), .B2(G77), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n740), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G97), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n445), .A2(G179), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G20), .A3(G190), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n752), .B(new_n755), .C1(new_n409), .C2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n756), .A2(G20), .A3(new_n339), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n317), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n749), .A2(new_n758), .A3(new_n375), .A4(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n754), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  INV_X1    g0563(.A(new_n750), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT33), .B(G317), .Z(new_n765));
  OAI221_X1 g0565(.A(new_n375), .B1(new_n762), .B2(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  INV_X1    g0567(.A(G329), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n759), .A2(new_n767), .B1(new_n768), .B2(new_n741), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(G326), .B2(new_n747), .ZN(new_n770));
  INV_X1    g0570(.A(G303), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(new_n757), .ZN(new_n772));
  INV_X1    g0572(.A(new_n751), .ZN(new_n773));
  INV_X1    g0573(.A(G311), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n739), .A2(G322), .ZN(new_n776));
  NOR4_X1   g0576(.A1(new_n766), .A2(new_n772), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n734), .B1(new_n761), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n727), .A2(new_n719), .A3(new_n736), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT99), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n723), .A2(new_n780), .ZN(G396));
  NAND2_X1  g0581(.A1(new_n329), .A2(new_n647), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n331), .B1(new_n446), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n330), .A2(new_n647), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n724), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G150), .A2(new_n750), .B1(new_n751), .B2(G159), .ZN(new_n788));
  INV_X1    g0588(.A(new_n739), .ZN(new_n789));
  INV_X1    g0589(.A(G143), .ZN(new_n790));
  INV_X1    g0590(.A(G137), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n788), .B1(new_n789), .B2(new_n790), .C1(new_n791), .C2(new_n748), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT34), .Z(new_n793));
  INV_X1    g0593(.A(new_n728), .ZN(new_n794));
  INV_X1    g0594(.A(new_n757), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(G50), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G132), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n759), .A2(new_n203), .B1(new_n797), .B2(new_n741), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n796), .B(new_n799), .C1(new_n202), .C2(new_n762), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT101), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n793), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G283), .A2(new_n750), .B1(new_n751), .B2(G116), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(KEYINPUT100), .B1(G303), .B2(new_n747), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n755), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n759), .A2(new_n409), .B1(new_n774), .B2(new_n741), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n807), .B(new_n375), .C1(new_n317), .C2(new_n757), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n789), .A2(new_n763), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n805), .A2(new_n808), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n734), .B1(new_n802), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n734), .A2(new_n724), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n275), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n787), .A2(new_n719), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n674), .B(new_n786), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(new_n714), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n815), .B1(new_n817), .B2(new_n719), .ZN(G384));
  NAND4_X1  g0618(.A1(new_n704), .A2(new_n708), .A3(KEYINPUT31), .A4(new_n647), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n690), .A2(new_n711), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n290), .A2(new_n685), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n310), .A2(new_n821), .B1(new_n309), .B2(new_n685), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n820), .A2(new_n785), .A3(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n645), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n384), .B1(new_n391), .B2(new_n203), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n371), .B1(new_n825), .B2(new_n386), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n392), .B1(new_n826), .B2(KEYINPUT103), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT103), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n828), .B(new_n371), .C1(new_n825), .C2(new_n386), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n404), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n435), .A2(new_n824), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT37), .ZN(new_n832));
  INV_X1    g0632(.A(new_n432), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n830), .B2(new_n824), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n830), .A2(new_n416), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n405), .B1(new_n416), .B2(new_n824), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n837), .A2(new_n832), .A3(new_n432), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(KEYINPUT38), .B(new_n831), .C1(new_n836), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n421), .A2(new_n645), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n435), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n421), .B1(new_n420), .B2(new_n645), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT37), .B1(new_n833), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n838), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n823), .A2(KEYINPUT40), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n820), .A2(new_n785), .A3(new_n822), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n830), .A2(new_n824), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(new_n835), .A3(new_n432), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n839), .B1(new_n853), .B2(KEYINPUT37), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n435), .A2(new_n824), .A3(new_n830), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n847), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n851), .B1(new_n840), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n858));
  OAI211_X1 g0658(.A(new_n850), .B(G330), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n453), .A2(G330), .A3(new_n820), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n856), .A2(new_n840), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n823), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n858), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n865), .A2(new_n453), .A3(new_n820), .A4(new_n850), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n453), .A2(new_n686), .A3(new_n688), .A4(new_n677), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(new_n638), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n867), .B(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n840), .A2(new_n848), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT104), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n856), .B2(new_n840), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI211_X1 g0675(.A(KEYINPUT104), .B(new_n871), .C1(new_n856), .C2(new_n840), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT105), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n309), .A2(new_n647), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT104), .ZN(new_n879));
  INV_X1    g0679(.A(new_n392), .ZN(new_n880));
  INV_X1    g0680(.A(new_n384), .ZN(new_n881));
  INV_X1    g0681(.A(new_n378), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT74), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n375), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n253), .A2(KEYINPUT74), .ZN(new_n885));
  AOI21_X1  g0685(.A(G20), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n882), .B1(new_n886), .B2(KEYINPUT7), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n881), .B1(new_n887), .B2(G68), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n271), .B1(new_n888), .B2(KEYINPUT16), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n880), .B1(new_n889), .B2(new_n828), .ZN(new_n890));
  INV_X1    g0690(.A(new_n829), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n403), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n432), .B1(new_n892), .B2(new_n645), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n420), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n838), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n896), .B2(new_n831), .ZN(new_n897));
  INV_X1    g0697(.A(new_n840), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n879), .B(KEYINPUT39), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n899), .B(new_n900), .C1(new_n874), .C2(new_n873), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n877), .A2(new_n878), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n423), .A2(new_n824), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n784), .B(KEYINPUT102), .Z(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n674), .B2(new_n786), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n905), .A2(new_n822), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n903), .B1(new_n906), .B2(new_n862), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n870), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n207), .B2(new_n641), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n503), .B1(new_n590), .B2(KEYINPUT35), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n231), .C1(KEYINPUT35), .C2(new_n590), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n234), .A2(G77), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n381), .A2(new_n382), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n914), .A2(new_n915), .B1(G50), .B2(new_n203), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(G1), .A3(new_n640), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n910), .A2(new_n913), .A3(new_n917), .ZN(G367));
  NAND4_X1  g0718(.A1(new_n616), .A2(new_n617), .A3(new_n620), .A4(new_n661), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n596), .A2(new_n673), .A3(new_n597), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n919), .B1(new_n606), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT108), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n922), .A2(new_n502), .A3(new_n648), .A4(new_n659), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT42), .Z(new_n924));
  INV_X1    g0724(.A(new_n922), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n603), .B1(new_n925), .B2(new_n498), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n673), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n562), .A2(new_n647), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n612), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT107), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n556), .A2(new_n562), .A3(new_n647), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(KEYINPUT107), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n924), .A2(new_n927), .B1(KEYINPUT43), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n658), .A2(new_n925), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n937), .B(new_n938), .Z(new_n939));
  INV_X1    g0739(.A(KEYINPUT45), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n925), .B2(new_n662), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n663), .A2(KEYINPUT45), .A3(new_n922), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n925), .A2(KEYINPUT44), .A3(new_n662), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT44), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n663), .B2(new_n922), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT109), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(new_n949), .A3(new_n658), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n658), .A2(new_n949), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n651), .A2(KEYINPUT109), .A3(new_n657), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n943), .A2(new_n947), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n660), .B1(new_n651), .B2(new_n659), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n657), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n718), .B(new_n660), .C1(new_n651), .C2(new_n659), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(new_n714), .A3(new_n689), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n716), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n666), .B(KEYINPUT41), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n207), .B1(new_n641), .B2(G45), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n939), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(G150), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n748), .A2(new_n790), .B1(new_n789), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G68), .B2(new_n754), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n742), .A2(G137), .ZN(new_n971));
  INV_X1    g0771(.A(new_n759), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n750), .A2(G159), .B1(G77), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n757), .A2(new_n202), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n375), .B(new_n974), .C1(G50), .C2(new_n751), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n970), .A2(new_n971), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n773), .A2(new_n767), .B1(new_n762), .B2(new_n317), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n742), .A2(G317), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n794), .B(new_n978), .C1(new_n507), .C2(new_n759), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT111), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n977), .B(new_n980), .C1(G294), .C2(new_n750), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT110), .B1(new_n795), .B2(G116), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT46), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(new_n774), .C2(new_n748), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n789), .A2(new_n771), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n976), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT112), .Z(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n734), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n931), .A2(new_n726), .A3(new_n932), .A4(new_n933), .ZN(new_n990));
  INV_X1    g0790(.A(new_n729), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n735), .B1(new_n211), .B2(new_n326), .C1(new_n991), .C2(new_n242), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n989), .A2(new_n719), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n967), .A2(new_n993), .ZN(G387));
  INV_X1    g0794(.A(KEYINPUT114), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n960), .B2(new_n667), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n959), .A2(KEYINPUT114), .A3(new_n666), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(new_n716), .C2(new_n958), .ZN(new_n998));
  INV_X1    g0798(.A(new_n965), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n958), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n742), .A2(G326), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G311), .A2(new_n750), .B1(new_n739), .B2(G317), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT113), .B(G322), .Z(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n771), .B2(new_n773), .C1(new_n748), .C2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n754), .A2(G283), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n795), .A2(G294), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1001), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1008), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n794), .B1(new_n1011), .B2(KEYINPUT49), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G116), .C2(new_n972), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n751), .A2(G68), .B1(G97), .B2(new_n972), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n275), .B2(new_n757), .C1(new_n401), .C2(new_n764), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n728), .B1(new_n968), .B2(new_n741), .C1(new_n789), .C2(new_n201), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n762), .A2(new_n326), .ZN(new_n1017));
  INV_X1    g0817(.A(G159), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n748), .A2(new_n1018), .ZN(new_n1019));
  NOR4_X1   g0819(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n734), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n649), .A2(new_n650), .A3(new_n726), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n324), .A2(new_n201), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n203), .A2(new_n275), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1024), .A2(G45), .A3(new_n1025), .A4(new_n669), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n729), .B1(new_n239), .B2(new_n477), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n669), .A2(new_n211), .A3(new_n253), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n211), .A2(G107), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n735), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1021), .A2(new_n719), .A3(new_n1022), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n998), .A2(new_n1000), .A3(new_n1032), .ZN(G393));
  NAND3_X1  g0833(.A1(new_n950), .A2(new_n959), .A3(new_n953), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n667), .B1(new_n1034), .B2(KEYINPUT116), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT116), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n950), .A2(new_n959), .A3(new_n1036), .A4(new_n953), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n961), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT117), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(KEYINPUT117), .A3(new_n961), .A4(new_n1037), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n954), .B(KEYINPUT115), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n999), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n925), .A2(new_n726), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n735), .B1(new_n507), .B2(new_n211), .C1(new_n991), .C2(new_n246), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n759), .A2(new_n409), .B1(new_n757), .B2(new_n203), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n773), .A2(new_n401), .B1(new_n790), .B2(new_n741), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G50), .C2(new_n750), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G150), .A2(new_n747), .B1(new_n739), .B2(G159), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT51), .Z(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1051), .A3(new_n728), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n762), .A2(new_n275), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G317), .A2(new_n747), .B1(new_n739), .B2(G311), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  OAI22_X1  g0855(.A1(new_n773), .A2(new_n763), .B1(new_n757), .B2(new_n767), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G303), .B2(new_n750), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n375), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n760), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n741), .B2(new_n1003), .C1(new_n503), .C2(new_n762), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1052), .A2(new_n1053), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n734), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1045), .A2(new_n719), .A3(new_n1046), .A4(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1042), .A2(new_n1044), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT118), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1063), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT118), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n1044), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1065), .A2(new_n1069), .ZN(G390));
  AOI21_X1  g0870(.A(new_n878), .B1(new_n905), .B2(new_n822), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(KEYINPUT104), .A3(new_n872), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n900), .B1(new_n1074), .B2(new_n899), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n901), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n713), .A2(G330), .A3(new_n785), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n822), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n878), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n783), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n684), .A2(new_n685), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n784), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1081), .B(new_n849), .C1(new_n1085), .C2(new_n1079), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1077), .A2(new_n1080), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n823), .A2(G330), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1071), .B1(new_n877), .B2(new_n901), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1085), .A2(new_n1079), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n849), .A2(new_n1081), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1089), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1087), .A2(new_n1094), .A3(new_n999), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n724), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n375), .B1(new_n748), .B2(new_n767), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1053), .B(new_n1097), .C1(G97), .C2(new_n751), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n759), .A2(new_n203), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n789), .A2(new_n503), .B1(new_n409), .B2(new_n757), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(G107), .C2(new_n750), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1098), .B(new_n1101), .C1(new_n763), .C2(new_n741), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G128), .A2(new_n747), .B1(new_n739), .B2(G132), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT119), .Z(new_n1104));
  OAI221_X1 g0904(.A(new_n253), .B1(new_n759), .B2(new_n201), .C1(new_n764), .C2(new_n791), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT53), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n757), .B2(new_n968), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n795), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n742), .A2(G125), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n773), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1104), .A2(new_n1109), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n762), .A2(new_n1018), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1102), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n734), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n401), .A2(new_n813), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1096), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1095), .B1(new_n720), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n868), .A2(new_n638), .A3(new_n860), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n905), .B1(new_n1089), .B2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n820), .A2(G330), .A3(new_n785), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1085), .B(new_n1080), .C1(new_n822), .C2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1120), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1087), .A2(new_n1094), .A3(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1126), .A2(new_n666), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1087), .A2(new_n1094), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1119), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(G378));
  AND3_X1   g0932(.A1(new_n363), .A2(KEYINPUT89), .A3(new_n368), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT89), .B1(new_n363), .B2(new_n368), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n438), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n353), .A2(new_n356), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n824), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1140));
  NAND3_X1  g0940(.A1(new_n637), .A2(new_n438), .A3(new_n1137), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1140), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n859), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT122), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1140), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(KEYINPUT122), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1153), .A2(G330), .A3(new_n865), .A4(new_n850), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1145), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n908), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1145), .A2(new_n1154), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n902), .A3(new_n907), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n999), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1153), .A2(new_n724), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n739), .A2(G128), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n757), .B2(new_n1111), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n747), .A2(G125), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n968), .B2(new_n762), .C1(new_n764), .C2(new_n797), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G137), .C2(new_n751), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT121), .ZN(new_n1167));
  XOR2_X1   g0967(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1168));
  XNOR2_X1  g0968(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(G41), .B1(new_n742), .B2(G124), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n272), .C1(new_n1018), .C2(new_n759), .ZN(new_n1171));
  AOI21_X1  g0971(.A(G41), .B1(new_n728), .B2(G33), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1169), .A2(new_n1171), .B1(G50), .B2(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n762), .A2(new_n203), .B1(new_n767), .B2(new_n741), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n542), .B2(new_n751), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G41), .B1(new_n972), .B2(G58), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n275), .C2(new_n757), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n728), .B(new_n1177), .C1(G116), .C2(new_n747), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n507), .B2(new_n764), .C1(new_n317), .C2(new_n789), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT58), .Z(new_n1180));
  OAI21_X1  g0980(.A(new_n734), .B1(new_n1173), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n813), .A2(new_n201), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1161), .A2(new_n719), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1160), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1120), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1126), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1157), .A2(KEYINPUT123), .A3(new_n902), .A4(new_n907), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT123), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1156), .A2(new_n1189), .A3(new_n1158), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(KEYINPUT57), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1126), .A2(new_n1186), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n666), .B1(new_n1193), .B2(KEYINPUT57), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1185), .B1(new_n1192), .B2(new_n1194), .ZN(G375));
  NAND2_X1  g0995(.A1(new_n1079), .A2(new_n724), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n253), .B1(new_n750), .B2(G116), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n507), .B2(new_n757), .C1(new_n789), .C2(new_n767), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1017), .B1(G107), .B2(new_n751), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n275), .B2(new_n759), .C1(new_n771), .C2(new_n741), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(G294), .C2(new_n747), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n751), .A2(G150), .B1(G58), .B2(new_n972), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n742), .A2(G128), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n739), .A2(G137), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n728), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n748), .A2(new_n797), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n764), .A2(new_n1111), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n762), .A2(new_n201), .B1(new_n757), .B2(new_n1018), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n734), .B1(new_n1201), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n813), .A2(new_n203), .ZN(new_n1211));
  AND4_X1   g1011(.A1(new_n719), .A2(new_n1196), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1124), .A2(new_n1122), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n999), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1213), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1120), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n963), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1217), .B2(new_n1125), .ZN(G381));
  INV_X1    g1018(.A(new_n993), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n939), .B2(new_n966), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1065), .A2(new_n1220), .A3(new_n1069), .ZN(new_n1221));
  OR2_X1    g1021(.A1(G381), .A2(G384), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1221), .A2(G396), .A3(G393), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1187), .A2(new_n1159), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT57), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n667), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1184), .B1(new_n1226), .B2(new_n1191), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n1131), .A3(new_n1227), .ZN(G407));
  NOR2_X1   g1028(.A1(new_n1223), .A2(new_n646), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1131), .ZN(new_n1230));
  OAI21_X1  g1030(.A(G213), .B1(new_n1229), .B2(new_n1230), .ZN(G409));
  NAND2_X1  g1031(.A1(new_n646), .A2(G213), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1190), .A2(new_n999), .A3(new_n1188), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1183), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT124), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1193), .A2(new_n963), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT124), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1233), .A2(new_n1237), .A3(new_n1183), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1131), .A3(new_n1236), .A4(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1232), .B(new_n1239), .C1(new_n1227), .C2(new_n1131), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1129), .B(new_n666), .C1(new_n1216), .C2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT60), .B1(new_n1215), .B2(new_n1120), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1214), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  XOR2_X1   g1044(.A(G384), .B(KEYINPUT125), .Z(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1214), .B(new_n1247), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT62), .B1(new_n1240), .B2(new_n1250), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n646), .A2(G213), .A3(G2897), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1246), .A2(new_n1252), .A3(new_n1248), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT61), .B1(new_n1240), .B2(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G375), .A2(G378), .B1(G213), .B2(new_n646), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1239), .A4(new_n1249), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1067), .A2(new_n1068), .A3(new_n1044), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1068), .B1(new_n1067), .B2(new_n1044), .ZN(new_n1262));
  OAI21_X1  g1062(.A(G387), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  XOR2_X1   g1063(.A(G393), .B(G396), .Z(new_n1264));
  AND3_X1   g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1221), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1263), .B2(new_n1221), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1260), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1264), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1065), .A2(new_n1220), .A3(new_n1069), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1220), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1263), .A2(new_n1221), .A3(new_n1264), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1240), .A2(new_n1255), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT127), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1240), .A2(new_n1278), .A3(new_n1255), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1274), .A2(new_n1276), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT126), .B1(new_n1240), .B2(new_n1250), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT63), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  OAI211_X1 g1083(.A(KEYINPUT126), .B(new_n1283), .C1(new_n1240), .C2(new_n1250), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1268), .B1(new_n1280), .B2(new_n1285), .ZN(G405));
  NAND2_X1  g1086(.A1(G375), .A2(G378), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1230), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1250), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1230), .A2(new_n1287), .A3(new_n1249), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1267), .B(new_n1291), .ZN(G402));
endmodule


