

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U558 ( .A(n667), .ZN(n635) );
  NOR2_X1 U559 ( .A1(G651), .A2(n534), .ZN(n806) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n729) );
  NAND2_X2 U561 ( .A1(n729), .A2(n728), .ZN(n667) );
  XNOR2_X1 U562 ( .A(n610), .B(KEYINPUT31), .ZN(n611) );
  NOR2_X1 U563 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U564 ( .A1(n674), .A2(n673), .ZN(n676) );
  XNOR2_X1 U565 ( .A(KEYINPUT105), .B(n774), .ZN(n524) );
  OR2_X1 U566 ( .A1(n773), .A2(n761), .ZN(n525) );
  XOR2_X1 U567 ( .A(n727), .B(KEYINPUT102), .Z(n526) );
  INV_X1 U568 ( .A(KEYINPUT94), .ZN(n644) );
  XNOR2_X1 U569 ( .A(n645), .B(n644), .ZN(n653) );
  INV_X1 U570 ( .A(KEYINPUT98), .ZN(n610) );
  INV_X1 U571 ( .A(KEYINPUT96), .ZN(n662) );
  XNOR2_X1 U572 ( .A(n612), .B(n611), .ZN(n665) );
  INV_X1 U573 ( .A(KEYINPUT32), .ZN(n675) );
  NAND2_X1 U574 ( .A1(G8), .A2(n667), .ZN(n710) );
  NOR2_X1 U575 ( .A1(n1000), .A2(n689), .ZN(n690) );
  NOR2_X1 U576 ( .A1(n555), .A2(G2104), .ZN(n902) );
  AND2_X1 U577 ( .A1(n555), .A2(G2104), .ZN(n907) );
  NOR2_X1 U578 ( .A1(n600), .A2(n599), .ZN(G160) );
  XNOR2_X1 U579 ( .A(n776), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U580 ( .A(G651), .ZN(n533) );
  NOR2_X1 U581 ( .A1(n533), .A2(G543), .ZN(n527) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n527), .Z(n624) );
  BUF_X1 U583 ( .A(n624), .Z(n801) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n534) );
  NAND2_X1 U585 ( .A1(G49), .A2(n806), .ZN(n529) );
  NAND2_X1 U586 ( .A1(G74), .A2(G651), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U588 ( .A1(n801), .A2(n530), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n534), .A2(G87), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(G288) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n802) );
  NAND2_X1 U592 ( .A1(G88), .A2(n802), .ZN(n536) );
  NOR2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n805) );
  NAND2_X1 U594 ( .A1(G75), .A2(n805), .ZN(n535) );
  NAND2_X1 U595 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U596 ( .A(KEYINPUT78), .B(n537), .ZN(n540) );
  NAND2_X1 U597 ( .A1(G62), .A2(n801), .ZN(n538) );
  XNOR2_X1 U598 ( .A(KEYINPUT77), .B(n538), .ZN(n539) );
  NOR2_X1 U599 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n806), .A2(G50), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(G303) );
  NAND2_X1 U602 ( .A1(G64), .A2(n801), .ZN(n544) );
  NAND2_X1 U603 ( .A1(G52), .A2(n806), .ZN(n543) );
  NAND2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U605 ( .A(KEYINPUT65), .B(n545), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n802), .A2(G90), .ZN(n546) );
  XNOR2_X1 U607 ( .A(n546), .B(KEYINPUT66), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G77), .A2(n805), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n549) );
  XNOR2_X1 U611 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U613 ( .A(KEYINPUT68), .B(n553), .ZN(G301) );
  NOR2_X1 U614 ( .A1(G2105), .A2(G2104), .ZN(n554) );
  XOR2_X2 U615 ( .A(KEYINPUT17), .B(n554), .Z(n906) );
  NAND2_X1 U616 ( .A1(G138), .A2(n906), .ZN(n561) );
  INV_X1 U617 ( .A(G2105), .ZN(n555) );
  AND2_X1 U618 ( .A1(G102), .A2(n907), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G126), .A2(n902), .ZN(n557) );
  AND2_X1 U620 ( .A1(G2105), .A2(G2104), .ZN(n903) );
  NAND2_X1 U621 ( .A1(G114), .A2(n903), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  AND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(G164) );
  NAND2_X1 U625 ( .A1(n802), .A2(G89), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G76), .A2(n805), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G63), .A2(n801), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G51), .A2(n806), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U636 ( .A1(G78), .A2(n805), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT70), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G65), .A2(n801), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G53), .A2(n806), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G91), .A2(n802), .ZN(n575) );
  XNOR2_X1 U642 ( .A(KEYINPUT69), .B(n575), .ZN(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(G299) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U646 ( .A1(G48), .A2(n806), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT76), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G61), .A2(n801), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G86), .A2(n802), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n805), .A2(G73), .ZN(n583) );
  XOR2_X1 U652 ( .A(KEYINPUT2), .B(n583), .Z(n584) );
  NOR2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U655 ( .A1(G85), .A2(n802), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G72), .A2(n805), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U658 ( .A1(G60), .A2(n801), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G47), .A2(n806), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n592) );
  OR2_X1 U661 ( .A1(n593), .A2(n592), .ZN(G290) );
  AND2_X1 U662 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  NOR2_X1 U663 ( .A1(G1971), .A2(G303), .ZN(n688) );
  XOR2_X1 U664 ( .A(G2078), .B(KEYINPUT25), .Z(n970) );
  NAND2_X1 U665 ( .A1(n902), .A2(G125), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G101), .A2(n907), .ZN(n594) );
  XOR2_X1 U667 ( .A(KEYINPUT23), .B(n594), .Z(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G137), .A2(n906), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G113), .A2(n903), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X1 U672 ( .A1(G160), .A2(G40), .ZN(n728) );
  NOR2_X1 U673 ( .A1(n970), .A2(n667), .ZN(n602) );
  XOR2_X1 U674 ( .A(G1961), .B(KEYINPUT91), .Z(n1014) );
  NOR2_X1 U675 ( .A1(n635), .A2(n1014), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n659) );
  AND2_X1 U677 ( .A1(G301), .A2(n659), .ZN(n609) );
  XOR2_X1 U678 ( .A(KEYINPUT97), .B(KEYINPUT30), .Z(n606) );
  NOR2_X1 U679 ( .A1(G2084), .A2(n667), .ZN(n677) );
  NOR2_X1 U680 ( .A1(n710), .A2(G1966), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT90), .ZN(n681) );
  NOR2_X1 U682 ( .A1(n677), .A2(n681), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n604), .A2(G8), .ZN(n605) );
  XNOR2_X1 U684 ( .A(n606), .B(n605), .ZN(n607) );
  NOR2_X1 U685 ( .A1(G168), .A2(n607), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n635), .A2(G1348), .ZN(n614) );
  NOR2_X1 U687 ( .A1(G2067), .A2(n667), .ZN(n613) );
  NOR2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n623) );
  NAND2_X1 U689 ( .A1(G66), .A2(n624), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G92), .A2(n802), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U692 ( .A(KEYINPUT72), .B(n617), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G79), .A2(n805), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G54), .A2(n806), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U697 ( .A(KEYINPUT15), .B(n622), .Z(n992) );
  INV_X1 U698 ( .A(n992), .ZN(n780) );
  OR2_X1 U699 ( .A1(n623), .A2(n780), .ZN(n643) );
  NAND2_X1 U700 ( .A1(n780), .A2(n623), .ZN(n641) );
  NAND2_X1 U701 ( .A1(n624), .A2(G56), .ZN(n625) );
  XNOR2_X1 U702 ( .A(KEYINPUT14), .B(n625), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n802), .A2(G81), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n626), .B(KEYINPUT12), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G68), .A2(n805), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U707 ( .A(KEYINPUT13), .B(n629), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT71), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n806), .A2(G43), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n999) );
  NAND2_X1 U712 ( .A1(n635), .A2(G1996), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n636), .B(KEYINPUT26), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n667), .A2(G1341), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U716 ( .A1(n999), .A2(n639), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n645) );
  INV_X1 U719 ( .A(G2072), .ZN(n939) );
  NOR2_X1 U720 ( .A1(n667), .A2(n939), .ZN(n648) );
  XOR2_X1 U721 ( .A(KEYINPUT93), .B(KEYINPUT27), .Z(n646) );
  XNOR2_X1 U722 ( .A(KEYINPUT92), .B(n646), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n648), .B(n647), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n667), .A2(G1956), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(n654) );
  NOR2_X1 U726 ( .A1(G299), .A2(n654), .ZN(n651) );
  XNOR2_X1 U727 ( .A(KEYINPUT95), .B(n651), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U729 ( .A1(G299), .A2(n654), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n655), .B(KEYINPUT28), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(KEYINPUT29), .ZN(n661) );
  NOR2_X1 U733 ( .A1(G301), .A2(n659), .ZN(n660) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n679) );
  AND2_X1 U737 ( .A1(G286), .A2(G8), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n679), .A2(n666), .ZN(n674) );
  INV_X1 U739 ( .A(G8), .ZN(n672) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n710), .ZN(n669) );
  NOR2_X1 U741 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(G303), .ZN(n671) );
  OR2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U745 ( .A(n676), .B(n675), .ZN(n685) );
  NAND2_X1 U746 ( .A1(G8), .A2(n677), .ZN(n678) );
  XOR2_X1 U747 ( .A(KEYINPUT89), .B(n678), .Z(n683) );
  INV_X1 U748 ( .A(n679), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n709) );
  NOR2_X1 U752 ( .A1(G288), .A2(G1976), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n686), .B(KEYINPUT99), .ZN(n719) );
  NAND2_X1 U754 ( .A1(n709), .A2(n719), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n690), .B(KEYINPUT64), .ZN(n693) );
  INV_X1 U757 ( .A(n710), .ZN(n691) );
  AND2_X1 U758 ( .A1(n691), .A2(KEYINPUT100), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n716) );
  INV_X1 U760 ( .A(KEYINPUT100), .ZN(n694) );
  INV_X1 U761 ( .A(KEYINPUT33), .ZN(n696) );
  OR2_X1 U762 ( .A1(n694), .A2(n696), .ZN(n703) );
  XNOR2_X1 U763 ( .A(G1981), .B(KEYINPUT101), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n695), .B(G305), .ZN(n989) );
  INV_X1 U765 ( .A(n989), .ZN(n702) );
  NAND2_X1 U766 ( .A1(n696), .A2(KEYINPUT64), .ZN(n700) );
  NOR2_X1 U767 ( .A1(KEYINPUT100), .A2(n719), .ZN(n697) );
  NAND2_X1 U768 ( .A1(KEYINPUT33), .A2(n697), .ZN(n698) );
  NAND2_X1 U769 ( .A1(n698), .A2(n691), .ZN(n699) );
  NAND2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n701) );
  OR2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n718) );
  AND2_X1 U772 ( .A1(n703), .A2(n718), .ZN(n714) );
  NOR2_X1 U773 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XOR2_X1 U774 ( .A(n704), .B(KEYINPUT88), .Z(n705) );
  XNOR2_X1 U775 ( .A(KEYINPUT24), .B(n705), .ZN(n706) );
  OR2_X1 U776 ( .A1(n710), .A2(n706), .ZN(n713) );
  NOR2_X1 U777 ( .A1(G2090), .A2(G303), .ZN(n707) );
  NAND2_X1 U778 ( .A1(G8), .A2(n707), .ZN(n708) );
  NAND2_X1 U779 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n717) );
  AND2_X1 U782 ( .A1(n714), .A2(n717), .ZN(n715) );
  NAND2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n726) );
  INV_X1 U784 ( .A(n717), .ZN(n724) );
  INV_X1 U785 ( .A(n718), .ZN(n722) );
  INV_X1 U786 ( .A(n719), .ZN(n1001) );
  NAND2_X1 U787 ( .A1(n1001), .A2(KEYINPUT33), .ZN(n720) );
  AND2_X1 U788 ( .A1(n720), .A2(n989), .ZN(n721) );
  OR2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n723) );
  OR2_X1 U790 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n727) );
  INV_X1 U792 ( .A(n728), .ZN(n730) );
  NOR2_X1 U793 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U794 ( .A(n731), .B(KEYINPUT83), .ZN(n773) );
  NAND2_X1 U795 ( .A1(G141), .A2(n906), .ZN(n732) );
  XNOR2_X1 U796 ( .A(n732), .B(KEYINPUT87), .ZN(n735) );
  NAND2_X1 U797 ( .A1(G129), .A2(n902), .ZN(n733) );
  XOR2_X1 U798 ( .A(KEYINPUT84), .B(n733), .Z(n734) );
  NOR2_X1 U799 ( .A1(n735), .A2(n734), .ZN(n742) );
  XOR2_X1 U800 ( .A(KEYINPUT86), .B(KEYINPUT38), .Z(n737) );
  NAND2_X1 U801 ( .A1(G105), .A2(n907), .ZN(n736) );
  XNOR2_X1 U802 ( .A(n737), .B(n736), .ZN(n740) );
  NAND2_X1 U803 ( .A1(G117), .A2(n903), .ZN(n738) );
  XNOR2_X1 U804 ( .A(KEYINPUT85), .B(n738), .ZN(n739) );
  NOR2_X1 U805 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U806 ( .A1(n742), .A2(n741), .ZN(n927) );
  NAND2_X1 U807 ( .A1(G1996), .A2(n927), .ZN(n750) );
  NAND2_X1 U808 ( .A1(G131), .A2(n906), .ZN(n744) );
  NAND2_X1 U809 ( .A1(G95), .A2(n907), .ZN(n743) );
  NAND2_X1 U810 ( .A1(n744), .A2(n743), .ZN(n748) );
  NAND2_X1 U811 ( .A1(G119), .A2(n902), .ZN(n746) );
  NAND2_X1 U812 ( .A1(G107), .A2(n903), .ZN(n745) );
  NAND2_X1 U813 ( .A1(n746), .A2(n745), .ZN(n747) );
  OR2_X1 U814 ( .A1(n748), .A2(n747), .ZN(n920) );
  NAND2_X1 U815 ( .A1(G1991), .A2(n920), .ZN(n749) );
  NAND2_X1 U816 ( .A1(n750), .A2(n749), .ZN(n944) );
  XOR2_X1 U817 ( .A(G1986), .B(G290), .Z(n998) );
  XOR2_X1 U818 ( .A(G2067), .B(KEYINPUT37), .Z(n762) );
  NAND2_X1 U819 ( .A1(G128), .A2(n902), .ZN(n752) );
  NAND2_X1 U820 ( .A1(G116), .A2(n903), .ZN(n751) );
  NAND2_X1 U821 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U822 ( .A(n753), .B(KEYINPUT35), .ZN(n758) );
  NAND2_X1 U823 ( .A1(G140), .A2(n906), .ZN(n755) );
  NAND2_X1 U824 ( .A1(G104), .A2(n907), .ZN(n754) );
  NAND2_X1 U825 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U826 ( .A(KEYINPUT34), .B(n756), .Z(n757) );
  NAND2_X1 U827 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U828 ( .A(n759), .B(KEYINPUT36), .ZN(n928) );
  NAND2_X1 U829 ( .A1(n762), .A2(n928), .ZN(n954) );
  NAND2_X1 U830 ( .A1(n998), .A2(n954), .ZN(n760) );
  NOR2_X1 U831 ( .A1(n944), .A2(n760), .ZN(n761) );
  NAND2_X1 U832 ( .A1(n526), .A2(n525), .ZN(n775) );
  NOR2_X1 U833 ( .A1(n762), .A2(n928), .ZN(n945) );
  INV_X1 U834 ( .A(n954), .ZN(n770) );
  NOR2_X1 U835 ( .A1(G1996), .A2(n927), .ZN(n763) );
  XOR2_X1 U836 ( .A(KEYINPUT103), .B(n763), .Z(n957) );
  NOR2_X1 U837 ( .A1(G1986), .A2(G290), .ZN(n764) );
  NOR2_X1 U838 ( .A1(G1991), .A2(n920), .ZN(n952) );
  NOR2_X1 U839 ( .A1(n764), .A2(n952), .ZN(n765) );
  NOR2_X1 U840 ( .A1(n944), .A2(n765), .ZN(n766) );
  XNOR2_X1 U841 ( .A(n766), .B(KEYINPUT104), .ZN(n767) );
  NOR2_X1 U842 ( .A1(n957), .A2(n767), .ZN(n768) );
  XOR2_X1 U843 ( .A(KEYINPUT39), .B(n768), .Z(n769) );
  NOR2_X1 U844 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U845 ( .A1(n945), .A2(n771), .ZN(n772) );
  NOR2_X1 U846 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U847 ( .A1(n775), .A2(n524), .ZN(n776) );
  AND2_X1 U848 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U849 ( .A(G132), .ZN(G219) );
  INV_X1 U850 ( .A(G82), .ZN(G220) );
  INV_X1 U851 ( .A(G120), .ZN(G236) );
  INV_X1 U852 ( .A(G69), .ZN(G235) );
  INV_X1 U853 ( .A(G108), .ZN(G238) );
  NAND2_X1 U854 ( .A1(G7), .A2(G661), .ZN(n778) );
  XNOR2_X1 U855 ( .A(n778), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U856 ( .A(G223), .ZN(n855) );
  NAND2_X1 U857 ( .A1(n855), .A2(G567), .ZN(n779) );
  XOR2_X1 U858 ( .A(KEYINPUT11), .B(n779), .Z(G234) );
  INV_X1 U859 ( .A(G860), .ZN(n785) );
  OR2_X1 U860 ( .A1(n999), .A2(n785), .ZN(G153) );
  NAND2_X1 U861 ( .A1(G301), .A2(G868), .ZN(n782) );
  INV_X1 U862 ( .A(G868), .ZN(n822) );
  NAND2_X1 U863 ( .A1(n780), .A2(n822), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n782), .A2(n781), .ZN(G284) );
  NOR2_X1 U865 ( .A1(G286), .A2(n822), .ZN(n784) );
  NOR2_X1 U866 ( .A1(G868), .A2(G299), .ZN(n783) );
  NOR2_X1 U867 ( .A1(n784), .A2(n783), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n785), .A2(G559), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n786), .A2(n992), .ZN(n787) );
  XNOR2_X1 U870 ( .A(n787), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U871 ( .A1(G868), .A2(n999), .ZN(n790) );
  NAND2_X1 U872 ( .A1(G868), .A2(n992), .ZN(n788) );
  NOR2_X1 U873 ( .A1(G559), .A2(n788), .ZN(n789) );
  NOR2_X1 U874 ( .A1(n790), .A2(n789), .ZN(G282) );
  NAND2_X1 U875 ( .A1(G123), .A2(n902), .ZN(n791) );
  XNOR2_X1 U876 ( .A(n791), .B(KEYINPUT18), .ZN(n798) );
  NAND2_X1 U877 ( .A1(G135), .A2(n906), .ZN(n793) );
  NAND2_X1 U878 ( .A1(G111), .A2(n903), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G99), .A2(n907), .ZN(n794) );
  XNOR2_X1 U881 ( .A(KEYINPUT73), .B(n794), .ZN(n795) );
  NOR2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n949) );
  XNOR2_X1 U884 ( .A(G2096), .B(n949), .ZN(n799) );
  NOR2_X1 U885 ( .A1(G2100), .A2(n799), .ZN(n800) );
  XOR2_X1 U886 ( .A(KEYINPUT74), .B(n800), .Z(G156) );
  NAND2_X1 U887 ( .A1(G67), .A2(n801), .ZN(n804) );
  NAND2_X1 U888 ( .A1(G93), .A2(n802), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n804), .A2(n803), .ZN(n810) );
  NAND2_X1 U890 ( .A1(G80), .A2(n805), .ZN(n808) );
  NAND2_X1 U891 ( .A1(G55), .A2(n806), .ZN(n807) );
  NAND2_X1 U892 ( .A1(n808), .A2(n807), .ZN(n809) );
  OR2_X1 U893 ( .A1(n810), .A2(n809), .ZN(n823) );
  NAND2_X1 U894 ( .A1(n992), .A2(G559), .ZN(n820) );
  XNOR2_X1 U895 ( .A(n999), .B(n820), .ZN(n811) );
  NOR2_X1 U896 ( .A1(G860), .A2(n811), .ZN(n812) );
  XOR2_X1 U897 ( .A(KEYINPUT75), .B(n812), .Z(n813) );
  XOR2_X1 U898 ( .A(n823), .B(n813), .Z(G145) );
  INV_X1 U899 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U900 ( .A(n823), .B(KEYINPUT19), .ZN(n814) );
  XNOR2_X1 U901 ( .A(G288), .B(n814), .ZN(n817) );
  XNOR2_X1 U902 ( .A(G166), .B(G299), .ZN(n815) );
  XNOR2_X1 U903 ( .A(n815), .B(G305), .ZN(n816) );
  XNOR2_X1 U904 ( .A(n817), .B(n816), .ZN(n818) );
  XNOR2_X1 U905 ( .A(n818), .B(G290), .ZN(n819) );
  XNOR2_X1 U906 ( .A(n999), .B(n819), .ZN(n864) );
  XNOR2_X1 U907 ( .A(n820), .B(n864), .ZN(n821) );
  NAND2_X1 U908 ( .A1(n821), .A2(G868), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U910 ( .A1(n825), .A2(n824), .ZN(G295) );
  NAND2_X1 U911 ( .A1(G2084), .A2(G2078), .ZN(n826) );
  XOR2_X1 U912 ( .A(KEYINPUT20), .B(n826), .Z(n827) );
  NAND2_X1 U913 ( .A1(G2090), .A2(n827), .ZN(n829) );
  XOR2_X1 U914 ( .A(KEYINPUT79), .B(KEYINPUT21), .Z(n828) );
  XNOR2_X1 U915 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U916 ( .A1(G2072), .A2(n830), .ZN(G158) );
  XNOR2_X1 U917 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U918 ( .A1(G235), .A2(G236), .ZN(n831) );
  XNOR2_X1 U919 ( .A(n831), .B(KEYINPUT81), .ZN(n832) );
  NOR2_X1 U920 ( .A1(G238), .A2(n832), .ZN(n833) );
  NAND2_X1 U921 ( .A1(G57), .A2(n833), .ZN(n861) );
  NAND2_X1 U922 ( .A1(G567), .A2(n861), .ZN(n839) );
  NOR2_X1 U923 ( .A1(G220), .A2(G219), .ZN(n834) );
  XOR2_X1 U924 ( .A(KEYINPUT22), .B(n834), .Z(n835) );
  NOR2_X1 U925 ( .A1(G218), .A2(n835), .ZN(n836) );
  XNOR2_X1 U926 ( .A(KEYINPUT80), .B(n836), .ZN(n837) );
  NAND2_X1 U927 ( .A1(n837), .A2(G96), .ZN(n862) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n862), .ZN(n838) );
  NAND2_X1 U929 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U930 ( .A(KEYINPUT82), .B(n840), .Z(G319) );
  INV_X1 U931 ( .A(G319), .ZN(n842) );
  NAND2_X1 U932 ( .A1(G661), .A2(G483), .ZN(n841) );
  NOR2_X1 U933 ( .A1(n842), .A2(n841), .ZN(n860) );
  NAND2_X1 U934 ( .A1(n860), .A2(G36), .ZN(G176) );
  XNOR2_X1 U935 ( .A(G1348), .B(G1341), .ZN(n843) );
  XNOR2_X1 U936 ( .A(n843), .B(KEYINPUT106), .ZN(n853) );
  XOR2_X1 U937 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n845) );
  XNOR2_X1 U938 ( .A(G2443), .B(G2446), .ZN(n844) );
  XNOR2_X1 U939 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U940 ( .A(G2435), .B(G2438), .Z(n847) );
  XNOR2_X1 U941 ( .A(G2454), .B(G2430), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U943 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U944 ( .A(G2451), .B(G2427), .ZN(n850) );
  XNOR2_X1 U945 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U946 ( .A(n853), .B(n852), .ZN(n854) );
  NAND2_X1 U947 ( .A1(n854), .A2(G14), .ZN(n933) );
  XNOR2_X1 U948 ( .A(KEYINPUT109), .B(n933), .ZN(G401) );
  NAND2_X1 U949 ( .A1(G2106), .A2(n855), .ZN(G217) );
  INV_X1 U950 ( .A(G661), .ZN(n857) );
  NAND2_X1 U951 ( .A1(G2), .A2(G15), .ZN(n856) );
  NOR2_X1 U952 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U953 ( .A(KEYINPUT110), .B(n858), .Z(G259) );
  NAND2_X1 U954 ( .A1(G3), .A2(G1), .ZN(n859) );
  NAND2_X1 U955 ( .A1(n860), .A2(n859), .ZN(G188) );
  INV_X1 U957 ( .A(G96), .ZN(G221) );
  NOR2_X1 U958 ( .A1(n862), .A2(n861), .ZN(G325) );
  INV_X1 U959 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U960 ( .A(G301), .B(n992), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n863), .B(G286), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n866) );
  NOR2_X1 U963 ( .A1(G37), .A2(n866), .ZN(G397) );
  XOR2_X1 U964 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n868) );
  XNOR2_X1 U965 ( .A(G2678), .B(KEYINPUT111), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U967 ( .A(KEYINPUT43), .B(G2090), .Z(n870) );
  XNOR2_X1 U968 ( .A(G2067), .B(G2072), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U970 ( .A(n872), .B(n871), .Z(n874) );
  XNOR2_X1 U971 ( .A(G2096), .B(G2100), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n876) );
  XOR2_X1 U973 ( .A(G2084), .B(G2078), .Z(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(G227) );
  XOR2_X1 U975 ( .A(G2474), .B(G1981), .Z(n878) );
  XNOR2_X1 U976 ( .A(G1986), .B(G1961), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U978 ( .A(n879), .B(KEYINPUT114), .Z(n881) );
  XNOR2_X1 U979 ( .A(G1996), .B(G1991), .ZN(n880) );
  XNOR2_X1 U980 ( .A(n881), .B(n880), .ZN(n885) );
  XOR2_X1 U981 ( .A(G1976), .B(G1971), .Z(n883) );
  XNOR2_X1 U982 ( .A(G1966), .B(G1956), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(n885), .B(n884), .Z(n887) );
  XNOR2_X1 U985 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(G229) );
  NAND2_X1 U987 ( .A1(n902), .A2(G124), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n888), .B(KEYINPUT44), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G112), .A2(n903), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G136), .A2(n906), .ZN(n892) );
  NAND2_X1 U992 ( .A1(G100), .A2(n907), .ZN(n891) );
  NAND2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(G162) );
  NAND2_X1 U995 ( .A1(G139), .A2(n906), .ZN(n896) );
  NAND2_X1 U996 ( .A1(G103), .A2(n907), .ZN(n895) );
  NAND2_X1 U997 ( .A1(n896), .A2(n895), .ZN(n901) );
  NAND2_X1 U998 ( .A1(G127), .A2(n902), .ZN(n898) );
  NAND2_X1 U999 ( .A1(G115), .A2(n903), .ZN(n897) );
  NAND2_X1 U1000 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U1001 ( .A(KEYINPUT47), .B(n899), .Z(n900) );
  NOR2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n940) );
  NAND2_X1 U1003 ( .A1(G130), .A2(n902), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(G118), .A2(n903), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n912) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n906), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(G106), .A2(n907), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1009 ( .A(KEYINPUT45), .B(n910), .Z(n911) );
  NOR2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n922) );
  XOR2_X1 U1011 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(KEYINPUT118), .B(n915), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n949), .B(KEYINPUT117), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1017 ( .A(G164), .B(n918), .Z(n919) );
  XNOR2_X1 U1018 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1019 ( .A(n922), .B(n921), .Z(n924) );
  XNOR2_X1 U1020 ( .A(G160), .B(G162), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1022 ( .A(n940), .B(n925), .Z(n926) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(n929), .B(n928), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(G37), .A2(n930), .ZN(G395) );
  NOR2_X1 U1026 ( .A1(G227), .A2(G229), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT49), .B(n931), .Z(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(G397), .A2(n934), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(G319), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n936), .A2(G395), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(n937), .B(KEYINPUT119), .ZN(G225) );
  INV_X1 U1033 ( .A(G225), .ZN(G308) );
  INV_X1 U1034 ( .A(G301), .ZN(G171) );
  INV_X1 U1035 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1036 ( .A(G164), .B(G2078), .Z(n938) );
  XNOR2_X1 U1037 ( .A(KEYINPUT122), .B(n938), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(n940), .B(n939), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(KEYINPUT50), .B(n943), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n962) );
  XNOR2_X1 U1043 ( .A(G160), .B(G2084), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(n948), .B(KEYINPUT120), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(n955), .B(KEYINPUT121), .ZN(n960) );
  XOR2_X1 U1049 ( .A(G2090), .B(G162), .Z(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1051 ( .A(KEYINPUT51), .B(n958), .Z(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(KEYINPUT52), .B(n963), .ZN(n964) );
  INV_X1 U1055 ( .A(KEYINPUT55), .ZN(n985) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n985), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n965), .A2(G29), .ZN(n1043) );
  XOR2_X1 U1058 ( .A(G2090), .B(G35), .Z(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT123), .B(n966), .ZN(n979) );
  XOR2_X1 U1060 ( .A(G1991), .B(G25), .Z(n967) );
  NAND2_X1 U1061 ( .A1(n967), .A2(G28), .ZN(n976) );
  XNOR2_X1 U1062 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(G33), .B(G2072), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(G1996), .B(G32), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G27), .B(n970), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n977), .B(KEYINPUT53), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n980), .B(KEYINPUT124), .ZN(n983) );
  XOR2_X1 U1073 ( .A(G2084), .B(G34), .Z(n981) );
  XNOR2_X1 U1074 ( .A(KEYINPUT54), .B(n981), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(n985), .B(n984), .ZN(n987) );
  INV_X1 U1077 ( .A(G29), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(G11), .A2(n988), .ZN(n1041) );
  XNOR2_X1 U1080 ( .A(G16), .B(KEYINPUT56), .ZN(n1013) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G168), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n991), .B(KEYINPUT57), .ZN(n1011) );
  XNOR2_X1 U1084 ( .A(G1348), .B(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(G171), .B(G1961), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G299), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1009) );
  XOR2_X1 U1090 ( .A(n999), .B(G1341), .Z(n1007) );
  XNOR2_X1 U1091 ( .A(G303), .B(G1971), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT125), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT126), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1039) );
  INV_X1 U1100 ( .A(G16), .ZN(n1037) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(n1014), .B(G5), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1027) );
  XNOR2_X1 U1104 ( .A(KEYINPUT59), .B(KEYINPUT127), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(n1017), .B(G4), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G1348), .B(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G1981), .B(G6), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(G1956), .B(G20), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(G19), .B(G1341), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1113 ( .A(KEYINPUT60), .B(n1025), .Z(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1034) );
  XNOR2_X1 U1115 ( .A(G1986), .B(G24), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(G1971), .B(G22), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  XOR2_X1 U1118 ( .A(G1976), .B(G23), .Z(n1030) );
  NAND2_X1 U1119 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1120 ( .A(KEYINPUT58), .B(n1032), .ZN(n1033) );
  NOR2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1122 ( .A(KEYINPUT61), .B(n1035), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1126 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1127 ( .A(KEYINPUT62), .B(n1044), .Z(G311) );
  INV_X1 U1128 ( .A(G311), .ZN(G150) );
endmodule

