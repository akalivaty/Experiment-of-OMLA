//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G567), .ZN(new_n460));
  INV_X1    g035(.A(G2106), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT66), .Z(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(KEYINPUT67), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n468), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n464), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n470), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n476), .A2(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n477), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n468), .A2(new_n473), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n500), .A3(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n495), .A2(new_n496), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n496), .B1(new_n495), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(KEYINPUT69), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n510), .B2(G50), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT70), .B(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n515), .A2(new_n525), .ZN(G166));
  XOR2_X1   g101(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n518), .A2(new_n519), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n519), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n531), .A2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n523), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT72), .B(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n532), .A2(new_n540), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n539), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AOI22_X1  g119(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n523), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT73), .B(G43), .Z(new_n548));
  OAI22_X1  g123(.A1(new_n532), .A2(new_n547), .B1(new_n534), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  XNOR2_X1  g130(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n534), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n510), .A2(G53), .A3(new_n559), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n558), .A2(KEYINPUT75), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(KEYINPUT75), .B1(new_n558), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n520), .A2(G91), .ZN(new_n564));
  INV_X1    g139(.A(G78), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT76), .B1(new_n565), .B2(new_n507), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n567), .A2(G78), .A3(G543), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n518), .A2(G65), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n569), .A2(new_n570), .ZN(new_n573));
  NOR3_X1   g148(.A1(new_n572), .A2(KEYINPUT78), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  INV_X1    g150(.A(new_n573), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n523), .B1(new_n569), .B2(new_n570), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n563), .B(new_n564), .C1(new_n574), .C2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(G166), .ZN(G303));
  OR2_X1    g156(.A1(new_n518), .A2(G74), .ZN(new_n582));
  AOI22_X1  g157(.A1(G651), .A2(new_n582), .B1(new_n520), .B2(G87), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n534), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n510), .A2(KEYINPUT79), .A3(G49), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n583), .A2(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n523), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n520), .A2(G86), .B1(G48), .B2(new_n510), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n520), .A2(G85), .B1(G47), .B2(new_n510), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n523), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT80), .ZN(G290));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NOR2_X1   g173(.A1(G301), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n518), .A2(new_n519), .A3(G92), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(new_n518), .ZN(new_n603));
  XOR2_X1   g178(.A(KEYINPUT81), .B(G66), .Z(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT82), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT83), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n601), .A2(new_n606), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT82), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n599), .B1(new_n614), .B2(new_n598), .ZN(G284));
  AOI21_X1  g190(.A(new_n599), .B1(new_n614), .B2(new_n598), .ZN(G321));
  AOI21_X1  g191(.A(G868), .B1(G299), .B2(KEYINPUT85), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(KEYINPUT85), .B2(G299), .ZN(new_n618));
  NOR2_X1   g193(.A1(G168), .A2(new_n598), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT84), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(G297));
  NAND2_X1  g196(.A1(new_n618), .A2(new_n620), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n614), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n477), .A2(G135), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT86), .ZN(new_n633));
  AOI211_X1 g208(.A(new_n631), .B(new_n633), .C1(G123), .C2(new_n484), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2096), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n468), .A2(new_n473), .A3(new_n479), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT87), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n659), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n639), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(G2096), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n673), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n673), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  OR2_X1    g263(.A1(G6), .A2(G16), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(G305), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT32), .B(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(G23), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G288), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT33), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT90), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n697), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n693), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n690), .A2(G22), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n690), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1971), .ZN(new_n703));
  OAI21_X1  g278(.A(KEYINPUT34), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT91), .Z(new_n705));
  INV_X1    g280(.A(KEYINPUT36), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n484), .A2(G119), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT88), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n477), .A2(G131), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n464), .A2(G107), .ZN(new_n710));
  OAI21_X1  g285(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n708), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G25), .B(new_n712), .S(G29), .Z(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n690), .A2(G24), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G290), .B2(G16), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT89), .B(G1986), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n715), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n700), .A2(new_n703), .A3(KEYINPUT34), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n705), .A2(new_n706), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n706), .B1(new_n705), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G19), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n550), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT92), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1341), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G26), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n484), .A2(G128), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n738));
  INV_X1    g313(.A(G116), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G2105), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n477), .B2(G140), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n734), .B1(new_n743), .B2(new_n732), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2067), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n731), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n690), .B1(new_n609), .B2(new_n613), .ZN(new_n747));
  NOR2_X1   g322(.A1(G4), .A2(G16), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n747), .A2(G1348), .A3(new_n748), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n746), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT94), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(KEYINPUT94), .B(new_n746), .C1(new_n751), .C2(new_n752), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT25), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n477), .A2(G139), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n468), .A2(new_n473), .A3(G127), .ZN(new_n761));
  NAND2_X1  g336(.A1(G115), .A2(G2104), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n464), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G33), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(G29), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(G2072), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT95), .Z(new_n770));
  OR2_X1    g345(.A1(G29), .A2(G32), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT98), .B(KEYINPUT26), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(KEYINPUT26), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT26), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n773), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n775), .A2(new_n780), .B1(G105), .B2(new_n479), .ZN(new_n781));
  AOI22_X1  g356(.A1(G129), .A2(new_n484), .B1(new_n477), .B2(G141), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT99), .ZN(new_n783));
  AOI21_X1  g358(.A(KEYINPUT99), .B1(new_n781), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT100), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n771), .B1(new_n786), .B2(new_n732), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT27), .B(G1996), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n770), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G11), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT31), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(KEYINPUT31), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n795), .A2(G28), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n732), .B1(new_n795), .B2(G28), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n793), .B(new_n794), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n634), .B2(G29), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n690), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n690), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G1961), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G1966), .ZN(new_n804));
  INV_X1    g379(.A(G21), .ZN(new_n805));
  AOI21_X1  g380(.A(KEYINPUT101), .B1(new_n690), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G286), .B2(new_n690), .ZN(new_n807));
  NAND3_X1  g382(.A1(G168), .A2(KEYINPUT101), .A3(G16), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n801), .A2(G1961), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n803), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n732), .A2(G35), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G162), .B2(new_n732), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT29), .ZN(new_n814));
  INV_X1    g389(.A(G2090), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(KEYINPUT29), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n815), .B1(new_n814), .B2(new_n816), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT24), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n732), .B1(new_n819), .B2(G34), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT96), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(KEYINPUT96), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n819), .A2(G34), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT97), .Z(new_n825));
  INV_X1    g400(.A(G160), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n732), .ZN(new_n827));
  INV_X1    g402(.A(G2084), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n817), .A2(new_n818), .A3(new_n829), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n768), .A2(G2072), .B1(new_n828), .B2(new_n827), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n811), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(G299), .A2(G16), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n690), .A2(G20), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT104), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT23), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1956), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n807), .A2(new_n804), .A3(new_n808), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT102), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n732), .A2(G27), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT103), .Z(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(G164), .B2(new_n732), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n443), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NOR4_X1   g420(.A1(new_n791), .A2(new_n832), .A3(new_n838), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n755), .A2(new_n756), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n727), .A2(new_n847), .ZN(G311));
  OAI21_X1  g423(.A(KEYINPUT105), .B1(new_n727), .B2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n705), .A2(new_n723), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT36), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n724), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n846), .A2(new_n756), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n755), .A4(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n849), .A2(new_n855), .ZN(G150));
  INV_X1    g431(.A(G93), .ZN(new_n857));
  INV_X1    g432(.A(G55), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n532), .A2(new_n857), .B1(new_n534), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT108), .ZN(new_n860));
  NAND2_X1  g435(.A1(G80), .A2(G543), .ZN(new_n861));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n603), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT107), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n523), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n614), .A2(G559), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT109), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n870), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n550), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n860), .A2(new_n550), .A3(new_n866), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n873), .B(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n879));
  INV_X1    g454(.A(G860), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n878), .B2(KEYINPUT39), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n869), .B1(new_n879), .B2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(G160), .B(G162), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n634), .B(new_n883), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n477), .A2(G142), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n484), .A2(G130), .ZN(new_n887));
  OR2_X1    g462(.A1(G106), .A2(G2105), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n888), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n502), .B1(new_n492), .B2(new_n494), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n783), .B2(new_n784), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n781), .A2(new_n782), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n495), .A2(new_n503), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT99), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n894), .A2(new_n900), .A3(new_n743), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n743), .B1(new_n894), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n892), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n783), .A2(new_n784), .A3(new_n893), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n742), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n894), .A2(new_n900), .A3(new_n743), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(KEYINPUT100), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n765), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n765), .A3(new_n907), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT110), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI211_X1 g487(.A(KEYINPUT110), .B(new_n765), .C1(new_n903), .C2(new_n908), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n891), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n712), .B(new_n637), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n901), .A2(new_n902), .A3(new_n892), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT100), .B1(new_n906), .B2(new_n907), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n916), .B(new_n764), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n890), .C1(new_n909), .C2(new_n911), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n915), .B1(new_n914), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n885), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n915), .ZN(new_n924));
  INV_X1    g499(.A(new_n920), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n764), .B1(new_n917), .B2(new_n918), .ZN(new_n926));
  INV_X1    g501(.A(new_n911), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n890), .B1(new_n928), .B2(new_n919), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n924), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n884), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n923), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g510(.A1(G299), .A2(new_n610), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT78), .B1(new_n572), .B2(new_n573), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n576), .A2(new_n575), .A3(new_n577), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n937), .A2(new_n938), .B1(G91), .B2(new_n520), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n607), .B1(new_n939), .B2(new_n563), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT41), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT41), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n936), .B2(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n614), .A2(new_n623), .A3(new_n877), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n877), .B1(new_n614), .B2(new_n623), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n948), .ZN(new_n950));
  INV_X1    g525(.A(new_n941), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n954));
  XNOR2_X1  g529(.A(G290), .B(G305), .ZN(new_n955));
  XOR2_X1   g530(.A(G166), .B(G288), .Z(new_n956));
  XNOR2_X1  g531(.A(new_n955), .B(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n949), .A2(new_n952), .A3(new_n959), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n954), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n958), .B1(new_n954), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g537(.A(G868), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n867), .A2(new_n598), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(G295));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n964), .ZN(G331));
  NAND3_X1  g541(.A1(new_n875), .A2(G301), .A3(new_n876), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G301), .B1(new_n875), .B2(new_n876), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n968), .A2(new_n969), .A3(G286), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n877), .A2(G171), .ZN(new_n971));
  AOI21_X1  g546(.A(G168), .B1(new_n971), .B2(new_n967), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n941), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(G286), .B1(new_n968), .B2(new_n969), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(G168), .A3(new_n967), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n942), .A3(new_n975), .A4(new_n944), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n976), .A3(new_n957), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n933), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n957), .B1(new_n973), .B2(new_n976), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n973), .A2(new_n976), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT112), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n973), .A2(new_n976), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n958), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n978), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(KEYINPUT44), .B(new_n980), .C1(new_n987), .C2(KEYINPUT43), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n985), .B2(new_n986), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n978), .A2(KEYINPUT43), .A3(new_n979), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n993));
  OAI21_X1  g568(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(G397));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n476), .A2(new_n995), .A3(new_n481), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n893), .B2(G1384), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1996), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1001), .A2(new_n785), .A3(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT113), .Z(new_n1004));
  INV_X1    g579(.A(G2067), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n742), .B(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n786), .B2(G1996), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n712), .B(new_n714), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n1001), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(G290), .B(G1986), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1000), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n898), .A2(KEYINPUT114), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n893), .B2(G1384), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n898), .A2(KEYINPUT68), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n893), .A2(new_n496), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1018), .B(new_n996), .C1(new_n1021), .C2(new_n1017), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n998), .A2(G1384), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n898), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n996), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1013), .B1(new_n504), .B2(new_n505), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(new_n998), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1022), .A2(G2090), .B1(new_n1027), .B2(G1971), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1028), .A2(G8), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G166), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(KEYINPUT115), .B2(KEYINPUT55), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT63), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1028), .A2(G8), .A3(new_n1034), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g612(.A(G1981), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n591), .A2(new_n592), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n591), .B2(new_n592), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1041), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1014), .A2(new_n996), .A3(new_n1016), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .A4(G8), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n583), .A2(new_n588), .A3(G1976), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1047), .A3(G8), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT116), .B(G1976), .Z(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(G288), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1045), .A2(new_n1051), .A3(G8), .A4(new_n1047), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1046), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1036), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1035), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G286), .A2(new_n1030), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1023), .B1(new_n504), .B2(new_n505), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n996), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT45), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1057), .B(new_n804), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1062), .A2(new_n828), .A3(new_n996), .A4(new_n1018), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT114), .B1(new_n898), .B2(new_n1013), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n893), .A2(new_n1015), .A3(G1384), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n998), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n996), .A3(new_n1058), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1057), .B1(new_n1068), .B2(new_n804), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1056), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT118), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(new_n1056), .C1(new_n1064), .C2(new_n1069), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1055), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n997), .B1(new_n1021), .B2(new_n1017), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1017), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n815), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n996), .A2(new_n1024), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1021), .B2(KEYINPUT45), .ZN(new_n1081));
  INV_X1    g656(.A(G1971), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1034), .B1(new_n1084), .B2(G8), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1054), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1074), .A2(KEYINPUT119), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT63), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT119), .B1(new_n1074), .B2(new_n1086), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1075), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1030), .B1(new_n1093), .B2(G168), .ZN(new_n1094));
  OAI21_X1  g669(.A(G286), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1068), .A2(new_n804), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT117), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1098), .A2(G168), .A3(new_n1063), .A4(new_n1061), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1099), .A2(new_n1092), .A3(G8), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT62), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(G8), .A3(new_n1095), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT51), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1094), .A2(new_n1092), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1081), .B2(G2078), .ZN(new_n1108));
  INV_X1    g683(.A(G1961), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1022), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1108), .B(new_n1110), .C1(new_n1068), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G171), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1113), .A2(new_n1054), .A3(new_n1085), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1101), .A2(new_n1106), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1045), .A2(G8), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G288), .A2(G1976), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1046), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1116), .B1(new_n1118), .B2(new_n1039), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1036), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(new_n1053), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1091), .A2(new_n1115), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1112), .A2(G171), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1107), .A2(G2078), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1080), .A2(new_n1127), .A3(new_n999), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1108), .A2(new_n1110), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(G301), .B1(new_n1129), .B2(KEYINPUT127), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(KEYINPUT127), .B2(new_n1129), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1113), .B1(G171), .B2(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1125), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1123), .A2(new_n1132), .A3(new_n1086), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n1136));
  INV_X1    g711(.A(G1956), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n996), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1137), .B1(new_n1138), .B2(new_n1077), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT57), .B1(new_n558), .B2(new_n560), .ZN(new_n1140));
  AOI22_X1  g715(.A1(G299), .A2(KEYINPUT57), .B1(new_n939), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1027), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1139), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1141), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1136), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT58), .B(G1341), .Z(new_n1147));
  NAND2_X1  g722(.A1(new_n1045), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1080), .B(new_n1002), .C1(new_n1021), .C2(KEYINPUT45), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1045), .A2(KEYINPUT122), .A3(new_n1147), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1150), .A2(new_n1151), .A3(KEYINPUT123), .A4(new_n1152), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n874), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1146), .B1(new_n1157), .B2(KEYINPUT59), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1045), .A2(G2067), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1022), .B2(new_n750), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT60), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT125), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(new_n1165), .A3(KEYINPUT60), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1164), .A2(new_n611), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1162), .A2(KEYINPUT60), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1165), .B1(new_n1162), .B2(KEYINPUT60), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1169), .B2(new_n608), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT126), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1144), .A2(KEYINPUT124), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1145), .A2(KEYINPUT121), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1136), .B1(new_n1144), .B2(KEYINPUT124), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1145), .A2(KEYINPUT121), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1167), .A2(new_n1170), .A3(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1160), .A2(new_n1172), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1144), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1162), .A2(new_n608), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT120), .Z(new_n1183));
  NAND2_X1  g758(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1181), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1135), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1012), .B1(new_n1122), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1001), .B1(new_n1006), .B2(new_n785), .ZN(new_n1188));
  OR3_X1    g763(.A1(new_n1001), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1189));
  OAI21_X1  g764(.A(KEYINPUT46), .B1(new_n1001), .B2(G1996), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT47), .Z(new_n1192));
  NOR3_X1   g767(.A1(new_n1001), .A2(G290), .A3(G1986), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT48), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1192), .B1(new_n1010), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n714), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n712), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1008), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n743), .A2(new_n1005), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1001), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1195), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1187), .A2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g777(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1204));
  OAI211_X1 g778(.A(new_n934), .B(new_n1204), .C1(new_n990), .C2(new_n991), .ZN(G225));
  INV_X1    g779(.A(G225), .ZN(G308));
endmodule


