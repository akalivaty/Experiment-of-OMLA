
module locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, 
        G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, 
        G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, 
        G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, 
        G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, 
        G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, 
        G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, 
        G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, 
        G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, 
        G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, 
        G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, 
        G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, 
        G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, 
        G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, 
        G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, 
        G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, 
        G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, 
        G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, 
        G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, G350, 
        G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, 
        G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, 
        G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, 
        G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, 
        G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, 
        G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, 
        KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, 
        KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, 
        KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, 
        KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, 
        KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, 
        KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, 
        KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, 
        KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, 
        KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, 
        KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G321, G280, G323, G331, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G284 = G321;
  assign G297 = G280;
  assign G282 = G323;
  assign G295 = G331;

  NAND2_X1 U494 ( .A1(n624), .A2(n623), .ZN(n668) );
  NOR2_X2 U495 ( .A1(n690), .A2(n681), .ZN(n682) );
  NOR2_X1 U496 ( .A1(G164), .A2(G1384), .ZN(n624) );
  NOR2_X1 U497 ( .A1(n668), .A2(n825), .ZN(n633) );
  NOR2_X1 U498 ( .A1(n861), .A2(n636), .ZN(n642) );
  NOR2_X1 U499 ( .A1(G651), .A2(G543), .ZN(n561) );
  NOR2_X1 U500 ( .A1(G651), .A2(n547), .ZN(n558) );
  NOR2_X1 U501 ( .A1(n466), .A2(n465), .ZN(G160) );
  INV_X1 U502 ( .A(G2104), .ZN(n458) );
  AND2_X1 U503 ( .A1(n458), .A2(G2105), .ZN(n768) );
  NAND2_X1 U504 ( .A1(n768), .A2(G125), .ZN(n461) );
  NOR2_X2 U505 ( .A1(G2105), .A2(n458), .ZN(n764) );
  NAND2_X1 U506 ( .A1(G101), .A2(n764), .ZN(n459) );
  XOR2_X1 U507 ( .A(KEYINPUT23), .B(n459), .Z(n460) );
  NAND2_X1 U508 ( .A1(n461), .A2(n460), .ZN(n466) );
  AND2_X1 U509 ( .A1(G2104), .A2(G2105), .ZN(n769) );
  NAND2_X1 U510 ( .A1(G113), .A2(n769), .ZN(n464) );
  NOR2_X1 U511 ( .A1(G2104), .A2(G2105), .ZN(n462) );
  XOR2_X1 U512 ( .A(KEYINPUT17), .B(n462), .Z(n765) );
  NAND2_X1 U513 ( .A1(G137), .A2(n765), .ZN(n463) );
  NAND2_X1 U514 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U515 ( .A1(G85), .A2(n561), .ZN(n468) );
  XOR2_X1 U516 ( .A(KEYINPUT0), .B(G543), .Z(n547) );
  INV_X1 U517 ( .A(G651), .ZN(n469) );
  NOR2_X1 U518 ( .A1(n547), .A2(n469), .ZN(n562) );
  NAND2_X1 U519 ( .A1(G72), .A2(n562), .ZN(n467) );
  NAND2_X1 U520 ( .A1(n468), .A2(n467), .ZN(n474) );
  NOR2_X1 U521 ( .A1(G543), .A2(n469), .ZN(n470) );
  XOR2_X1 U522 ( .A(KEYINPUT1), .B(n470), .Z(n557) );
  NAND2_X1 U523 ( .A1(G60), .A2(n557), .ZN(n472) );
  NAND2_X1 U524 ( .A1(G47), .A2(n558), .ZN(n471) );
  NAND2_X1 U525 ( .A1(n472), .A2(n471), .ZN(n473) );
  OR2_X1 U526 ( .A1(n474), .A2(n473), .ZN(G290) );
  NAND2_X1 U527 ( .A1(G64), .A2(n557), .ZN(n476) );
  NAND2_X1 U528 ( .A1(G52), .A2(n558), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n476), .A2(n475), .ZN(n481) );
  NAND2_X1 U530 ( .A1(G90), .A2(n561), .ZN(n478) );
  NAND2_X1 U531 ( .A1(G77), .A2(n562), .ZN(n477) );
  NAND2_X1 U532 ( .A1(n478), .A2(n477), .ZN(n479) );
  XOR2_X1 U533 ( .A(KEYINPUT9), .B(n479), .Z(n480) );
  NOR2_X1 U534 ( .A1(n481), .A2(n480), .ZN(G171) );
  AND2_X1 U535 ( .A1(G94), .A2(G452), .ZN(G173) );
  NAND2_X1 U536 ( .A1(G91), .A2(n561), .ZN(n483) );
  NAND2_X1 U537 ( .A1(G78), .A2(n562), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n483), .A2(n482), .ZN(n487) );
  NAND2_X1 U539 ( .A1(G65), .A2(n557), .ZN(n485) );
  NAND2_X1 U540 ( .A1(G53), .A2(n558), .ZN(n484) );
  NAND2_X1 U541 ( .A1(n485), .A2(n484), .ZN(n486) );
  NOR2_X1 U542 ( .A1(n487), .A2(n486), .ZN(n849) );
  INV_X1 U543 ( .A(n849), .ZN(G299) );
  INV_X1 U544 ( .A(G57), .ZN(G237) );
  INV_X1 U545 ( .A(G132), .ZN(G219) );
  INV_X1 U546 ( .A(G82), .ZN(G220) );
  NAND2_X1 U547 ( .A1(G7), .A2(G661), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U549 ( .A(G223), .ZN(n723) );
  NAND2_X1 U550 ( .A1(n723), .A2(G567), .ZN(n489) );
  XOR2_X1 U551 ( .A(KEYINPUT11), .B(n489), .Z(G234) );
  NAND2_X1 U552 ( .A1(G56), .A2(n557), .ZN(n490) );
  XOR2_X1 U553 ( .A(KEYINPUT14), .B(n490), .Z(n496) );
  NAND2_X1 U554 ( .A1(n561), .A2(G81), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n491), .B(KEYINPUT12), .ZN(n493) );
  NAND2_X1 U556 ( .A1(G68), .A2(n562), .ZN(n492) );
  NAND2_X1 U557 ( .A1(n493), .A2(n492), .ZN(n494) );
  XOR2_X1 U558 ( .A(KEYINPUT13), .B(n494), .Z(n495) );
  NOR2_X1 U559 ( .A1(n496), .A2(n495), .ZN(n498) );
  NAND2_X1 U560 ( .A1(n558), .A2(G43), .ZN(n497) );
  NAND2_X1 U561 ( .A1(n498), .A2(n497), .ZN(n861) );
  INV_X1 U562 ( .A(G860), .ZN(n521) );
  OR2_X1 U563 ( .A1(n861), .A2(n521), .ZN(G153) );
  INV_X1 U564 ( .A(G171), .ZN(G301) );
  NAND2_X1 U565 ( .A1(G868), .A2(G301), .ZN(n507) );
  NAND2_X1 U566 ( .A1(G66), .A2(n557), .ZN(n500) );
  NAND2_X1 U567 ( .A1(G92), .A2(n561), .ZN(n499) );
  NAND2_X1 U568 ( .A1(n500), .A2(n499), .ZN(n504) );
  NAND2_X1 U569 ( .A1(G79), .A2(n562), .ZN(n502) );
  NAND2_X1 U570 ( .A1(G54), .A2(n558), .ZN(n501) );
  NAND2_X1 U571 ( .A1(n502), .A2(n501), .ZN(n503) );
  NOR2_X1 U572 ( .A1(n504), .A2(n503), .ZN(n505) );
  XOR2_X1 U573 ( .A(KEYINPUT15), .B(n505), .Z(n846) );
  OR2_X1 U574 ( .A1(n846), .A2(G868), .ZN(n506) );
  NAND2_X1 U575 ( .A1(n507), .A2(n506), .ZN(G321) );
  NAND2_X1 U576 ( .A1(n561), .A2(G89), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n508), .B(KEYINPUT4), .ZN(n510) );
  NAND2_X1 U578 ( .A1(G76), .A2(n562), .ZN(n509) );
  NAND2_X1 U579 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n511), .B(KEYINPUT5), .ZN(n516) );
  NAND2_X1 U581 ( .A1(G63), .A2(n557), .ZN(n513) );
  NAND2_X1 U582 ( .A1(G51), .A2(n558), .ZN(n512) );
  NAND2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X1 U584 ( .A(KEYINPUT6), .B(n514), .Z(n515) );
  NAND2_X1 U585 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n517), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U587 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U588 ( .A(G868), .ZN(n518) );
  NOR2_X1 U589 ( .A1(G286), .A2(n518), .ZN(n520) );
  NOR2_X1 U590 ( .A1(G868), .A2(G299), .ZN(n519) );
  NOR2_X1 U591 ( .A1(n520), .A2(n519), .ZN(G280) );
  NAND2_X1 U592 ( .A1(n521), .A2(G559), .ZN(n522) );
  NAND2_X1 U593 ( .A1(n522), .A2(n846), .ZN(n523) );
  XNOR2_X1 U594 ( .A(n523), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U595 ( .A1(G868), .A2(n861), .ZN(n526) );
  NAND2_X1 U596 ( .A1(G868), .A2(n846), .ZN(n524) );
  NOR2_X1 U597 ( .A1(G559), .A2(n524), .ZN(n525) );
  NOR2_X1 U598 ( .A1(n526), .A2(n525), .ZN(G323) );
  NAND2_X1 U599 ( .A1(n768), .A2(G123), .ZN(n527) );
  XNOR2_X1 U600 ( .A(n527), .B(KEYINPUT18), .ZN(n529) );
  NAND2_X1 U601 ( .A1(G135), .A2(n765), .ZN(n528) );
  NAND2_X1 U602 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U603 ( .A1(G111), .A2(n769), .ZN(n531) );
  NAND2_X1 U604 ( .A1(G99), .A2(n764), .ZN(n530) );
  NAND2_X1 U605 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U606 ( .A1(n533), .A2(n532), .ZN(n796) );
  XNOR2_X1 U607 ( .A(n796), .B(G2096), .ZN(n535) );
  INV_X1 U608 ( .A(G2100), .ZN(n534) );
  NAND2_X1 U609 ( .A1(n535), .A2(n534), .ZN(G156) );
  NAND2_X1 U610 ( .A1(n846), .A2(G559), .ZN(n573) );
  XNOR2_X1 U611 ( .A(n861), .B(n573), .ZN(n536) );
  NOR2_X1 U612 ( .A1(n536), .A2(G860), .ZN(n543) );
  NAND2_X1 U613 ( .A1(G93), .A2(n561), .ZN(n538) );
  NAND2_X1 U614 ( .A1(G80), .A2(n562), .ZN(n537) );
  NAND2_X1 U615 ( .A1(n538), .A2(n537), .ZN(n542) );
  NAND2_X1 U616 ( .A1(G67), .A2(n557), .ZN(n540) );
  NAND2_X1 U617 ( .A1(G55), .A2(n558), .ZN(n539) );
  NAND2_X1 U618 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U619 ( .A1(n542), .A2(n541), .ZN(n575) );
  XNOR2_X1 U620 ( .A(n543), .B(n575), .ZN(G145) );
  NAND2_X1 U621 ( .A1(G49), .A2(n558), .ZN(n545) );
  NAND2_X1 U622 ( .A1(G74), .A2(G651), .ZN(n544) );
  NAND2_X1 U623 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U624 ( .A1(n557), .A2(n546), .ZN(n549) );
  NAND2_X1 U625 ( .A1(n547), .A2(G87), .ZN(n548) );
  NAND2_X1 U626 ( .A1(n549), .A2(n548), .ZN(G288) );
  NAND2_X1 U627 ( .A1(G61), .A2(n557), .ZN(n551) );
  NAND2_X1 U628 ( .A1(G86), .A2(n561), .ZN(n550) );
  NAND2_X1 U629 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U630 ( .A1(n562), .A2(G73), .ZN(n552) );
  XOR2_X1 U631 ( .A(KEYINPUT2), .B(n552), .Z(n553) );
  NOR2_X1 U632 ( .A1(n554), .A2(n553), .ZN(n556) );
  NAND2_X1 U633 ( .A1(n558), .A2(G48), .ZN(n555) );
  NAND2_X1 U634 ( .A1(n556), .A2(n555), .ZN(G305) );
  NAND2_X1 U635 ( .A1(G62), .A2(n557), .ZN(n560) );
  NAND2_X1 U636 ( .A1(G50), .A2(n558), .ZN(n559) );
  NAND2_X1 U637 ( .A1(n560), .A2(n559), .ZN(n566) );
  NAND2_X1 U638 ( .A1(G88), .A2(n561), .ZN(n564) );
  NAND2_X1 U639 ( .A1(G75), .A2(n562), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U641 ( .A1(n566), .A2(n565), .ZN(G166) );
  XOR2_X1 U642 ( .A(G290), .B(n861), .Z(n567) );
  XNOR2_X1 U643 ( .A(G288), .B(n567), .ZN(n570) );
  XNOR2_X1 U644 ( .A(KEYINPUT19), .B(G299), .ZN(n568) );
  XNOR2_X1 U645 ( .A(n568), .B(G305), .ZN(n569) );
  XOR2_X1 U646 ( .A(n570), .B(n569), .Z(n572) );
  XNOR2_X1 U647 ( .A(G166), .B(n575), .ZN(n571) );
  XNOR2_X1 U648 ( .A(n572), .B(n571), .ZN(n786) );
  XOR2_X1 U649 ( .A(n786), .B(n573), .Z(n574) );
  NAND2_X1 U650 ( .A1(G868), .A2(n574), .ZN(n577) );
  OR2_X1 U651 ( .A1(n575), .A2(G868), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(G331) );
  NAND2_X1 U653 ( .A1(G2078), .A2(G2084), .ZN(n578) );
  XOR2_X1 U654 ( .A(KEYINPUT20), .B(n578), .Z(n579) );
  NAND2_X1 U655 ( .A1(G2090), .A2(n579), .ZN(n580) );
  XNOR2_X1 U656 ( .A(KEYINPUT21), .B(n580), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n581), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U658 ( .A(KEYINPUT3), .B(G44), .ZN(G218) );
  NOR2_X1 U659 ( .A1(G220), .A2(G219), .ZN(n582) );
  XOR2_X1 U660 ( .A(KEYINPUT22), .B(n582), .Z(n583) );
  NOR2_X1 U661 ( .A1(G218), .A2(n583), .ZN(n584) );
  NAND2_X1 U662 ( .A1(G96), .A2(n584), .ZN(n727) );
  NAND2_X1 U663 ( .A1(n727), .A2(G2106), .ZN(n588) );
  NAND2_X1 U664 ( .A1(G69), .A2(G120), .ZN(n585) );
  NOR2_X1 U665 ( .A1(G237), .A2(n585), .ZN(n586) );
  NAND2_X1 U666 ( .A1(G108), .A2(n586), .ZN(n728) );
  NAND2_X1 U667 ( .A1(n728), .A2(G567), .ZN(n587) );
  NAND2_X1 U668 ( .A1(n588), .A2(n587), .ZN(n729) );
  NAND2_X1 U669 ( .A1(G483), .A2(G661), .ZN(n589) );
  NOR2_X1 U670 ( .A1(n729), .A2(n589), .ZN(n726) );
  NAND2_X1 U671 ( .A1(n726), .A2(G36), .ZN(G176) );
  NAND2_X1 U672 ( .A1(G126), .A2(n768), .ZN(n591) );
  NAND2_X1 U673 ( .A1(G114), .A2(n769), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U675 ( .A1(G102), .A2(n764), .ZN(n593) );
  NAND2_X1 U676 ( .A1(G138), .A2(n765), .ZN(n592) );
  NAND2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U678 ( .A1(n595), .A2(n594), .ZN(G164) );
  INV_X1 U679 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U680 ( .A(G1986), .B(G290), .ZN(n858) );
  NAND2_X1 U681 ( .A1(G160), .A2(G40), .ZN(n622) );
  NOR2_X1 U682 ( .A1(n624), .A2(n622), .ZN(n709) );
  NAND2_X1 U683 ( .A1(n858), .A2(n709), .ZN(n699) );
  XNOR2_X1 U684 ( .A(G2067), .B(KEYINPUT37), .ZN(n707) );
  NAND2_X1 U685 ( .A1(G104), .A2(n764), .ZN(n597) );
  NAND2_X1 U686 ( .A1(G140), .A2(n765), .ZN(n596) );
  NAND2_X1 U687 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U688 ( .A(KEYINPUT34), .B(n598), .ZN(n603) );
  NAND2_X1 U689 ( .A1(G128), .A2(n768), .ZN(n600) );
  NAND2_X1 U690 ( .A1(G116), .A2(n769), .ZN(n599) );
  NAND2_X1 U691 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U692 ( .A(KEYINPUT35), .B(n601), .Z(n602) );
  NOR2_X1 U693 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U694 ( .A(KEYINPUT36), .B(n604), .ZN(n776) );
  NOR2_X1 U695 ( .A1(n707), .A2(n776), .ZN(n801) );
  NAND2_X1 U696 ( .A1(n709), .A2(n801), .ZN(n705) );
  NAND2_X1 U697 ( .A1(G119), .A2(n768), .ZN(n606) );
  NAND2_X1 U698 ( .A1(G107), .A2(n769), .ZN(n605) );
  NAND2_X1 U699 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U700 ( .A1(G95), .A2(n764), .ZN(n608) );
  NAND2_X1 U701 ( .A1(G131), .A2(n765), .ZN(n607) );
  NAND2_X1 U702 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U703 ( .A1(n610), .A2(n609), .ZN(n779) );
  INV_X1 U704 ( .A(G1991), .ZN(n820) );
  NOR2_X1 U705 ( .A1(n779), .A2(n820), .ZN(n619) );
  NAND2_X1 U706 ( .A1(G129), .A2(n768), .ZN(n612) );
  NAND2_X1 U707 ( .A1(G117), .A2(n769), .ZN(n611) );
  NAND2_X1 U708 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U709 ( .A1(n764), .A2(G105), .ZN(n613) );
  XOR2_X1 U710 ( .A(KEYINPUT38), .B(n613), .Z(n614) );
  NOR2_X1 U711 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U712 ( .A1(n765), .A2(G141), .ZN(n616) );
  NAND2_X1 U713 ( .A1(n617), .A2(n616), .ZN(n761) );
  AND2_X1 U714 ( .A1(G1996), .A2(n761), .ZN(n618) );
  NOR2_X1 U715 ( .A1(n619), .A2(n618), .ZN(n803) );
  INV_X1 U716 ( .A(n709), .ZN(n620) );
  NOR2_X1 U717 ( .A1(n803), .A2(n620), .ZN(n702) );
  INV_X1 U718 ( .A(n702), .ZN(n621) );
  NAND2_X1 U719 ( .A1(n705), .A2(n621), .ZN(n697) );
  INV_X1 U720 ( .A(n622), .ZN(n623) );
  NAND2_X1 U721 ( .A1(G8), .A2(n668), .ZN(n690) );
  NOR2_X1 U722 ( .A1(G1981), .A2(G305), .ZN(n625) );
  XOR2_X1 U723 ( .A(n625), .B(KEYINPUT24), .Z(n626) );
  NOR2_X1 U724 ( .A1(n690), .A2(n626), .ZN(n695) );
  NOR2_X1 U725 ( .A1(G2084), .A2(n668), .ZN(n653) );
  NAND2_X1 U726 ( .A1(G8), .A2(n653), .ZN(n666) );
  NOR2_X1 U727 ( .A1(G1966), .A2(n690), .ZN(n664) );
  INV_X1 U728 ( .A(G1961), .ZN(n868) );
  NAND2_X1 U729 ( .A1(n668), .A2(n868), .ZN(n628) );
  INV_X1 U730 ( .A(n668), .ZN(n637) );
  XNOR2_X1 U731 ( .A(KEYINPUT25), .B(G2078), .ZN(n824) );
  NAND2_X1 U732 ( .A1(n637), .A2(n824), .ZN(n627) );
  NAND2_X1 U733 ( .A1(n628), .A2(n627), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n657), .A2(G171), .ZN(n652) );
  NAND2_X1 U735 ( .A1(n637), .A2(G2072), .ZN(n629) );
  XNOR2_X1 U736 ( .A(n629), .B(KEYINPUT27), .ZN(n631) );
  INV_X1 U737 ( .A(G1956), .ZN(n869) );
  NOR2_X1 U738 ( .A1(n869), .A2(n637), .ZN(n630) );
  NOR2_X1 U739 ( .A1(n631), .A2(n630), .ZN(n645) );
  NOR2_X1 U740 ( .A1(n645), .A2(n849), .ZN(n632) );
  XOR2_X1 U741 ( .A(n632), .B(KEYINPUT28), .Z(n649) );
  INV_X1 U742 ( .A(G1996), .ZN(n825) );
  XOR2_X1 U743 ( .A(n633), .B(KEYINPUT26), .Z(n635) );
  NAND2_X1 U744 ( .A1(n668), .A2(G1341), .ZN(n634) );
  NAND2_X1 U745 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U746 ( .A1(n846), .A2(n642), .ZN(n641) );
  NAND2_X1 U747 ( .A1(G1348), .A2(n668), .ZN(n639) );
  NAND2_X1 U748 ( .A1(G2067), .A2(n637), .ZN(n638) );
  NAND2_X1 U749 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U750 ( .A1(n641), .A2(n640), .ZN(n644) );
  OR2_X1 U751 ( .A1(n846), .A2(n642), .ZN(n643) );
  NAND2_X1 U752 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U753 ( .A1(n645), .A2(n849), .ZN(n646) );
  NAND2_X1 U754 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U755 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U756 ( .A(KEYINPUT29), .B(n650), .Z(n651) );
  NAND2_X1 U757 ( .A1(n652), .A2(n651), .ZN(n662) );
  NOR2_X1 U758 ( .A1(n664), .A2(n653), .ZN(n654) );
  NAND2_X1 U759 ( .A1(G8), .A2(n654), .ZN(n655) );
  XNOR2_X1 U760 ( .A(KEYINPUT30), .B(n655), .ZN(n656) );
  NOR2_X1 U761 ( .A1(G168), .A2(n656), .ZN(n659) );
  NOR2_X1 U762 ( .A1(G171), .A2(n657), .ZN(n658) );
  NOR2_X1 U763 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U764 ( .A(KEYINPUT31), .B(n660), .Z(n661) );
  NAND2_X1 U765 ( .A1(n662), .A2(n661), .ZN(n667) );
  INV_X1 U766 ( .A(n667), .ZN(n663) );
  NOR2_X1 U767 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U768 ( .A1(n666), .A2(n665), .ZN(n677) );
  NAND2_X1 U769 ( .A1(G286), .A2(n667), .ZN(n673) );
  NOR2_X1 U770 ( .A1(G1971), .A2(n690), .ZN(n670) );
  NOR2_X1 U771 ( .A1(G2090), .A2(n668), .ZN(n669) );
  NOR2_X1 U772 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U773 ( .A1(n671), .A2(G303), .ZN(n672) );
  NAND2_X1 U774 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U775 ( .A1(n674), .A2(G8), .ZN(n675) );
  XNOR2_X1 U776 ( .A(KEYINPUT32), .B(n675), .ZN(n676) );
  NAND2_X1 U777 ( .A1(n677), .A2(n676), .ZN(n689) );
  NOR2_X1 U778 ( .A1(G1976), .A2(G288), .ZN(n850) );
  NOR2_X1 U779 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U780 ( .A1(n850), .A2(n678), .ZN(n679) );
  NAND2_X1 U781 ( .A1(n689), .A2(n679), .ZN(n680) );
  NAND2_X1 U782 ( .A1(G1976), .A2(G288), .ZN(n851) );
  NAND2_X1 U783 ( .A1(n680), .A2(n851), .ZN(n681) );
  NOR2_X1 U784 ( .A1(KEYINPUT33), .A2(n682), .ZN(n685) );
  NAND2_X1 U785 ( .A1(n850), .A2(KEYINPUT33), .ZN(n683) );
  NOR2_X1 U786 ( .A1(n683), .A2(n690), .ZN(n684) );
  NOR2_X1 U787 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U788 ( .A(G1981), .B(G305), .Z(n843) );
  NAND2_X1 U789 ( .A1(n686), .A2(n843), .ZN(n693) );
  NOR2_X1 U790 ( .A1(G2090), .A2(G303), .ZN(n687) );
  NAND2_X1 U791 ( .A1(G8), .A2(n687), .ZN(n688) );
  NAND2_X1 U792 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U793 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U794 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U795 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U796 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U797 ( .A1(n699), .A2(n698), .ZN(n712) );
  NOR2_X1 U798 ( .A1(G1996), .A2(n761), .ZN(n805) );
  NOR2_X1 U799 ( .A1(G1986), .A2(G290), .ZN(n700) );
  AND2_X1 U800 ( .A1(n820), .A2(n779), .ZN(n797) );
  NOR2_X1 U801 ( .A1(n700), .A2(n797), .ZN(n701) );
  NOR2_X1 U802 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U803 ( .A1(n805), .A2(n703), .ZN(n704) );
  XNOR2_X1 U804 ( .A(n704), .B(KEYINPUT39), .ZN(n706) );
  NAND2_X1 U805 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n707), .A2(n776), .ZN(n809) );
  NAND2_X1 U807 ( .A1(n708), .A2(n809), .ZN(n710) );
  NAND2_X1 U808 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U810 ( .A(KEYINPUT40), .B(n713), .ZN(G329) );
  XOR2_X1 U811 ( .A(G2446), .B(G2451), .Z(n715) );
  XNOR2_X1 U812 ( .A(G2427), .B(G2443), .ZN(n714) );
  XNOR2_X1 U813 ( .A(n715), .B(n714), .ZN(n721) );
  XOR2_X1 U814 ( .A(G2430), .B(G2454), .Z(n717) );
  XNOR2_X1 U815 ( .A(G1348), .B(G1341), .ZN(n716) );
  XNOR2_X1 U816 ( .A(n717), .B(n716), .ZN(n719) );
  XOR2_X1 U817 ( .A(G2438), .B(G2435), .Z(n718) );
  XNOR2_X1 U818 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U819 ( .A(n721), .B(n720), .Z(n722) );
  NAND2_X1 U820 ( .A1(G14), .A2(n722), .ZN(n790) );
  INV_X1 U821 ( .A(n790), .ZN(G401) );
  NAND2_X1 U822 ( .A1(G2106), .A2(n723), .ZN(G217) );
  AND2_X1 U823 ( .A1(G2), .A2(G15), .ZN(n724) );
  NAND2_X1 U824 ( .A1(G661), .A2(n724), .ZN(G259) );
  NAND2_X1 U825 ( .A1(G1), .A2(G3), .ZN(n725) );
  NAND2_X1 U826 ( .A1(n726), .A2(n725), .ZN(G188) );
  INV_X1 U828 ( .A(G120), .ZN(G236) );
  INV_X1 U829 ( .A(G96), .ZN(G221) );
  INV_X1 U830 ( .A(G69), .ZN(G235) );
  NOR2_X1 U831 ( .A1(n728), .A2(n727), .ZN(G325) );
  INV_X1 U832 ( .A(G325), .ZN(G261) );
  INV_X1 U833 ( .A(n729), .ZN(G319) );
  XOR2_X1 U834 ( .A(G2100), .B(G2096), .Z(n731) );
  XNOR2_X1 U835 ( .A(G2678), .B(KEYINPUT43), .ZN(n730) );
  XNOR2_X1 U836 ( .A(n731), .B(n730), .ZN(n735) );
  XOR2_X1 U837 ( .A(KEYINPUT42), .B(G2090), .Z(n733) );
  XNOR2_X1 U838 ( .A(G2067), .B(G2072), .ZN(n732) );
  XNOR2_X1 U839 ( .A(n733), .B(n732), .ZN(n734) );
  XOR2_X1 U840 ( .A(n735), .B(n734), .Z(n737) );
  XNOR2_X1 U841 ( .A(G2078), .B(G2084), .ZN(n736) );
  XNOR2_X1 U842 ( .A(n737), .B(n736), .ZN(G227) );
  XOR2_X1 U843 ( .A(G1976), .B(G1981), .Z(n739) );
  XNOR2_X1 U844 ( .A(G1966), .B(G1956), .ZN(n738) );
  XNOR2_X1 U845 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U846 ( .A(n740), .B(G2474), .Z(n742) );
  XNOR2_X1 U847 ( .A(G1996), .B(G1991), .ZN(n741) );
  XNOR2_X1 U848 ( .A(n742), .B(n741), .ZN(n746) );
  XOR2_X1 U849 ( .A(KEYINPUT41), .B(G1971), .Z(n744) );
  XNOR2_X1 U850 ( .A(G1986), .B(G1961), .ZN(n743) );
  XNOR2_X1 U851 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U852 ( .A(n746), .B(n745), .ZN(G229) );
  NAND2_X1 U853 ( .A1(n768), .A2(G124), .ZN(n747) );
  XNOR2_X1 U854 ( .A(n747), .B(KEYINPUT44), .ZN(n749) );
  NAND2_X1 U855 ( .A1(G136), .A2(n765), .ZN(n748) );
  NAND2_X1 U856 ( .A1(n749), .A2(n748), .ZN(n753) );
  NAND2_X1 U857 ( .A1(G112), .A2(n769), .ZN(n751) );
  NAND2_X1 U858 ( .A1(G100), .A2(n764), .ZN(n750) );
  NAND2_X1 U859 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U860 ( .A1(n753), .A2(n752), .ZN(G162) );
  NAND2_X1 U861 ( .A1(G130), .A2(n768), .ZN(n755) );
  NAND2_X1 U862 ( .A1(G118), .A2(n769), .ZN(n754) );
  NAND2_X1 U863 ( .A1(n755), .A2(n754), .ZN(n760) );
  NAND2_X1 U864 ( .A1(G106), .A2(n764), .ZN(n757) );
  NAND2_X1 U865 ( .A1(G142), .A2(n765), .ZN(n756) );
  NAND2_X1 U866 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U867 ( .A(n758), .B(KEYINPUT45), .Z(n759) );
  NOR2_X1 U868 ( .A1(n760), .A2(n759), .ZN(n762) );
  XNOR2_X1 U869 ( .A(n762), .B(n761), .ZN(n763) );
  XNOR2_X1 U870 ( .A(G162), .B(n763), .ZN(n778) );
  NAND2_X1 U871 ( .A1(G103), .A2(n764), .ZN(n767) );
  NAND2_X1 U872 ( .A1(G139), .A2(n765), .ZN(n766) );
  NAND2_X1 U873 ( .A1(n767), .A2(n766), .ZN(n774) );
  NAND2_X1 U874 ( .A1(G127), .A2(n768), .ZN(n771) );
  NAND2_X1 U875 ( .A1(G115), .A2(n769), .ZN(n770) );
  NAND2_X1 U876 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U877 ( .A(KEYINPUT47), .B(n772), .Z(n773) );
  NOR2_X1 U878 ( .A1(n774), .A2(n773), .ZN(n811) );
  XOR2_X1 U879 ( .A(G160), .B(n811), .Z(n775) );
  XNOR2_X1 U880 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U881 ( .A(n778), .B(n777), .ZN(n784) );
  XOR2_X1 U882 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n781) );
  XNOR2_X1 U883 ( .A(n779), .B(n796), .ZN(n780) );
  XNOR2_X1 U884 ( .A(n781), .B(n780), .ZN(n782) );
  XOR2_X1 U885 ( .A(G164), .B(n782), .Z(n783) );
  XNOR2_X1 U886 ( .A(n784), .B(n783), .ZN(n785) );
  NOR2_X1 U887 ( .A1(G37), .A2(n785), .ZN(G395) );
  XNOR2_X1 U888 ( .A(n846), .B(G286), .ZN(n787) );
  XNOR2_X1 U889 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U890 ( .A(n788), .B(G171), .ZN(n789) );
  NOR2_X1 U891 ( .A1(G37), .A2(n789), .ZN(G397) );
  NAND2_X1 U892 ( .A1(G319), .A2(n790), .ZN(n793) );
  NOR2_X1 U893 ( .A1(G227), .A2(G229), .ZN(n791) );
  XNOR2_X1 U894 ( .A(KEYINPUT49), .B(n791), .ZN(n792) );
  NOR2_X1 U895 ( .A1(n793), .A2(n792), .ZN(n795) );
  NOR2_X1 U896 ( .A1(G395), .A2(G397), .ZN(n794) );
  NAND2_X1 U897 ( .A1(n795), .A2(n794), .ZN(G225) );
  INV_X1 U898 ( .A(G225), .ZN(G308) );
  INV_X1 U899 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U900 ( .A(G160), .B(G2084), .ZN(n799) );
  NOR2_X1 U901 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U902 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U903 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U904 ( .A1(n803), .A2(n802), .ZN(n808) );
  XOR2_X1 U905 ( .A(G2090), .B(G162), .Z(n804) );
  NOR2_X1 U906 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U907 ( .A(n806), .B(KEYINPUT51), .ZN(n807) );
  NOR2_X1 U908 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U909 ( .A1(n810), .A2(n809), .ZN(n816) );
  XOR2_X1 U910 ( .A(G2072), .B(n811), .Z(n813) );
  XOR2_X1 U911 ( .A(G164), .B(G2078), .Z(n812) );
  NOR2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U913 ( .A(KEYINPUT50), .B(n814), .Z(n815) );
  NOR2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U915 ( .A(KEYINPUT52), .B(n817), .ZN(n818) );
  INV_X1 U916 ( .A(KEYINPUT55), .ZN(n839) );
  NAND2_X1 U917 ( .A1(n818), .A2(n839), .ZN(n819) );
  NAND2_X1 U918 ( .A1(n819), .A2(G29), .ZN(n897) );
  XNOR2_X1 U919 ( .A(G2090), .B(G35), .ZN(n834) );
  XNOR2_X1 U920 ( .A(G25), .B(n820), .ZN(n821) );
  NAND2_X1 U921 ( .A1(n821), .A2(G28), .ZN(n831) );
  XNOR2_X1 U922 ( .A(G2067), .B(G26), .ZN(n823) );
  XNOR2_X1 U923 ( .A(G33), .B(G2072), .ZN(n822) );
  NOR2_X1 U924 ( .A1(n823), .A2(n822), .ZN(n829) );
  XOR2_X1 U925 ( .A(n824), .B(G27), .Z(n827) );
  XOR2_X1 U926 ( .A(n825), .B(G32), .Z(n826) );
  NOR2_X1 U927 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U928 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U929 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U930 ( .A(KEYINPUT53), .B(n832), .ZN(n833) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n837) );
  XOR2_X1 U932 ( .A(G2084), .B(KEYINPUT54), .Z(n835) );
  XNOR2_X1 U933 ( .A(G34), .B(n835), .ZN(n836) );
  NAND2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n841) );
  INV_X1 U936 ( .A(G29), .ZN(n840) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(n842) );
  NAND2_X1 U938 ( .A1(G11), .A2(n842), .ZN(n895) );
  XNOR2_X1 U939 ( .A(G16), .B(KEYINPUT56), .ZN(n867) );
  XNOR2_X1 U940 ( .A(G1966), .B(G168), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n845), .B(KEYINPUT57), .ZN(n865) );
  XOR2_X1 U943 ( .A(G1348), .B(n846), .Z(n848) );
  XOR2_X1 U944 ( .A(G171), .B(G1961), .Z(n847) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n860) );
  XNOR2_X1 U946 ( .A(n849), .B(G1956), .ZN(n856) );
  INV_X1 U947 ( .A(n850), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n852), .A2(n851), .ZN(n854) );
  XNOR2_X1 U949 ( .A(G1971), .B(G303), .ZN(n853) );
  NOR2_X1 U950 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U951 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U952 ( .A1(n858), .A2(n857), .ZN(n859) );
  NAND2_X1 U953 ( .A1(n860), .A2(n859), .ZN(n863) );
  XNOR2_X1 U954 ( .A(G1341), .B(n861), .ZN(n862) );
  NOR2_X1 U955 ( .A1(n863), .A2(n862), .ZN(n864) );
  NAND2_X1 U956 ( .A1(n865), .A2(n864), .ZN(n866) );
  NAND2_X1 U957 ( .A1(n867), .A2(n866), .ZN(n893) );
  INV_X1 U958 ( .A(G16), .ZN(n891) );
  XNOR2_X1 U959 ( .A(G5), .B(n868), .ZN(n881) );
  XNOR2_X1 U960 ( .A(G20), .B(n869), .ZN(n873) );
  XNOR2_X1 U961 ( .A(G1341), .B(G19), .ZN(n871) );
  XNOR2_X1 U962 ( .A(G1981), .B(G6), .ZN(n870) );
  NOR2_X1 U963 ( .A1(n871), .A2(n870), .ZN(n872) );
  NAND2_X1 U964 ( .A1(n873), .A2(n872), .ZN(n876) );
  XOR2_X1 U965 ( .A(KEYINPUT59), .B(G1348), .Z(n874) );
  XNOR2_X1 U966 ( .A(G4), .B(n874), .ZN(n875) );
  NOR2_X1 U967 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U968 ( .A(KEYINPUT60), .B(n877), .Z(n879) );
  XNOR2_X1 U969 ( .A(G1966), .B(G21), .ZN(n878) );
  NOR2_X1 U970 ( .A1(n879), .A2(n878), .ZN(n880) );
  NAND2_X1 U971 ( .A1(n881), .A2(n880), .ZN(n888) );
  XNOR2_X1 U972 ( .A(G1971), .B(G22), .ZN(n883) );
  XNOR2_X1 U973 ( .A(G23), .B(G1976), .ZN(n882) );
  NOR2_X1 U974 ( .A1(n883), .A2(n882), .ZN(n885) );
  XOR2_X1 U975 ( .A(G1986), .B(G24), .Z(n884) );
  NAND2_X1 U976 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U977 ( .A(KEYINPUT58), .B(n886), .ZN(n887) );
  NOR2_X1 U978 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U979 ( .A(KEYINPUT61), .B(n889), .ZN(n890) );
  NAND2_X1 U980 ( .A1(n891), .A2(n890), .ZN(n892) );
  NAND2_X1 U981 ( .A1(n893), .A2(n892), .ZN(n894) );
  NOR2_X1 U982 ( .A1(n895), .A2(n894), .ZN(n896) );
  NAND2_X1 U983 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U984 ( .A(KEYINPUT62), .B(n898), .Z(G311) );
  INV_X1 U985 ( .A(G311), .ZN(G150) );
endmodule

