//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n888, new_n889, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G141gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n203), .A2(G148gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT77), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n203), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(G148gat), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(new_n209), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n225), .A2(new_n214), .A3(new_n216), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n223), .A2(KEYINPUT80), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT80), .B1(new_n223), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n218), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT81), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT81), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n231), .B(new_n218), .C1(new_n227), .C2(new_n228), .ZN(new_n232));
  INV_X1    g031(.A(G134gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT68), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(KEYINPUT1), .ZN(new_n236));
  INV_X1    g035(.A(G120gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G113gat), .ZN(new_n238));
  INV_X1    g037(.A(G113gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G120gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n233), .ZN(new_n243));
  INV_X1    g042(.A(G127gat), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n236), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n244), .B1(new_n236), .B2(new_n243), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n232), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT82), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n226), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT80), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n226), .A3(KEYINPUT80), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n252), .A2(new_n253), .B1(new_n217), .B2(new_n212), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n243), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G127gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n243), .A3(new_n244), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n249), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n248), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n230), .A2(new_n249), .A3(new_n232), .A4(new_n247), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT83), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT83), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n260), .A2(new_n266), .A3(new_n262), .A4(new_n263), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n268));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n245), .B2(new_n246), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n256), .A2(KEYINPUT69), .A3(new_n257), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n254), .A2(new_n270), .A3(new_n271), .A4(KEYINPUT4), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n229), .B2(new_n247), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n272), .A2(new_n274), .A3(new_n261), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n230), .A2(KEYINPUT3), .A3(new_n232), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n277), .B(new_n218), .C1(new_n227), .C2(new_n228), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n247), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n268), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n267), .A3(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n229), .A2(new_n247), .A3(new_n273), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n254), .A2(new_n270), .A3(new_n271), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n273), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n268), .A2(new_n261), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n279), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G1gat), .B(G29gat), .Z(new_n288));
  XNOR2_X1  g087(.A(G57gat), .B(G85gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n290), .B(new_n291), .Z(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(KEYINPUT6), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT89), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n287), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n281), .A2(KEYINPUT89), .A3(new_n286), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n286), .A2(new_n292), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n295), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G228gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT22), .ZN(new_n313));
  OR2_X1    g112(.A1(KEYINPUT73), .A2(G197gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(KEYINPUT73), .A2(G197gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G204gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(G204gat), .A3(new_n315), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n309), .B1(new_n320), .B2(KEYINPUT74), .ZN(new_n321));
  INV_X1    g120(.A(new_n319), .ZN(new_n322));
  AOI21_X1  g121(.A(G204gat), .B1(new_n314), .B2(new_n315), .ZN(new_n323));
  OAI22_X1  g122(.A1(new_n322), .A2(new_n323), .B1(KEYINPUT22), .B2(new_n312), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n308), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n277), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n230), .A3(new_n232), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n278), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT88), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n327), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n331), .A2(new_n332), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n307), .B(new_n329), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n327), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n330), .B1(new_n320), .B2(new_n309), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n324), .A2(new_n308), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n277), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(KEYINPUT87), .A3(new_n229), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT87), .B1(new_n340), .B2(new_n229), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n306), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(KEYINPUT31), .B(G50gat), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n336), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n336), .B2(new_n344), .ZN(new_n349));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(G22gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n344), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n345), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n351), .B1(new_n355), .B2(new_n347), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT67), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT27), .B(G183gat), .ZN(new_n359));
  INV_X1    g158(.A(G190gat), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT28), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(KEYINPUT28), .ZN(new_n364));
  NOR2_X1   g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT26), .ZN(new_n366));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n365), .A2(KEYINPUT26), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n363), .A2(new_n364), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT23), .B1(new_n365), .B2(KEYINPUT65), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT65), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n374), .B(new_n375), .C1(G169gat), .C2(G176gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n369), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n379));
  AND2_X1   g178(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n367), .A2(new_n379), .B1(new_n380), .B2(G190gat), .ZN(new_n381));
  OR3_X1    g180(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n373), .A2(new_n369), .A3(new_n376), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(KEYINPUT64), .A3(G190gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n367), .ZN(new_n385));
  NAND3_X1  g184(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT64), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT25), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n382), .B1(new_n390), .B2(KEYINPUT66), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT66), .B(new_n378), .C1(new_n392), .C2(new_n377), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n372), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n270), .A2(new_n271), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT70), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n378), .B1(new_n392), .B2(new_n377), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT66), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n364), .A2(new_n371), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n401), .A2(new_n393), .B1(new_n363), .B2(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n270), .A2(new_n271), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT70), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n395), .A2(new_n396), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n397), .A2(new_n406), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT34), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT32), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n397), .A2(new_n406), .A3(new_n408), .ZN(new_n412));
  INV_X1    g211(.A(new_n407), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT33), .B1(new_n412), .B2(new_n413), .ZN(new_n415));
  XNOR2_X1  g214(.A(G15gat), .B(G43gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT71), .ZN(new_n417));
  XNOR2_X1  g216(.A(G71gat), .B(G99gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n419), .A2(KEYINPUT72), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(KEYINPUT72), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT33), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n410), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n414), .A2(new_n419), .ZN(new_n427));
  INV_X1    g226(.A(new_n415), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n410), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n424), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n357), .A2(new_n426), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  AOI22_X1  g234(.A1(new_n395), .A2(new_n330), .B1(G226gat), .B2(G233gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(G226gat), .A2(G233gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n403), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n327), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n403), .B2(KEYINPUT29), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n395), .A2(G226gat), .A3(G233gat), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n327), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n435), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n439), .B1(new_n436), .B2(new_n438), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n327), .A3(new_n442), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n435), .B(KEYINPUT75), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI22_X1  g249(.A1(new_n444), .A2(new_n445), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT76), .B1(new_n448), .B2(new_n435), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT76), .ZN(new_n453));
  INV_X1    g252(.A(new_n435), .ZN(new_n454));
  AOI211_X1 g253(.A(new_n453), .B(new_n454), .C1(new_n446), .C2(new_n447), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n451), .B1(new_n456), .B2(new_n445), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT35), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n305), .A2(new_n432), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n292), .B1(new_n281), .B2(new_n286), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n294), .B1(new_n303), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n462), .A2(new_n457), .A3(KEYINPUT86), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT86), .B1(new_n462), .B2(new_n457), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n463), .A2(new_n464), .A3(new_n432), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n460), .B1(new_n465), .B2(new_n458), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n353), .A2(new_n356), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n463), .B2(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n299), .A2(new_n304), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n448), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n446), .A2(KEYINPUT37), .A3(new_n447), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n449), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n444), .A2(new_n453), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n454), .B1(new_n446), .B2(new_n447), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT76), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n435), .B1(new_n448), .B2(new_n470), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n472), .B1(new_n479), .B2(new_n473), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n469), .A2(new_n481), .A3(new_n294), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n284), .A2(new_n279), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n262), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n260), .A2(new_n263), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n261), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(KEYINPUT39), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n261), .B1(new_n284), .B2(new_n279), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT39), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n293), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n487), .A2(new_n490), .A3(KEYINPUT40), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT40), .B1(new_n487), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n477), .A3(new_n445), .ZN(new_n494));
  INV_X1    g293(.A(new_n448), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n495), .A2(new_n449), .B1(new_n476), .B2(KEYINPUT30), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n299), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n357), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n426), .A2(new_n431), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n426), .A2(new_n431), .A3(KEYINPUT36), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n468), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n466), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G57gat), .B(G64gat), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT9), .ZN(new_n508));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT95), .ZN(new_n514));
  INV_X1    g313(.A(new_n509), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT21), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(new_n244), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT16), .ZN(new_n524));
  AOI21_X1  g323(.A(G1gat), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(KEYINPUT92), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT93), .B(G8gat), .Z(new_n528));
  OR2_X1    g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(KEYINPUT93), .B2(G8gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n512), .A2(new_n516), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(KEYINPUT21), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n522), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(new_n215), .ZN(new_n536));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n534), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G29gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n542));
  AND2_X1   g341(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n542), .B1(new_n545), .B2(G36gat), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n548));
  XNOR2_X1  g347(.A(G43gat), .B(G50gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n548), .A2(new_n549), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT91), .ZN(new_n555));
  INV_X1    g354(.A(new_n552), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT17), .ZN(new_n557));
  NAND3_X1  g356(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G99gat), .B(G106gat), .Z(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n555), .A2(new_n557), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n552), .A2(new_n568), .B1(KEYINPUT41), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n575), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n532), .A2(new_n568), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n517), .A2(new_n569), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n532), .A2(KEYINPUT10), .A3(new_n568), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n582), .A2(new_n584), .ZN(new_n590));
  INV_X1    g389(.A(new_n588), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G120gat), .B(G148gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT97), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n589), .A2(new_n592), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n540), .A2(new_n581), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT13), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n531), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n556), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n531), .A2(new_n552), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n555), .A2(new_n607), .A3(new_n557), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(new_n604), .A3(new_n609), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT18), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n604), .A4(new_n609), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G169gat), .B(G197gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n614), .A2(new_n615), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n603), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n506), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT98), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n506), .A2(new_n631), .A3(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n462), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g435(.A(new_n457), .B1(new_n630), .B2(new_n632), .ZN(new_n637));
  INV_X1    g436(.A(G8gat), .ZN(new_n638));
  OR3_X1    g437(.A1(new_n637), .A2(KEYINPUT99), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT99), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT42), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n637), .A2(new_n641), .A3(new_n642), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n639), .B(new_n640), .C1(new_n643), .C2(new_n644), .ZN(G1325gat));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646));
  INV_X1    g445(.A(new_n503), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT36), .B1(new_n426), .B2(new_n431), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n502), .A2(KEYINPUT101), .A3(new_n503), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n633), .A2(G15gat), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n500), .ZN(new_n654));
  AOI21_X1  g453(.A(G15gat), .B1(new_n633), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n655), .A2(KEYINPUT100), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(KEYINPUT100), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n633), .A2(new_n467), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  AOI21_X1  g460(.A(new_n581), .B1(new_n466), .B2(new_n505), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n540), .A2(new_n627), .A3(new_n601), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n634), .A2(new_n541), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT102), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT45), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n292), .B1(new_n287), .B2(new_n296), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n303), .B1(new_n669), .B2(new_n298), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n471), .A2(new_n454), .A3(new_n473), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT38), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n456), .A3(new_n474), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n670), .A2(new_n673), .A3(new_n295), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n498), .A2(new_n357), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n504), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n462), .A2(new_n457), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT86), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n462), .A2(new_n457), .A3(KEYINPUT86), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n357), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n305), .A2(new_n432), .A3(new_n459), .ZN(new_n683));
  INV_X1    g482(.A(new_n432), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n679), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n683), .B1(new_n685), .B2(KEYINPUT35), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n580), .C1(new_n682), .C2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n468), .A2(new_n499), .A3(new_n649), .A4(new_n650), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n581), .B1(new_n466), .B2(new_n688), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n687), .B(new_n663), .C1(new_n689), .C2(KEYINPUT44), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n462), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n667), .A2(KEYINPUT45), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n668), .A2(new_n691), .A3(new_n692), .ZN(G1328gat));
  XNOR2_X1  g492(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n664), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n457), .A2(G36gat), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n664), .A2(G36gat), .A3(new_n457), .A4(new_n694), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n690), .B2(new_n457), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G36gat), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n690), .A2(new_n701), .A3(new_n457), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n700), .B(KEYINPUT105), .C1(new_n703), .C2(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1329gat));
  NOR2_X1   g508(.A1(new_n500), .A2(G43gat), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n664), .A2(KEYINPUT106), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT106), .B1(new_n664), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n690), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(new_n652), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT107), .B1(new_n690), .B2(new_n651), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G43gat), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n690), .A2(KEYINPUT107), .A3(new_n651), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT47), .B1(new_n664), .B2(new_n711), .ZN(new_n723));
  OAI22_X1  g522(.A1(new_n718), .A2(KEYINPUT47), .B1(new_n722), .B2(new_n723), .ZN(G1330gat));
  NOR3_X1   g523(.A1(new_n664), .A2(G50gat), .A3(new_n357), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(KEYINPUT108), .B2(new_n726), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n726), .A2(KEYINPUT108), .ZN(new_n728));
  OAI21_X1  g527(.A(G50gat), .B1(new_n690), .B2(new_n357), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  NAND4_X1  g531(.A1(new_n540), .A2(new_n627), .A3(new_n581), .A4(new_n601), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n466), .B2(new_n688), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n634), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n497), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  NAND2_X1  g539(.A1(new_n734), .A2(new_n652), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n500), .A2(G71gat), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n741), .A2(G71gat), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n467), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  OR2_X1    g545(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n540), .A2(new_n626), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n602), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n747), .A2(new_n687), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n462), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n689), .A2(new_n748), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT51), .B1(new_n689), .B2(new_n748), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n634), .A2(new_n563), .A3(new_n601), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n752), .B1(new_n757), .B2(new_n758), .ZN(G1336gat));
  NAND4_X1  g558(.A1(new_n747), .A2(new_n497), .A3(new_n687), .A4(new_n750), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n457), .A2(new_n602), .A3(G92gat), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n761), .B(new_n762), .C1(new_n757), .C2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n757), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n763), .B(KEYINPUT109), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n766), .A2(new_n767), .B1(G92gat), .B2(new_n760), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n768), .B2(new_n762), .ZN(G1337gat));
  NOR2_X1   g568(.A1(new_n751), .A2(new_n651), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT110), .B(G99gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n654), .A2(new_n601), .A3(new_n771), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n770), .A2(new_n771), .B1(new_n757), .B2(new_n772), .ZN(G1338gat));
  OAI21_X1  g572(.A(G106gat), .B1(new_n751), .B2(new_n357), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n357), .A2(new_n602), .A3(G106gat), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n757), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n774), .B(new_n779), .C1(new_n757), .C2(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1339gat));
  OR2_X1    g580(.A1(new_n603), .A2(new_n626), .ZN(new_n782));
  INV_X1    g581(.A(new_n540), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n585), .A2(new_n586), .A3(new_n591), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n589), .A2(KEYINPUT54), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n591), .B1(new_n585), .B2(new_n586), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n599), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(KEYINPUT55), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n600), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT55), .B1(new_n785), .B2(new_n788), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT111), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n791), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n600), .A4(new_n789), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n626), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n608), .A2(new_n609), .A3(new_n606), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n604), .B1(new_n611), .B2(new_n609), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n621), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n625), .A2(new_n601), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n580), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n625), .A2(new_n801), .ZN(new_n804));
  AND4_X1   g603(.A1(new_n580), .A2(new_n804), .A3(new_n792), .A4(new_n795), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n783), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n782), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n684), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n808), .A2(new_n462), .A3(new_n497), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n626), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n601), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT113), .B(G120gat), .Z(new_n813));
  XNOR2_X1  g612(.A(new_n812), .B(new_n813), .ZN(G1341gat));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n540), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT68), .B(G127gat), .Z(new_n816));
  XNOR2_X1  g615(.A(new_n815), .B(new_n816), .ZN(G1342gat));
  NOR2_X1   g616(.A1(new_n462), .A2(new_n497), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n580), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n808), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n233), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n233), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(KEYINPUT56), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(KEYINPUT114), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(KEYINPUT114), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(G1343gat));
  INV_X1    g626(.A(new_n790), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n785), .A2(new_n788), .ZN(new_n829));
  XOR2_X1   g628(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n614), .A2(new_n615), .A3(new_n624), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n624), .B1(new_n614), .B2(new_n615), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n828), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n802), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n625), .A2(KEYINPUT115), .A3(new_n601), .A4(new_n801), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n581), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n580), .A2(new_n804), .A3(new_n792), .A4(new_n795), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n540), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n603), .A2(new_n626), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n467), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT57), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n807), .A2(new_n845), .A3(new_n467), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n651), .A2(new_n818), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n844), .A2(new_n846), .A3(new_n626), .A4(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n221), .ZN(new_n849));
  NOR2_X1   g648(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n807), .A2(new_n467), .A3(new_n847), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n627), .A2(G141gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n853), .A2(KEYINPUT118), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(KEYINPUT117), .A3(KEYINPUT58), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n848), .A2(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(KEYINPUT118), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n860), .B2(new_n859), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n858), .B1(new_n861), .B2(new_n863), .ZN(G1344gat));
  NAND3_X1  g663(.A1(new_n854), .A2(new_n205), .A3(new_n601), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT119), .Z(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n807), .A2(new_n467), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n580), .A2(new_n804), .A3(new_n828), .A4(new_n793), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n540), .B1(new_n839), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n845), .B(new_n467), .C1(new_n871), .C2(new_n842), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n601), .A3(new_n847), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n867), .B1(new_n874), .B2(G148gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n602), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(KEYINPUT59), .A3(new_n205), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n866), .B1(new_n875), .B2(new_n878), .ZN(G1345gat));
  XOR2_X1   g678(.A(KEYINPUT79), .B(G155gat), .Z(new_n880));
  NAND3_X1  g679(.A1(new_n854), .A2(new_n540), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n876), .A2(new_n783), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n880), .ZN(G1346gat));
  NOR4_X1   g682(.A1(new_n868), .A2(G162gat), .A3(new_n652), .A4(new_n819), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT120), .Z(new_n885));
  OAI21_X1  g684(.A(G162gat), .B1(new_n876), .B2(new_n581), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1347gat));
  NOR3_X1   g686(.A1(new_n808), .A2(new_n634), .A3(new_n457), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n626), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n601), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g691(.A1(new_n634), .A2(new_n457), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n807), .A2(new_n684), .A3(new_n540), .A4(new_n893), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(new_n359), .ZN(new_n895));
  INV_X1    g694(.A(G183gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT122), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT60), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n895), .B2(new_n897), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903));
  OAI22_X1  g702(.A1(KEYINPUT121), .A2(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1350gat));
  NOR2_X1   g704(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n888), .B2(new_n580), .ZN(new_n907));
  NAND2_X1  g706(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n907), .B(new_n908), .Z(G1351gat));
  AND2_X1   g708(.A1(new_n651), .A2(new_n893), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n869), .A2(new_n872), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(G197gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(new_n627), .ZN(new_n913));
  AND4_X1   g712(.A1(new_n467), .A2(new_n807), .A3(new_n651), .A4(new_n893), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n626), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n913), .A2(new_n915), .ZN(G1352gat));
  NAND3_X1  g715(.A1(new_n873), .A2(new_n601), .A3(new_n910), .ZN(new_n917));
  XOR2_X1   g716(.A(KEYINPUT123), .B(G204gat), .Z(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n602), .A2(new_n918), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n922));
  NOR2_X1   g721(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n919), .B(new_n924), .C1(new_n922), .C2(new_n921), .ZN(G1353gat));
  NAND3_X1  g724(.A1(new_n914), .A2(new_n310), .A3(new_n540), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n869), .A2(new_n540), .A3(new_n872), .A4(new_n910), .ZN(new_n927));
  AND2_X1   g726(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n928));
  OAI21_X1  g727(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n928), .B1(new_n927), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n926), .B1(new_n932), .B2(new_n933), .ZN(G1354gat));
  OAI21_X1  g733(.A(G218gat), .B1(new_n911), .B2(new_n581), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n914), .A2(new_n311), .A3(new_n580), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT126), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1355gat));
endmodule


