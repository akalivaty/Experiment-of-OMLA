//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT67), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  AND3_X1   g012(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n213), .A2(new_n216), .A3(KEYINPUT68), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT68), .B1(new_n213), .B2(new_n216), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(KEYINPUT23), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n226), .B2(KEYINPUT23), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n207), .B1(new_n219), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n221), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT65), .B1(new_n221), .B2(KEYINPUT23), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n222), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(new_n208), .A3(new_n209), .ZN(new_n234));
  NAND2_X1  g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT24), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n234), .A2(new_n237), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n231), .A2(new_n207), .A3(new_n232), .A4(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(G190gat), .B1(new_n208), .B2(KEYINPUT27), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT27), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G183gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(KEYINPUT69), .B(new_n209), .C1(new_n243), .C2(G183gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n247), .B2(KEYINPUT28), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n242), .A2(new_n249), .A3(new_n250), .A4(new_n244), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT26), .B1(new_n223), .B2(new_n225), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT26), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n220), .B1(new_n221), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n235), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n241), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n228), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n206), .B1(new_n258), .B2(KEYINPUT29), .ZN(new_n259));
  INV_X1    g058(.A(new_n206), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n228), .B2(new_n257), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n230), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n221), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n265));
  AND4_X1   g064(.A1(new_n207), .A2(new_n240), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n251), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n246), .A2(new_n250), .B1(new_n242), .B2(new_n244), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n235), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n224), .A2(G169gat), .A3(G176gat), .ZN(new_n271));
  INV_X1    g070(.A(G169gat), .ZN(new_n272));
  INV_X1    g071(.A(G176gat), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT66), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n254), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n255), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n232), .A2(new_n266), .B1(new_n269), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n213), .A2(new_n216), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n213), .A2(new_n216), .A3(KEYINPUT68), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n227), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT25), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT77), .A3(new_n260), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n259), .A2(new_n263), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G197gat), .B(G204gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT22), .ZN(new_n289));
  NAND2_X1  g088(.A1(G211gat), .A2(G218gat), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  INV_X1    g090(.A(G218gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT22), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n290), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n288), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT79), .B1(new_n285), .B2(new_n260), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n302));
  AOI211_X1 g101(.A(new_n302), .B(new_n206), .C1(new_n278), .C2(new_n284), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n259), .B(new_n298), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(KEYINPUT78), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n287), .A2(new_n306), .A3(new_n299), .ZN(new_n307));
  AOI211_X1 g106(.A(KEYINPUT80), .B(new_n205), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT80), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(KEYINPUT78), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT77), .B1(new_n285), .B2(new_n260), .ZN(new_n311));
  AOI211_X1 g110(.A(new_n262), .B(new_n206), .C1(new_n278), .C2(new_n284), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n298), .B1(new_n313), .B2(new_n259), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n307), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n205), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n202), .B1(new_n308), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n305), .A2(new_n205), .A3(new_n307), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n205), .B1(new_n305), .B2(new_n307), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(KEYINPUT30), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT39), .ZN(new_n324));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G141gat), .ZN(new_n328));
  INV_X1    g127(.A(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G148gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT81), .B1(new_n334), .B2(new_n335), .ZN(new_n338));
  INV_X1    g137(.A(G155gat), .ZN(new_n339));
  INV_X1    g138(.A(G162gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n342));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(KEYINPUT2), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n338), .A2(new_n344), .A3(new_n331), .A4(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n346), .A2(KEYINPUT82), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(KEYINPUT82), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n337), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n351), .B(new_n337), .C1(new_n347), .C2(new_n348), .ZN(new_n352));
  XNOR2_X1  g151(.A(G113gat), .B(G120gat), .ZN(new_n353));
  INV_X1    g152(.A(G134gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(G127gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n356));
  AND2_X1   g155(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n357));
  NOR4_X1   g156(.A1(new_n353), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(G127gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361));
  INV_X1    g160(.A(G113gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(G120gat), .ZN(new_n363));
  INV_X1    g162(.A(G120gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(G113gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n361), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G127gat), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT70), .B1(new_n367), .B2(G134gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT70), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n354), .A3(G127gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(G134gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n366), .A2(new_n372), .A3(KEYINPUT71), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT71), .B1(new_n366), .B2(new_n372), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n360), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n350), .A2(new_n352), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT83), .A4(new_n376), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n348), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n346), .A2(KEYINPUT82), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n382), .A2(new_n383), .B1(new_n336), .B2(new_n333), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n372), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT71), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n387), .A2(new_n373), .B1(new_n359), .B2(new_n358), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n349), .B2(new_n376), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n324), .B(new_n326), .C1(new_n381), .C2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n349), .B(new_n376), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n394), .A2(new_n326), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n392), .B1(new_n379), .B2(new_n380), .ZN(new_n396));
  OAI211_X1 g195(.A(KEYINPUT39), .B(new_n395), .C1(new_n396), .C2(new_n325), .ZN(new_n397));
  XOR2_X1   g196(.A(KEYINPUT84), .B(KEYINPUT0), .Z(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT40), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n402), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n396), .A2(KEYINPUT5), .A3(new_n325), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n394), .B2(new_n326), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n396), .B2(new_n325), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n405), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n403), .A2(new_n404), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n403), .A2(KEYINPUT87), .A3(new_n404), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n323), .A2(new_n412), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT37), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n315), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n305), .A2(KEYINPUT37), .A3(new_n307), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n205), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n315), .A2(new_n316), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT80), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n321), .A2(new_n309), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n422), .A2(KEYINPUT38), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n402), .B1(new_n407), .B2(new_n410), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n396), .A2(KEYINPUT5), .A3(new_n325), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n326), .B(new_n392), .C1(new_n379), .C2(new_n380), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n428), .B(new_n406), .C1(new_n429), .C2(new_n409), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n406), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT38), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n287), .A2(new_n298), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n259), .B(new_n299), .C1(new_n301), .C2(new_n303), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(KEYINPUT37), .A3(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n420), .A2(new_n435), .A3(new_n205), .A4(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n426), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G22gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT29), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n298), .B1(new_n352), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(G228gat), .A2(G233gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n296), .A2(KEYINPUT85), .A3(new_n288), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n294), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT85), .B1(new_n296), .B2(new_n288), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n444), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n351), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n447), .B1(new_n452), .B2(new_n349), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT3), .B1(new_n298), .B2(new_n444), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n384), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n447), .B1(new_n456), .B2(new_n445), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n443), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT31), .B(G50gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(new_n457), .A3(new_n443), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n460), .ZN(new_n463));
  INV_X1    g262(.A(new_n461), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n458), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n418), .A2(new_n440), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n432), .A2(new_n433), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n318), .A3(new_n322), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n466), .B(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n376), .B1(new_n228), .B2(new_n257), .ZN(new_n473));
  INV_X1    g272(.A(G227gat), .ZN(new_n474));
  INV_X1    g273(.A(G233gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n278), .A2(new_n388), .A3(new_n284), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n479), .B(KEYINPUT34), .Z(new_n480));
  INV_X1    g279(.A(KEYINPUT74), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G43gat), .ZN(new_n482));
  INV_X1    g281(.A(G99gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT73), .B(G71gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n477), .B1(new_n473), .B2(new_n478), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(KEYINPUT33), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT32), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n481), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n228), .A2(new_n376), .A3(new_n257), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n388), .B1(new_n278), .B2(new_n284), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n476), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT32), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT33), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT74), .A4(new_n486), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT75), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n486), .A2(KEYINPUT33), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n490), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n494), .A2(KEYINPUT32), .A3(new_n501), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT75), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n480), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n499), .A2(new_n505), .A3(new_n480), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(KEYINPUT76), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n509), .A2(KEYINPUT76), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n507), .B(new_n508), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n499), .A2(new_n505), .A3(new_n480), .ZN(new_n513));
  OAI22_X1  g312(.A1(new_n513), .A2(new_n506), .B1(KEYINPUT76), .B2(new_n509), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n470), .A2(new_n472), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n468), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n513), .A2(new_n506), .A3(new_n466), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n517), .A2(new_n469), .A3(new_n318), .A4(new_n322), .ZN(new_n518));
  AND2_X1   g317(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n519));
  NOR2_X1   g318(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n319), .B1(new_n423), .B2(new_n202), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n424), .A2(new_n425), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(new_n202), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n525), .A2(new_n469), .A3(new_n519), .A4(new_n517), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n516), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n516), .A2(new_n527), .A3(KEYINPUT89), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT94), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G1gat), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n536), .A2(KEYINPUT16), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n533), .B(G8gat), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n536), .A2(new_n537), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(G8gat), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n533), .A2(G8gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n536), .A2(KEYINPUT16), .A3(new_n537), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G43gat), .B(G50gat), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G29gat), .ZN(new_n551));
  INV_X1    g350(.A(G36gat), .ZN(new_n552));
  OR3_X1    g351(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT91), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OAI221_X1 g355(.A(new_n550), .B1(new_n551), .B2(new_n552), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(KEYINPUT90), .A3(new_n555), .ZN(new_n558));
  OAI221_X1 g357(.A(new_n558), .B1(KEYINPUT90), .B2(new_n553), .C1(new_n551), .C2(new_n552), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n548), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n546), .B(new_n563), .C1(new_n564), .C2(new_n561), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n540), .A2(new_n561), .A3(new_n545), .ZN(new_n566));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT18), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n567), .B(KEYINPUT13), .Z(new_n571));
  INV_X1    g370(.A(new_n566), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n561), .B1(new_n540), .B2(new_n545), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n565), .A2(KEYINPUT18), .A3(new_n566), .A4(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G113gat), .B(G141gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G197gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT11), .B(G169gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT12), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n570), .A2(new_n574), .A3(new_n575), .A4(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G127gat), .B(G155gat), .Z(new_n586));
  XOR2_X1   g385(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n587));
  OR2_X1    g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT96), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n592), .A2(KEYINPUT9), .ZN(new_n593));
  XOR2_X1   g392(.A(G57gat), .B(G64gat), .Z(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n592), .A2(KEYINPUT95), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(KEYINPUT95), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n588), .A4(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT21), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n546), .A2(new_n208), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n208), .B1(new_n546), .B2(new_n601), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n587), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n546), .A2(new_n601), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(G183gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n587), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n602), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n600), .A2(KEYINPUT21), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n605), .B2(new_n609), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n586), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n605), .A2(new_n609), .ZN(new_n615));
  INV_X1    g414(.A(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n586), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT99), .B(G211gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT100), .ZN(new_n622));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n614), .A2(new_n619), .A3(new_n626), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G99gat), .A2(G106gat), .ZN(new_n631));
  INV_X1    g430(.A(G85gat), .ZN(new_n632));
  INV_X1    g431(.A(G92gat), .ZN(new_n633));
  AOI22_X1  g432(.A1(KEYINPUT8), .A2(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT102), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT101), .B(KEYINPUT7), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n632), .A2(new_n633), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G99gat), .B(G106gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT103), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(new_n635), .A3(new_n638), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n563), .B(new_n645), .C1(new_n564), .C2(new_n561), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n644), .ZN(new_n647));
  AND2_X1   g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n561), .A2(new_n647), .B1(KEYINPUT41), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n646), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n654));
  XNOR2_X1  g453(.A(G134gat), .B(G162gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n651), .B1(new_n646), .B2(new_n649), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n653), .B2(new_n658), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n647), .A2(new_n600), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n595), .A2(new_n599), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n642), .A3(new_n644), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G230gat), .A2(G233gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT104), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT106), .B(G120gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(G176gat), .B(G204gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(new_n672));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n662), .A2(new_n673), .A3(new_n664), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n647), .A2(new_n600), .A3(KEYINPUT10), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n667), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(KEYINPUT105), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n678), .B(new_n667), .C1(new_n674), .C2(new_n675), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n668), .B(new_n672), .C1(new_n677), .C2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n672), .ZN(new_n681));
  INV_X1    g480(.A(new_n668), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n676), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n630), .A2(new_n661), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n532), .A2(new_n585), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n469), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT107), .B(G1gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1324gat));
  NAND4_X1  g488(.A1(new_n532), .A2(new_n585), .A3(new_n323), .A4(new_n685), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  OR3_X1    g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(G8gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n691), .B1(new_n690), .B2(new_n692), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(G1325gat));
  INV_X1    g495(.A(G15gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n512), .A2(new_n514), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n686), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n507), .A2(new_n508), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n686), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n697), .B2(new_n701), .ZN(G1326gat));
  INV_X1    g501(.A(new_n472), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  INV_X1    g505(.A(new_n661), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n530), .A2(new_n531), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n522), .A2(new_n526), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n515), .B2(new_n468), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n708), .B1(new_n712), .B2(new_n707), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n628), .A2(new_n629), .ZN(new_n714));
  INV_X1    g513(.A(new_n585), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n714), .A2(new_n715), .A3(new_n684), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n710), .A2(new_n434), .A3(new_n713), .A4(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(G29gat), .A3(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n530), .A2(new_n531), .A3(new_n661), .A4(new_n716), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n551), .A3(new_n434), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n724), .A2(KEYINPUT45), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(KEYINPUT45), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n721), .B1(new_n725), .B2(new_n726), .ZN(G1328gat));
  NAND3_X1  g526(.A1(new_n723), .A2(new_n552), .A3(new_n323), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n728), .A2(KEYINPUT46), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(KEYINPUT46), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n710), .A2(new_n713), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n731), .A2(new_n323), .A3(new_n716), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n729), .B(new_n730), .C1(new_n552), .C2(new_n732), .ZN(G1329gat));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n722), .B2(new_n700), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n698), .A2(new_n734), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n710), .A2(new_n713), .A3(new_n716), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g538(.A1(new_n710), .A2(new_n466), .A3(new_n713), .A4(new_n716), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G50gat), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n722), .A2(G50gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n472), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n743), .A3(KEYINPUT48), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n710), .A2(new_n472), .A3(new_n713), .A4(new_n716), .ZN(new_n745));
  AOI22_X1  g544(.A1(G50gat), .A2(new_n745), .B1(new_n742), .B2(new_n472), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n746), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g546(.A1(new_n630), .A2(new_n661), .ZN(new_n748));
  INV_X1    g547(.A(new_n684), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n585), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n528), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n469), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(G57gat), .Z(G1332gat));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n750), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n516), .B2(new_n527), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT109), .B1(new_n757), .B2(new_n748), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n525), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n760), .B2(new_n761), .ZN(G1333gat));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n512), .B(new_n514), .C1(new_n755), .C2(new_n758), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G71gat), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n700), .B(KEYINPUT110), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n751), .A2(G71gat), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n765), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g571(.A(KEYINPUT50), .B(new_n770), .C1(new_n766), .C2(G71gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1334gat));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n703), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g575(.A1(new_n714), .A2(new_n585), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n528), .A2(new_n661), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT51), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n528), .A2(new_n780), .A3(new_n661), .A4(new_n777), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n779), .A2(new_n684), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n434), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n714), .A2(new_n585), .A3(new_n749), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n731), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(new_n632), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n783), .B1(new_n786), .B2(new_n434), .ZN(G1336gat));
  NAND4_X1  g586(.A1(new_n710), .A2(new_n323), .A3(new_n713), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G92gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n525), .A2(G92gat), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n779), .A2(new_n684), .A3(new_n781), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n794), .A3(KEYINPUT52), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n789), .B(new_n793), .C1(new_n790), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n785), .B2(new_n698), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n483), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n700), .B2(new_n800), .ZN(G1338gat));
  NOR2_X1   g600(.A1(new_n467), .A2(G106gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n782), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n710), .A2(new_n466), .A3(new_n713), .A4(new_n784), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G106gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n710), .A2(new_n472), .A3(new_n713), .A4(new_n784), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n782), .A2(new_n802), .B1(new_n808), .B2(G106gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(new_n804), .ZN(G1339gat));
  NAND3_X1  g609(.A1(new_n674), .A2(new_n667), .A3(new_n675), .ZN(new_n811));
  OAI211_X1 g610(.A(KEYINPUT54), .B(new_n811), .C1(new_n677), .C2(new_n679), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n672), .B1(new_n676), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n812), .A2(new_n814), .A3(KEYINPUT55), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n585), .A3(new_n680), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n567), .B1(new_n565), .B2(new_n566), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n572), .A2(new_n573), .A3(new_n571), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n580), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n684), .A2(new_n584), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n661), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n817), .A2(new_n680), .A3(new_n818), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n661), .A2(new_n584), .A3(new_n822), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n630), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n714), .A2(new_n715), .A3(new_n707), .A4(new_n749), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n517), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n323), .A2(new_n469), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n362), .A3(new_n585), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n703), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT112), .B1(new_n830), .B2(new_n703), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n323), .A2(new_n469), .A3(new_n700), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n585), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n841), .A2(new_n842), .A3(G113gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n841), .B2(G113gat), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n834), .B1(new_n843), .B2(new_n844), .ZN(G1340gat));
  NAND3_X1  g644(.A1(new_n833), .A2(new_n364), .A3(new_n684), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n839), .A2(new_n840), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n684), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n846), .B1(new_n849), .B2(new_n364), .ZN(G1341gat));
  NAND4_X1  g649(.A1(new_n847), .A2(KEYINPUT114), .A3(G127gat), .A4(new_n714), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n833), .A2(new_n714), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n833), .A2(new_n854), .A3(new_n714), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n367), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n839), .A2(G127gat), .A3(new_n840), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n630), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n851), .A2(new_n856), .A3(new_n859), .ZN(G1342gat));
  NAND4_X1  g659(.A1(new_n831), .A2(new_n354), .A3(new_n661), .A4(new_n832), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT56), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n861), .B(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n661), .B(new_n840), .C1(new_n837), .C2(new_n838), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G134gat), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n863), .A2(KEYINPUT116), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1343gat));
  NAND2_X1  g669(.A1(new_n830), .A2(new_n466), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n832), .A2(new_n698), .ZN(new_n872));
  NOR4_X1   g671(.A1(new_n871), .A2(G141gat), .A3(new_n715), .A4(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n830), .A2(KEYINPUT57), .A3(new_n472), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n874), .B(new_n703), .C1(new_n828), .C2(new_n829), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n872), .B1(new_n879), .B2(KEYINPUT117), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n585), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n873), .B1(new_n881), .B2(G141gat), .ZN(new_n882));
  XNOR2_X1  g681(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n882), .B(new_n884), .ZN(G1344gat));
  NOR2_X1   g684(.A1(new_n871), .A2(new_n872), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n327), .A3(new_n684), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n878), .A2(new_n880), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n749), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(KEYINPUT59), .A3(new_n327), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n871), .A2(KEYINPUT57), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n830), .A2(new_n874), .A3(new_n472), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n684), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G148gat), .B1(new_n893), .B2(new_n872), .ZN(new_n894));
  XOR2_X1   g693(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n887), .B1(new_n890), .B2(new_n896), .ZN(G1345gat));
  AOI21_X1  g696(.A(G155gat), .B1(new_n886), .B2(new_n714), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n888), .A2(new_n630), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g699(.A(G162gat), .B1(new_n886), .B2(new_n661), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n888), .A2(new_n340), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n661), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n525), .A2(new_n434), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n768), .B(new_n904), .C1(new_n837), .C2(new_n838), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n715), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n831), .A2(new_n904), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n272), .A3(new_n585), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1348gat));
  NOR2_X1   g708(.A1(new_n905), .A2(new_n273), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT120), .B1(new_n910), .B2(new_n684), .ZN(new_n911));
  AOI21_X1  g710(.A(G176gat), .B1(new_n907), .B2(new_n684), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n913));
  NOR4_X1   g712(.A1(new_n905), .A2(new_n913), .A3(new_n273), .A4(new_n749), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(G1349gat));
  OAI21_X1  g714(.A(G183gat), .B1(new_n905), .B2(new_n630), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917));
  AND4_X1   g716(.A1(new_n244), .A2(new_n831), .A3(new_n714), .A4(new_n904), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n208), .A2(KEYINPUT27), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n916), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n916), .B2(new_n920), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n209), .A3(new_n661), .ZN(new_n925));
  OAI21_X1  g724(.A(G190gat), .B1(new_n905), .B2(new_n707), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(KEYINPUT61), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n928), .B(G190gat), .C1(new_n905), .C2(new_n707), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n925), .B1(new_n927), .B2(new_n930), .ZN(G1351gat));
  XNOR2_X1  g730(.A(KEYINPUT124), .B(G197gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n904), .A2(new_n698), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n891), .A2(new_n892), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(new_n935), .B2(new_n715), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n871), .A2(new_n933), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(KEYINPUT123), .ZN(new_n938));
  INV_X1    g737(.A(new_n932), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(KEYINPUT123), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n938), .A2(new_n585), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n936), .B1(new_n943), .B2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(G204gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n937), .A2(new_n946), .A3(new_n684), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT126), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n950));
  OAI21_X1  g749(.A(G204gat), .B1(new_n893), .B2(new_n933), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(G1353gat));
  NAND4_X1  g751(.A1(new_n938), .A2(new_n291), .A3(new_n714), .A4(new_n940), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n891), .A2(new_n714), .A3(new_n892), .A4(new_n934), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n953), .B(KEYINPUT127), .C1(new_n955), .C2(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1354gat));
  NAND4_X1  g760(.A1(new_n938), .A2(new_n292), .A3(new_n661), .A4(new_n940), .ZN(new_n962));
  OAI21_X1  g761(.A(G218gat), .B1(new_n935), .B2(new_n707), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1355gat));
endmodule


