

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  OR2_X1 U324 ( .A1(n387), .A2(n386), .ZN(n388) );
  INV_X1 U325 ( .A(KEYINPUT74), .ZN(n359) );
  XNOR2_X1 U326 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U327 ( .A(n362), .B(n361), .ZN(n367) );
  XNOR2_X1 U328 ( .A(n462), .B(KEYINPUT122), .ZN(n463) );
  XNOR2_X1 U329 ( .A(n464), .B(n463), .ZN(G1350GAT) );
  XOR2_X1 U330 ( .A(G15GAT), .B(G127GAT), .Z(n452) );
  XOR2_X1 U331 ( .A(G64GAT), .B(n452), .Z(n293) );
  XOR2_X1 U332 ( .A(G1GAT), .B(G8GAT), .Z(n340) );
  XNOR2_X1 U333 ( .A(n340), .B(G71GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n299) );
  XOR2_X1 U335 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n295) );
  XNOR2_X1 U336 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n355) );
  XOR2_X1 U338 ( .A(n355), .B(KEYINPUT79), .Z(n297) );
  NAND2_X1 U339 ( .A1(G231GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U341 ( .A(n299), .B(n298), .Z(n301) );
  XNOR2_X1 U342 ( .A(G22GAT), .B(G155GAT), .ZN(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n309) );
  XOR2_X1 U344 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n303) );
  XNOR2_X1 U345 ( .A(G78GAT), .B(KEYINPUT15), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U347 ( .A(G211GAT), .B(KEYINPUT78), .Z(n305) );
  XNOR2_X1 U348 ( .A(G183GAT), .B(KEYINPUT14), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U350 ( .A(n307), .B(n306), .Z(n308) );
  XOR2_X1 U351 ( .A(n309), .B(n308), .Z(n559) );
  XOR2_X1 U352 ( .A(KEYINPUT89), .B(KEYINPUT18), .Z(n311) );
  XNOR2_X1 U353 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U355 ( .A(KEYINPUT19), .B(G183GAT), .Z(n313) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(G190GAT), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U358 ( .A(n315), .B(n314), .ZN(n448) );
  XOR2_X1 U359 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n317) );
  NAND2_X1 U360 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U361 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U362 ( .A(G92GAT), .B(G204GAT), .Z(n319) );
  XNOR2_X1 U363 ( .A(G36GAT), .B(G8GAT), .ZN(n318) );
  XNOR2_X1 U364 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U365 ( .A(n321), .B(n320), .Z(n327) );
  XOR2_X1 U366 ( .A(G176GAT), .B(G64GAT), .Z(n358) );
  XNOR2_X1 U367 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n322) );
  XNOR2_X1 U368 ( .A(n322), .B(KEYINPUT93), .ZN(n323) );
  XOR2_X1 U369 ( .A(n323), .B(KEYINPUT92), .Z(n325) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(G218GAT), .ZN(n324) );
  XNOR2_X1 U371 ( .A(n325), .B(n324), .ZN(n431) );
  XNOR2_X1 U372 ( .A(n358), .B(n431), .ZN(n326) );
  XNOR2_X1 U373 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U374 ( .A(n448), .B(n328), .Z(n529) );
  XOR2_X1 U375 ( .A(KEYINPUT30), .B(G15GAT), .Z(n330) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U378 ( .A(n331), .B(KEYINPUT67), .Z(n339) );
  XOR2_X1 U379 ( .A(G113GAT), .B(G43GAT), .Z(n333) );
  XNOR2_X1 U380 ( .A(G169GAT), .B(G50GAT), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U382 ( .A(G197GAT), .B(KEYINPUT29), .Z(n335) );
  XNOR2_X1 U383 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U385 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U386 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U387 ( .A(n341), .B(n340), .Z(n345) );
  XOR2_X1 U388 ( .A(G29GAT), .B(G36GAT), .Z(n343) );
  XNOR2_X1 U389 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n342) );
  XNOR2_X1 U390 ( .A(n343), .B(n342), .ZN(n374) );
  XOR2_X1 U391 ( .A(G141GAT), .B(G22GAT), .Z(n428) );
  XNOR2_X1 U392 ( .A(n374), .B(n428), .ZN(n344) );
  XOR2_X1 U393 ( .A(n345), .B(n344), .Z(n515) );
  INV_X1 U394 ( .A(n515), .ZN(n573) );
  XOR2_X1 U395 ( .A(G85GAT), .B(G92GAT), .Z(n371) );
  XNOR2_X1 U396 ( .A(G99GAT), .B(G120GAT), .ZN(n346) );
  XNOR2_X1 U397 ( .A(n346), .B(G71GAT), .ZN(n443) );
  XNOR2_X1 U398 ( .A(n371), .B(n443), .ZN(n347) );
  AND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  NAND2_X1 U400 ( .A1(n347), .A2(n348), .ZN(n352) );
  INV_X1 U401 ( .A(n347), .ZN(n350) );
  INV_X1 U402 ( .A(n348), .ZN(n349) );
  NAND2_X1 U403 ( .A1(n350), .A2(n349), .ZN(n351) );
  NAND2_X1 U404 ( .A1(n352), .A2(n351), .ZN(n354) );
  INV_X1 U405 ( .A(KEYINPUT31), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n357) );
  XNOR2_X1 U407 ( .A(n355), .B(KEYINPUT33), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n362) );
  XNOR2_X1 U409 ( .A(KEYINPUT32), .B(n358), .ZN(n360) );
  XOR2_X1 U410 ( .A(KEYINPUT72), .B(G204GAT), .Z(n364) );
  XNOR2_X1 U411 ( .A(KEYINPUT73), .B(G78GAT), .ZN(n363) );
  XNOR2_X1 U412 ( .A(n364), .B(n363), .ZN(n366) );
  XOR2_X1 U413 ( .A(G148GAT), .B(G106GAT), .Z(n365) );
  XOR2_X1 U414 ( .A(n366), .B(n365), .Z(n440) );
  XOR2_X1 U415 ( .A(n367), .B(n440), .Z(n392) );
  XNOR2_X1 U416 ( .A(n392), .B(KEYINPUT41), .ZN(n555) );
  NOR2_X1 U417 ( .A1(n573), .A2(n555), .ZN(n368) );
  XNOR2_X1 U418 ( .A(n368), .B(KEYINPUT46), .ZN(n387) );
  XOR2_X1 U419 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n370) );
  XNOR2_X1 U420 ( .A(G99GAT), .B(G106GAT), .ZN(n369) );
  XOR2_X1 U421 ( .A(n370), .B(n369), .Z(n385) );
  XOR2_X1 U422 ( .A(G50GAT), .B(G162GAT), .Z(n427) );
  XOR2_X1 U423 ( .A(G218GAT), .B(n427), .Z(n373) );
  XNOR2_X1 U424 ( .A(G190GAT), .B(n371), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U426 ( .A(KEYINPUT76), .B(n374), .Z(n376) );
  NAND2_X1 U427 ( .A1(G232GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U429 ( .A(n378), .B(n377), .Z(n383) );
  XOR2_X1 U430 ( .A(G43GAT), .B(G134GAT), .Z(n444) );
  XOR2_X1 U431 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n380) );
  XNOR2_X1 U432 ( .A(KEYINPUT77), .B(KEYINPUT11), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n444), .B(n381), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n385), .B(n384), .ZN(n567) );
  NAND2_X1 U437 ( .A1(n559), .A2(n567), .ZN(n386) );
  XNOR2_X1 U438 ( .A(n388), .B(KEYINPUT47), .ZN(n395) );
  XNOR2_X1 U439 ( .A(KEYINPUT36), .B(n567), .ZN(n584) );
  NOR2_X1 U440 ( .A1(n559), .A2(n584), .ZN(n390) );
  XNOR2_X1 U441 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n389) );
  XNOR2_X1 U442 ( .A(n390), .B(n389), .ZN(n391) );
  NAND2_X1 U443 ( .A1(n573), .A2(n391), .ZN(n393) );
  NOR2_X1 U444 ( .A1(n393), .A2(n392), .ZN(n394) );
  NOR2_X1 U445 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U446 ( .A(n396), .B(KEYINPUT48), .ZN(n537) );
  NOR2_X1 U447 ( .A1(n529), .A2(n537), .ZN(n398) );
  XNOR2_X1 U448 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n397) );
  XNOR2_X1 U449 ( .A(n398), .B(n397), .ZN(n425) );
  XOR2_X1 U450 ( .A(KEYINPUT96), .B(KEYINPUT1), .Z(n400) );
  XNOR2_X1 U451 ( .A(G127GAT), .B(G57GAT), .ZN(n399) );
  XNOR2_X1 U452 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U453 ( .A(KEYINPUT95), .B(KEYINPUT4), .Z(n402) );
  XNOR2_X1 U454 ( .A(KEYINPUT77), .B(G148GAT), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n404), .B(n403), .ZN(n418) );
  XOR2_X1 U457 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n406) );
  XNOR2_X1 U458 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n406), .B(n405), .ZN(n416) );
  XOR2_X1 U460 ( .A(G155GAT), .B(KEYINPUT94), .Z(n408) );
  XNOR2_X1 U461 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n432) );
  XOR2_X1 U463 ( .A(G1GAT), .B(n432), .Z(n410) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U466 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n412) );
  XNOR2_X1 U467 ( .A(G141GAT), .B(G120GAT), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U469 ( .A(n414), .B(n413), .Z(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U472 ( .A(G134GAT), .B(n419), .ZN(n424) );
  XOR2_X1 U473 ( .A(G162GAT), .B(G85GAT), .Z(n422) );
  XNOR2_X1 U474 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n420), .B(KEYINPUT81), .ZN(n456) );
  XNOR2_X1 U476 ( .A(G29GAT), .B(n456), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U478 ( .A(n424), .B(n423), .Z(n502) );
  INV_X1 U479 ( .A(n502), .ZN(n526) );
  NAND2_X1 U480 ( .A1(n425), .A2(n526), .ZN(n426) );
  XOR2_X1 U481 ( .A(KEYINPUT64), .B(n426), .Z(n572) );
  XOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n430) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n436) );
  XOR2_X1 U485 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n434) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U488 ( .A(n436), .B(n435), .Z(n438) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n478) );
  NAND2_X1 U492 ( .A1(n572), .A2(n478), .ZN(n442) );
  XOR2_X1 U493 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n461) );
  XOR2_X1 U495 ( .A(n443), .B(n444), .Z(n446) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n448), .B(n447), .ZN(n460) );
  XOR2_X1 U499 ( .A(KEYINPUT87), .B(KEYINPUT83), .Z(n450) );
  XNOR2_X1 U500 ( .A(KEYINPUT86), .B(KEYINPUT82), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U502 ( .A(n451), .B(KEYINPUT20), .Z(n454) );
  XNOR2_X1 U503 ( .A(n452), .B(G176GAT), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U505 ( .A(n455), .B(KEYINPUT84), .Z(n458) );
  XNOR2_X1 U506 ( .A(n456), .B(KEYINPUT85), .ZN(n457) );
  XNOR2_X1 U507 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X2 U508 ( .A(n460), .B(n459), .Z(n531) );
  INV_X1 U509 ( .A(n531), .ZN(n538) );
  NAND2_X1 U510 ( .A1(n461), .A2(n538), .ZN(n568) );
  NOR2_X1 U511 ( .A1(n559), .A2(n568), .ZN(n464) );
  INV_X1 U512 ( .A(G183GAT), .ZN(n462) );
  NOR2_X1 U513 ( .A1(n555), .A2(n568), .ZN(n467) );
  XNOR2_X1 U514 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n465) );
  XNOR2_X1 U515 ( .A(n465), .B(G176GAT), .ZN(n466) );
  XNOR2_X1 U516 ( .A(n467), .B(n466), .ZN(G1349GAT) );
  XOR2_X1 U517 ( .A(KEYINPUT107), .B(KEYINPUT34), .Z(n469) );
  XNOR2_X1 U518 ( .A(G1GAT), .B(KEYINPUT108), .ZN(n468) );
  XNOR2_X1 U519 ( .A(n469), .B(n468), .ZN(n490) );
  NOR2_X1 U520 ( .A1(n573), .A2(n392), .ZN(n500) );
  XOR2_X1 U521 ( .A(n531), .B(KEYINPUT90), .Z(n473) );
  XNOR2_X1 U522 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n470) );
  XOR2_X1 U523 ( .A(n470), .B(n478), .Z(n511) );
  INV_X1 U524 ( .A(n529), .ZN(n506) );
  XNOR2_X1 U525 ( .A(KEYINPUT27), .B(n506), .ZN(n475) );
  NAND2_X1 U526 ( .A1(n502), .A2(n475), .ZN(n536) );
  NOR2_X1 U527 ( .A1(n511), .A2(n536), .ZN(n471) );
  XNOR2_X1 U528 ( .A(KEYINPUT103), .B(n471), .ZN(n472) );
  NOR2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n486) );
  NOR2_X1 U530 ( .A1(n478), .A2(n538), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(KEYINPUT26), .ZN(n571) );
  NAND2_X1 U532 ( .A1(n475), .A2(n571), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(KEYINPUT104), .ZN(n482) );
  NOR2_X1 U534 ( .A1(n531), .A2(n529), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(KEYINPUT105), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT25), .B(n480), .Z(n481) );
  NAND2_X1 U538 ( .A1(n482), .A2(n481), .ZN(n483) );
  NAND2_X1 U539 ( .A1(n483), .A2(n526), .ZN(n484) );
  XOR2_X1 U540 ( .A(KEYINPUT106), .B(n484), .Z(n485) );
  NOR2_X1 U541 ( .A1(n486), .A2(n485), .ZN(n497) );
  INV_X1 U542 ( .A(n559), .ZN(n579) );
  NAND2_X1 U543 ( .A1(n567), .A2(n579), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT16), .B(n487), .ZN(n488) );
  NOR2_X1 U545 ( .A1(n497), .A2(n488), .ZN(n516) );
  NAND2_X1 U546 ( .A1(n500), .A2(n516), .ZN(n495) );
  NOR2_X1 U547 ( .A1(n526), .A2(n495), .ZN(n489) );
  XOR2_X1 U548 ( .A(n490), .B(n489), .Z(G1324GAT) );
  NOR2_X1 U549 ( .A1(n529), .A2(n495), .ZN(n492) );
  XNOR2_X1 U550 ( .A(G8GAT), .B(KEYINPUT109), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  NOR2_X1 U552 ( .A1(n531), .A2(n495), .ZN(n494) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  INV_X1 U555 ( .A(n511), .ZN(n540) );
  NOR2_X1 U556 ( .A1(n540), .A2(n495), .ZN(n496) );
  XOR2_X1 U557 ( .A(G22GAT), .B(n496), .Z(G1327GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT110), .B(KEYINPUT39), .Z(n504) );
  NOR2_X1 U559 ( .A1(n584), .A2(n497), .ZN(n498) );
  NAND2_X1 U560 ( .A1(n559), .A2(n498), .ZN(n499) );
  XNOR2_X1 U561 ( .A(KEYINPUT37), .B(n499), .ZN(n525) );
  NAND2_X1 U562 ( .A1(n525), .A2(n500), .ZN(n501) );
  XOR2_X1 U563 ( .A(KEYINPUT38), .B(n501), .Z(n512) );
  NAND2_X1 U564 ( .A1(n502), .A2(n512), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(n505), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n506), .A2(n512), .ZN(n507) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(n507), .ZN(G1329GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n509) );
  NAND2_X1 U570 ( .A1(n512), .A2(n538), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n510), .ZN(G1330GAT) );
  NAND2_X1 U573 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n513), .B(KEYINPUT112), .ZN(n514) );
  XNOR2_X1 U575 ( .A(G50GAT), .B(n514), .ZN(G1331GAT) );
  NOR2_X1 U576 ( .A1(n515), .A2(n555), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n524), .A2(n516), .ZN(n521) );
  NOR2_X1 U578 ( .A1(n526), .A2(n521), .ZN(n517) );
  XOR2_X1 U579 ( .A(G57GAT), .B(n517), .Z(n518) );
  XNOR2_X1 U580 ( .A(KEYINPUT42), .B(n518), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n529), .A2(n521), .ZN(n519) );
  XOR2_X1 U582 ( .A(G64GAT), .B(n519), .Z(G1333GAT) );
  NOR2_X1 U583 ( .A1(n531), .A2(n521), .ZN(n520) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n540), .A2(n521), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n533) );
  NOR2_X1 U589 ( .A1(n526), .A2(n533), .ZN(n528) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(G1336GAT) );
  NOR2_X1 U592 ( .A1(n529), .A2(n533), .ZN(n530) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n530), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n531), .A2(n533), .ZN(n532) );
  XOR2_X1 U595 ( .A(G99GAT), .B(n532), .Z(G1338GAT) );
  NOR2_X1 U596 ( .A1(n540), .A2(n533), .ZN(n534) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(n534), .Z(n535) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n553) );
  NAND2_X1 U600 ( .A1(n553), .A2(n538), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n539), .B(KEYINPUT115), .ZN(n541) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT116), .B(n542), .ZN(n550) );
  NOR2_X1 U604 ( .A1(n573), .A2(n550), .ZN(n543) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n543), .Z(G1340GAT) );
  NOR2_X1 U606 ( .A1(n550), .A2(n555), .ZN(n545) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n547) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n549) );
  NOR2_X1 U612 ( .A1(n559), .A2(n550), .ZN(n548) );
  XOR2_X1 U613 ( .A(n549), .B(n548), .Z(G1342GAT) );
  XNOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n552) );
  NOR2_X1 U615 ( .A1(n567), .A2(n550), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n553), .A2(n571), .ZN(n562) );
  NOR2_X1 U618 ( .A1(n573), .A2(n562), .ZN(n554) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  NOR2_X1 U620 ( .A1(n555), .A2(n562), .ZN(n557) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n559), .A2(n562), .ZN(n561) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n567), .A2(n562), .ZN(n563) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NOR2_X1 U629 ( .A1(n573), .A2(n568), .ZN(n564) );
  XOR2_X1 U630 ( .A(G169GAT), .B(n564), .Z(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n566) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(n570), .B(n569), .Z(G1351GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n583) );
  NOR2_X1 U637 ( .A1(n573), .A2(n583), .ZN(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  INV_X1 U642 ( .A(n583), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n580), .A2(n392), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  XOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT125), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G218GAT), .B(n587), .Z(G1355GAT) );
endmodule

