//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT65), .B(G238), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(new_n214), .A2(G68), .B1(G77), .B2(G244), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n215), .B(new_n216), .C1(new_n207), .C2(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR4_X1   g0024(.A1(new_n218), .A2(new_n219), .A3(new_n221), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G87), .A2(G250), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n212), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  INV_X1    g0028(.A(new_n212), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  INV_X1    g0032(.A(new_n203), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n234), .A2(new_n211), .A3(new_n235), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n228), .A2(new_n232), .A3(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  AOI21_X1  g0053(.A(new_n211), .B1(new_n201), .B2(new_n203), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n254), .B1(G150), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n211), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT8), .A2(G58), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT70), .A2(G58), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT70), .A2(G58), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n258), .B1(new_n261), .B2(KEYINPUT8), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n256), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n235), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n264), .A2(new_n266), .B1(new_n222), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n210), .A2(G20), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT71), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n267), .A2(new_n235), .A3(new_n265), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G50), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT9), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n269), .A2(new_n277), .A3(new_n274), .ZN(new_n278));
  AND2_X1   g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G223), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G1698), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G222), .B2(G1698), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(G77), .B2(new_n285), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT67), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G45), .ZN(new_n291));
  AOI21_X1  g0091(.A(G41), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT68), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n210), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n294), .B1(new_n300), .B2(new_n235), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n279), .A2(KEYINPUT68), .A3(new_n280), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G226), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n287), .A2(new_n297), .A3(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n305), .A2(KEYINPUT69), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(KEYINPUT69), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n276), .A2(new_n278), .B1(new_n308), .B2(G190), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(G200), .A3(new_n307), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n309), .A2(KEYINPUT72), .A3(KEYINPUT10), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(G190), .ZN(new_n312));
  INV_X1    g0112(.A(new_n278), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n277), .B1(new_n269), .B2(new_n274), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n312), .B(new_n310), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n316));
  OR2_X1    g0116(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n308), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(new_n275), .C1(G169), .C2(new_n308), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n311), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT76), .ZN(new_n323));
  INV_X1    g0123(.A(G13), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(G1), .ZN(new_n325));
  INV_X1    g0125(.A(G68), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(G20), .A3(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT12), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(KEYINPUT12), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n273), .A2(G68), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n326), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n202), .B2(new_n257), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n266), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT75), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n335), .A3(new_n266), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT74), .B(KEYINPUT11), .Z(new_n337));
  AND3_X1   g0137(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n334), .B2(new_n336), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n330), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n303), .A2(G238), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n223), .A2(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G33), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G33), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G97), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(G232), .A2(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n346), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT73), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n285), .A2(KEYINPUT73), .A3(new_n352), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n297), .B(new_n343), .C1(new_n357), .C2(new_n281), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT13), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n285), .A2(new_n344), .B1(G33), .B2(G97), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT73), .B1(new_n285), .B2(new_n352), .ZN(new_n361));
  AND4_X1   g0161(.A1(KEYINPUT73), .A2(new_n346), .A3(new_n348), .A4(new_n352), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n281), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(new_n297), .A4(new_n343), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n342), .B1(new_n368), .B2(G169), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  AOI211_X1 g0170(.A(KEYINPUT14), .B(new_n370), .C1(new_n359), .C2(new_n367), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n359), .A2(G179), .A3(new_n367), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n341), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G190), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n359), .B2(new_n367), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n376), .A2(new_n340), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n323), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n367), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n363), .A2(new_n364), .B1(G238), .B2(new_n303), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n366), .B1(new_n382), .B2(new_n297), .ZN(new_n383));
  OAI21_X1  g0183(.A(G169), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT14), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n368), .A2(new_n342), .A3(G169), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n373), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n379), .B1(new_n387), .B2(new_n340), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT76), .ZN(new_n389));
  INV_X1    g0189(.A(new_n273), .ZN(new_n390));
  NOR2_X1   g0190(.A1(G13), .A2(G33), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n229), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT15), .B(G87), .ZN(new_n393));
  AOI21_X1  g0193(.A(G20), .B1(new_n393), .B2(G33), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT8), .B(G58), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n235), .B1(new_n395), .B2(new_n345), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n392), .A2(G77), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(G77), .B2(new_n267), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n346), .A2(new_n348), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n207), .ZN(new_n400));
  NOR2_X1   g0200(.A1(G232), .A2(G1698), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n213), .B2(G1698), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n364), .B(new_n400), .C1(new_n402), .C2(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n303), .A2(G244), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n297), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n370), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n405), .A2(G179), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n398), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n322), .A2(new_n380), .A3(new_n389), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT81), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT77), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n345), .B2(KEYINPUT3), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n347), .A2(KEYINPUT77), .A3(G33), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n282), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n223), .A2(G1698), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n414), .A2(new_n346), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n296), .B1(new_n420), .B2(new_n364), .ZN(new_n421));
  INV_X1    g0221(.A(G232), .ZN(new_n422));
  AOI211_X1 g0222(.A(new_n422), .B(new_n299), .C1(new_n301), .C2(new_n302), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(G200), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n281), .B1(new_n418), .B2(new_n419), .ZN(new_n426));
  NOR4_X1   g0226(.A1(new_n426), .A2(new_n423), .A3(G190), .A4(new_n296), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n410), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n421), .A2(new_n375), .A3(new_n424), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n426), .A2(new_n423), .A3(new_n296), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(KEYINPUT81), .C1(G200), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n262), .A2(new_n268), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n390), .B2(new_n262), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT16), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT78), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT7), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n285), .B2(G20), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT7), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT78), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n399), .A2(new_n441), .A3(new_n211), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n326), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n255), .A2(G159), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n203), .B1(new_n261), .B2(G68), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n211), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n435), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(KEYINPUT79), .B(new_n435), .C1(new_n443), .C2(new_n446), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n347), .A2(KEYINPUT77), .A3(G33), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT77), .B1(new_n347), .B2(G33), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n346), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(new_n439), .A3(new_n211), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n347), .A2(G33), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n412), .B2(new_n413), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT7), .B1(new_n457), .B2(G20), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n458), .A3(G68), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT70), .B(G58), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n233), .B1(new_n460), .B2(new_n326), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n461), .A2(G20), .B1(G159), .B2(new_n255), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(KEYINPUT16), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n463), .A2(new_n266), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n434), .B1(new_n451), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n432), .A2(new_n465), .A3(KEYINPUT17), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT17), .B1(new_n432), .B2(new_n465), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(G169), .B1(new_n421), .B2(new_n424), .ZN(new_n469));
  NOR4_X1   g0269(.A1(new_n426), .A2(new_n423), .A3(G179), .A4(new_n296), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT80), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n421), .A2(new_n319), .A3(new_n424), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT80), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(G169), .C2(new_n430), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n451), .A2(new_n464), .ZN(new_n476));
  INV_X1    g0276(.A(new_n434), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n478), .A3(KEYINPUT18), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT18), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n471), .A2(new_n474), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n465), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n398), .B1(G200), .B2(new_n405), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n405), .A2(new_n375), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n468), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n288), .A2(G1), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n294), .A3(G274), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n301), .A2(new_n302), .B1(new_n488), .B2(new_n490), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(G257), .ZN(new_n494));
  INV_X1    g0294(.A(G244), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G1698), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n496), .B(new_n346), .C1(new_n452), .C2(new_n453), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT84), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT84), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n457), .A2(new_n500), .A3(new_n496), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g0303(.A(G250), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(new_n415), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n505), .A2(new_n285), .B1(G33), .B2(G283), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT85), .B1(new_n507), .B2(new_n364), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT85), .ZN(new_n509));
  AOI211_X1 g0309(.A(new_n509), .B(new_n281), .C1(new_n502), .C2(new_n506), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n319), .B(new_n494), .C1(new_n508), .C2(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n511), .A2(KEYINPUT87), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n267), .A2(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n438), .A2(new_n442), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G107), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT83), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g0317(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n518));
  NAND2_X1  g0318(.A1(new_n207), .A2(G97), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g0320(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n208), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(G20), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n255), .A2(G77), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n514), .A2(KEYINPUT83), .A3(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n517), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n513), .B1(new_n528), .B2(new_n266), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n272), .B1(new_n210), .B2(G33), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G97), .ZN(new_n531));
  INV_X1    g0331(.A(new_n494), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n507), .B2(new_n364), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n529), .A2(new_n531), .B1(new_n534), .B2(new_n370), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n511), .A2(KEYINPUT87), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n512), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n507), .A2(new_n364), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(G190), .A3(new_n494), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n529), .A2(new_n531), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n494), .B1(new_n508), .B2(new_n510), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G200), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(KEYINPUT86), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT86), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n537), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G238), .A2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n495), .B2(G1698), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n457), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n364), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT88), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n301), .A2(new_n302), .ZN(new_n553));
  INV_X1    g0353(.A(new_n490), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(G250), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n551), .A2(new_n552), .A3(new_n491), .A4(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n457), .A2(new_n547), .B1(G33), .B2(G116), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n491), .B(new_n555), .C1(new_n557), .C2(new_n281), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT88), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G190), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n257), .B2(new_n206), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n563), .B(KEYINPUT89), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n326), .A2(G20), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n211), .B1(new_n350), .B2(new_n562), .ZN(new_n566));
  OR3_X1    g0366(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n457), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n266), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n393), .A2(new_n268), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n530), .A2(G87), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n561), .B(new_n573), .C1(new_n377), .C2(new_n560), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n560), .A2(new_n319), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n556), .A2(new_n559), .A3(new_n370), .ZN(new_n576));
  XOR2_X1   g0376(.A(new_n393), .B(KEYINPUT90), .Z(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n530), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n570), .A2(new_n578), .A3(new_n571), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n220), .A2(new_n415), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n217), .A2(G1698), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n457), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  XOR2_X1   g0384(.A(KEYINPUT91), .B(G303), .Z(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n399), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n281), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(KEYINPUT5), .A2(G41), .ZN(new_n588));
  NOR2_X1   g0388(.A1(KEYINPUT5), .A2(G41), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n490), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n300), .A2(new_n294), .A3(new_n235), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT68), .B1(new_n279), .B2(new_n280), .ZN(new_n592));
  OAI211_X1 g0392(.A(G270), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NOR4_X1   g0394(.A1(new_n587), .A2(new_n594), .A3(new_n319), .A4(new_n492), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n530), .A2(G116), .ZN(new_n596));
  INV_X1    g0396(.A(G116), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n325), .A2(G20), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n265), .A2(new_n235), .B1(G20), .B2(new_n597), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G33), .A2(G283), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n600), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT20), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n599), .A2(KEYINPUT20), .A3(new_n601), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n596), .B(new_n598), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n587), .A2(new_n492), .A3(new_n594), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G190), .ZN(new_n607));
  INV_X1    g0407(.A(new_n604), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(new_n377), .C2(new_n606), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n584), .A2(new_n586), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n364), .ZN(new_n611));
  INV_X1    g0411(.A(new_n492), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(new_n593), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n613), .A2(KEYINPUT21), .A3(G169), .A4(new_n604), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n604), .A2(G169), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(new_n606), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n605), .A2(new_n609), .A3(new_n614), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n285), .A2(new_n211), .A3(G87), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT22), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT23), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n211), .B2(G107), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n619), .A2(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n457), .A2(KEYINPUT22), .A3(new_n211), .A4(G87), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT24), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n624), .A2(KEYINPUT24), .A3(new_n625), .A4(new_n626), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n266), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n530), .A2(G107), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n325), .A2(G20), .A3(new_n207), .ZN(new_n633));
  XOR2_X1   g0433(.A(new_n633), .B(KEYINPUT25), .Z(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n504), .A2(new_n415), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n220), .A2(G1698), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n457), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(G33), .A2(G294), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n364), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT92), .ZN(new_n642));
  OAI211_X1 g0442(.A(G264), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n281), .B1(new_n638), .B2(new_n639), .ZN(new_n645));
  INV_X1    g0445(.A(new_n643), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT92), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI211_X1 g0447(.A(new_n319), .B(new_n492), .C1(new_n644), .C2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n370), .B1(new_n649), .B2(new_n612), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n635), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n644), .A2(new_n647), .ZN(new_n653));
  AOI21_X1  g0453(.A(G200), .B1(new_n653), .B2(new_n612), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n641), .A2(new_n375), .A3(new_n612), .A4(new_n643), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT93), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n649), .A2(KEYINPUT93), .A3(new_n375), .A4(new_n612), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n652), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n581), .A2(new_n618), .A3(new_n651), .A4(new_n660), .ZN(new_n661));
  NOR4_X1   g0461(.A1(new_n409), .A2(new_n487), .A3(new_n545), .A4(new_n661), .ZN(G372));
  INV_X1    g0462(.A(new_n321), .ZN(new_n663));
  INV_X1    g0463(.A(new_n379), .ZN(new_n664));
  INV_X1    g0464(.A(new_n408), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n468), .B(new_n664), .C1(new_n374), .C2(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n666), .A2(KEYINPUT95), .A3(new_n483), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT95), .B1(new_n666), .B2(new_n483), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n311), .A2(new_n318), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n663), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n409), .A2(new_n487), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT86), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n541), .A2(G200), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n529), .A2(new_n531), .A3(new_n539), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n540), .A2(KEYINPUT86), .A3(new_n542), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT87), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n511), .B(new_n679), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n677), .A2(new_n678), .B1(new_n680), .B2(new_n535), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n560), .A2(G190), .B1(G200), .B2(new_n558), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT94), .ZN(new_n684));
  INV_X1    g0484(.A(new_n579), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n319), .B2(new_n560), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n558), .A2(new_n370), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n682), .A2(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n617), .A2(new_n614), .A3(new_n605), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n651), .A2(new_n689), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n688), .A2(new_n660), .A3(new_n690), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n681), .A2(new_n691), .B1(new_n686), .B2(new_n687), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n574), .A2(new_n580), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT26), .B1(new_n537), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT26), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n688), .A2(new_n680), .A3(new_n695), .A4(new_n535), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n673), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n672), .A2(new_n699), .ZN(G369));
  NOR3_X1   g0500(.A1(new_n324), .A2(G1), .A3(G20), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT96), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT27), .ZN(new_n703));
  OR3_X1    g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G213), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n701), .B2(new_n703), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n702), .B1(new_n701), .B2(new_n703), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT97), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT97), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(G343), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n635), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n714), .A2(KEYINPUT98), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(KEYINPUT98), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n715), .A2(new_n651), .A3(new_n660), .A4(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n651), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n713), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n689), .ZN(new_n721));
  INV_X1    g0521(.A(new_n713), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n722), .A2(new_n608), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n721), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n689), .A2(new_n609), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(new_n725), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n717), .A2(new_n723), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n718), .A2(new_n722), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(G399));
  NAND2_X1  g0534(.A1(new_n686), .A2(new_n687), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT100), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n680), .A2(new_n581), .A3(new_n695), .A4(new_n535), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n688), .A2(new_n660), .A3(new_n690), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n736), .B(new_n737), .C1(new_n545), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n684), .A2(new_n682), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n735), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n537), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n695), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT29), .B(new_n722), .C1(new_n739), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n713), .B1(new_n692), .B2(new_n697), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n745), .B2(KEYINPUT29), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n560), .A2(new_n533), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n642), .B1(new_n641), .B2(new_n643), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n645), .A2(KEYINPUT92), .A3(new_n646), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n595), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n747), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n611), .A2(G179), .A3(new_n612), .A4(new_n593), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n647), .B2(new_n644), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n754), .A2(KEYINPUT30), .A3(new_n533), .A4(new_n560), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n541), .A2(new_n319), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n612), .B1(new_n749), .B2(new_n750), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n613), .A3(new_n558), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n752), .B(new_n755), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n713), .ZN(new_n760));
  AOI21_X1  g0560(.A(KEYINPUT31), .B1(new_n759), .B2(new_n713), .ZN(new_n761));
  OAI21_X1  g0561(.A(KEYINPUT99), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n713), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT31), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT99), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n713), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n660), .A2(new_n651), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(new_n727), .A3(new_n693), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n677), .A2(new_n678), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n770), .A2(new_n537), .A3(new_n771), .A4(new_n722), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n762), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G330), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n746), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(KEYINPUT101), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(KEYINPUT101), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n777), .A2(new_n210), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n230), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G41), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n567), .A2(G116), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n782), .A2(G1), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n234), .B2(new_n782), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n779), .A2(new_n786), .ZN(G364));
  INV_X1    g0587(.A(new_n729), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n728), .A2(G330), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n324), .A2(G20), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G45), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n782), .A2(G1), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n788), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n391), .B(KEYINPUT102), .Z(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n235), .B1(G20), .B2(new_n370), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n249), .A2(G45), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n230), .A2(new_n454), .ZN(new_n801));
  INV_X1    g0601(.A(new_n234), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n289), .A2(new_n291), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n800), .A2(new_n805), .B1(new_n597), .B2(new_n780), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n230), .A2(G355), .A3(new_n285), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n799), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n375), .A2(G200), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n319), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G97), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n211), .A2(G179), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G190), .A2(G200), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G159), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT32), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n812), .A2(new_n285), .A3(new_n817), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n211), .A2(new_n319), .A3(KEYINPUT103), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT103), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G20), .B2(G179), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n377), .A2(G190), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n813), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n825), .A2(new_n326), .B1(new_n207), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n375), .A2(new_n377), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n818), .B(new_n827), .C1(G50), .C2(new_n830), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n822), .A2(G190), .A3(G200), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(G77), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n828), .A2(new_n813), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(G87), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n815), .A2(KEYINPUT32), .A3(new_n816), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT104), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n823), .B2(new_n809), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n822), .A2(KEYINPUT104), .A3(new_n375), .A4(G200), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n837), .B1(new_n842), .B2(new_n261), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n831), .A2(new_n833), .A3(new_n836), .A4(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n830), .A2(G326), .B1(G294), .B2(new_n811), .ZN(new_n845));
  INV_X1    g0645(.A(G311), .ZN(new_n846));
  INV_X1    g0646(.A(new_n832), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT105), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n835), .A2(G303), .ZN(new_n850));
  INV_X1    g0650(.A(new_n815), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G329), .ZN(new_n852));
  XNOR2_X1  g0652(.A(KEYINPUT106), .B(KEYINPUT33), .ZN(new_n853));
  INV_X1    g0653(.A(G317), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n399), .B1(new_n825), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n842), .B2(G322), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n849), .A2(new_n850), .A3(new_n852), .A4(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G283), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n826), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n844), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n808), .B1(new_n861), .B2(new_n797), .ZN(new_n862));
  INV_X1    g0662(.A(new_n792), .ZN(new_n863));
  INV_X1    g0663(.A(new_n796), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n862), .B(new_n863), .C1(new_n728), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n793), .A2(new_n865), .ZN(G396));
  INV_X1    g0666(.A(new_n825), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G137), .A2(new_n830), .B1(new_n867), .B2(G150), .ZN(new_n868));
  XNOR2_X1  g0668(.A(KEYINPUT107), .B(G143), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n868), .B1(new_n816), .B2(new_n847), .C1(new_n841), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT34), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(G132), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n457), .B1(new_n874), .B2(new_n815), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n871), .B2(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n811), .A2(new_n261), .ZN(new_n877));
  INV_X1    g0677(.A(new_n826), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G50), .A2(new_n835), .B1(new_n878), .B2(G68), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n873), .A2(new_n876), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n842), .A2(G294), .B1(G311), .B2(new_n851), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n830), .A2(G303), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n881), .A2(new_n812), .A3(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n883), .B(new_n399), .C1(new_n597), .C2(new_n847), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n878), .A2(G87), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n885), .B1(new_n207), .B2(new_n834), .C1(new_n825), .C2(new_n859), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n880), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT108), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n888), .A2(new_n797), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n797), .A2(new_n391), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n202), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n408), .A2(new_n713), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n484), .A2(new_n485), .B1(new_n398), .B2(new_n713), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(new_n665), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n863), .B(new_n891), .C1(new_n896), .C2(new_n795), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n745), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n895), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT109), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n735), .B1(new_n545), .B2(new_n738), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n694), .A2(new_n696), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n722), .B(new_n896), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n899), .A2(KEYINPUT109), .A3(new_n895), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(new_n774), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n898), .B1(new_n908), .B2(new_n792), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(G384));
  NOR2_X1   g0710(.A1(new_n760), .A2(new_n761), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n772), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n673), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT113), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n713), .A2(new_n340), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n388), .A2(new_n915), .B1(new_n374), .B2(new_n713), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n895), .B(new_n916), .C1(new_n772), .C2(new_n911), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT112), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT37), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n478), .B1(new_n475), .B2(new_n712), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n432), .A2(new_n465), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n463), .A2(new_n266), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n449), .B2(new_n450), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n471), .B(new_n474), .C1(new_n925), .C2(new_n434), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n712), .B1(new_n925), .B2(new_n434), .ZN(new_n927));
  AND4_X1   g0727(.A1(new_n920), .A2(new_n926), .A3(new_n922), .A4(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n919), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n927), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT18), .B1(new_n475), .B2(new_n478), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n481), .A2(new_n465), .A3(new_n480), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT17), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n922), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n432), .A2(new_n465), .A3(KEYINPUT17), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n930), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n465), .B1(new_n481), .B2(new_n711), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n432), .A2(new_n465), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT37), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n926), .A2(new_n922), .A3(new_n927), .A4(new_n920), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(KEYINPUT112), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n929), .A2(new_n938), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT38), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n459), .A2(new_n462), .ZN(new_n947));
  NOR2_X1   g0747(.A1(KEYINPUT111), .A2(KEYINPUT16), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n947), .B(new_n948), .Z(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n266), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n477), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n712), .B(new_n951), .C1(new_n933), .C2(new_n937), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n481), .A2(new_n711), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n940), .B1(new_n953), .B2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n942), .B1(new_n954), .B2(new_n920), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(KEYINPUT38), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n918), .B1(new_n946), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n916), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n895), .B1(new_n772), .B2(new_n911), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n952), .A2(KEYINPUT38), .A3(new_n955), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT38), .B1(new_n952), .B2(new_n955), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n958), .B(new_n959), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n917), .A2(new_n957), .B1(new_n962), .B2(new_n918), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n914), .B(new_n963), .Z(new_n964));
  AND2_X1   g0764(.A1(new_n964), .A2(G330), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n916), .B1(new_n904), .B2(new_n893), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n961), .B2(new_n960), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n483), .A2(new_n712), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n961), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(KEYINPUT39), .A3(new_n956), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n960), .B1(new_n945), .B2(new_n944), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n971), .B1(new_n972), .B2(KEYINPUT39), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n387), .A2(new_n340), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n713), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n967), .B(new_n969), .C1(new_n973), .C2(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n744), .B(new_n673), .C1(new_n745), .C2(KEYINPUT29), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n672), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n977), .B(new_n979), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n965), .B1(KEYINPUT114), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n980), .B(KEYINPUT114), .Z(new_n982));
  OAI221_X1 g0782(.A(new_n981), .B1(new_n210), .B2(new_n790), .C1(new_n982), .C2(new_n965), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT35), .B1(new_n520), .B2(new_n523), .ZN(new_n984));
  NOR4_X1   g0784(.A1(new_n984), .A2(new_n211), .A3(new_n597), .A4(new_n235), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT110), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n520), .A2(KEYINPUT35), .A3(new_n523), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT36), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n802), .B1(new_n460), .B2(new_n326), .ZN(new_n990));
  INV_X1    g0790(.A(new_n201), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n990), .A2(new_n202), .B1(new_n326), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(G1), .A3(new_n324), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n983), .A2(new_n989), .A3(new_n993), .ZN(G367));
  NOR2_X1   g0794(.A1(new_n731), .A2(new_n545), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n529), .A2(new_n531), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n681), .B1(new_n997), .B2(new_n722), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n537), .B1(new_n998), .B2(new_n651), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT115), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(KEYINPUT115), .B(new_n537), .C1(new_n998), .C2(new_n651), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1001), .A2(new_n722), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n996), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n722), .A2(new_n684), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(new_n686), .A3(new_n687), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n741), .B2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(KEYINPUT43), .B2(new_n1007), .ZN(new_n1010));
  AOI211_X1 g0810(.A(KEYINPUT43), .B(new_n1007), .C1(new_n996), .C2(new_n1003), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n730), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT116), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n680), .A2(new_n535), .A3(new_n713), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n998), .A2(new_n1015), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1014), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1010), .A2(new_n1012), .A3(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n996), .A2(new_n1003), .B1(KEYINPUT43), .B2(new_n1007), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1018), .B1(new_n1023), .B2(new_n1011), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n791), .A2(G1), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n731), .A2(new_n733), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n1016), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT45), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1029), .A2(new_n1016), .A3(KEYINPUT45), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT44), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n1029), .B2(new_n1016), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1028), .A2(KEYINPUT44), .A3(new_n998), .A4(new_n1015), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n788), .A2(new_n723), .A3(new_n720), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n732), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n777), .A2(new_n778), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n781), .B(KEYINPUT41), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1027), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1025), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n834), .A2(new_n597), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT117), .B1(new_n1048), .B2(KEYINPUT46), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G317), .B2(new_n851), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n457), .B1(new_n811), .B2(G107), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n878), .A2(G97), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1048), .A2(KEYINPUT117), .A3(KEYINPUT46), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G294), .A2(new_n867), .B1(new_n830), .B2(G311), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(KEYINPUT46), .B2(new_n1048), .C1(new_n859), .C2(new_n847), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(new_n585), .C2(new_n842), .ZN(new_n1057));
  INV_X1    g0857(.A(G137), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n811), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n285), .B1(new_n815), .B2(new_n1058), .C1(new_n1059), .C2(new_n326), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n830), .A2(new_n869), .B1(G77), .B2(new_n878), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n832), .A2(new_n991), .B1(new_n261), .B2(new_n835), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n816), .C2(new_n825), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1060), .B(new_n1063), .C1(G150), .C2(new_n842), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1057), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT47), .Z(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n797), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1007), .A2(new_n864), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n798), .B1(new_n230), .B2(new_n393), .C1(new_n245), .C2(new_n801), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1067), .A2(new_n863), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1047), .A2(new_n1070), .ZN(G387));
  INV_X1    g0871(.A(new_n778), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1042), .B1(new_n1072), .B2(new_n776), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n777), .A2(new_n778), .A3(new_n1041), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n1074), .A3(new_n781), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n720), .A2(new_n796), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT50), .B1(new_n395), .B2(G50), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1077), .A2(new_n783), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(G68), .A2(G77), .ZN(new_n1079));
  OR3_X1    g0879(.A1(new_n395), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1078), .A2(new_n288), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n801), .B1(new_n242), .B2(new_n803), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n780), .A2(new_n783), .A3(new_n399), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n780), .A2(new_n207), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n799), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(G150), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n834), .A2(new_n202), .B1(new_n815), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT118), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n454), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n1052), .C1(new_n1089), .C2(new_n1088), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT119), .Z(new_n1092));
  OAI22_X1  g0892(.A1(new_n841), .A2(new_n222), .B1(new_n326), .B2(new_n847), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n867), .A2(new_n262), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n830), .A2(G159), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n577), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n1059), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n867), .A2(G311), .B1(new_n585), .B2(new_n832), .ZN(new_n1101));
  INV_X1    g0901(.A(G322), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n829), .C1(new_n854), .C2(new_n841), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT48), .ZN(new_n1104));
  INV_X1    g0904(.A(G294), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1104), .B1(new_n859), .B2(new_n1059), .C1(new_n1105), .C2(new_n834), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT49), .Z(new_n1107));
  INV_X1    g0907(.A(G326), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n454), .B1(new_n597), .B2(new_n826), .C1(new_n1108), .C2(new_n815), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1100), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1076), .B(new_n1086), .C1(new_n1110), .C2(new_n797), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n863), .A2(new_n1111), .B1(new_n1042), .B2(new_n1026), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1075), .A2(new_n1112), .ZN(G393));
  OAI211_X1 g0913(.A(new_n1042), .B(new_n1039), .C1(new_n1072), .C2(new_n776), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1073), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1039), .A2(new_n1013), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n730), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n781), .B(new_n1114), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n998), .A2(new_n796), .A3(new_n1015), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n798), .B1(new_n206), .B2(new_n230), .C1(new_n252), .C2(new_n801), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n842), .A2(G159), .B1(G150), .B2(new_n830), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT120), .B(KEYINPUT51), .Z(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1122), .A2(new_n1124), .B1(new_n326), .B2(new_n834), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n811), .A2(G77), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n885), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n454), .B(new_n1128), .C1(new_n867), .C2(new_n991), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1126), .B(new_n1129), .C1(new_n395), .C2(new_n847), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1125), .B(new_n1130), .C1(new_n851), .C2(new_n869), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n867), .A2(new_n585), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n597), .B2(new_n1059), .C1(new_n1105), .C2(new_n847), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT121), .Z(new_n1134));
  OAI22_X1  g0934(.A1(new_n841), .A2(new_n846), .B1(new_n854), .B2(new_n829), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT52), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n826), .A2(new_n207), .B1(new_n815), .B2(new_n1102), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n285), .B(new_n1137), .C1(G283), .C2(new_n835), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n797), .B1(new_n1131), .B2(new_n1140), .ZN(new_n1141));
  AND4_X1   g0941(.A1(new_n863), .A2(new_n1120), .A3(new_n1121), .A4(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1118), .B2(new_n1026), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1119), .A2(new_n1143), .ZN(G390));
  AOI21_X1  g0944(.A(KEYINPUT39), .B1(new_n946), .B2(new_n956), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT39), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n960), .A2(new_n961), .A3(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1145), .A2(new_n1147), .B1(new_n966), .B2(new_n975), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n894), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n408), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n722), .B(new_n1150), .C1(new_n739), .C2(new_n743), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n893), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n958), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n975), .B1(new_n946), .B2(new_n956), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n773), .A2(G330), .A3(new_n896), .A4(new_n958), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1148), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n904), .A2(new_n893), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n976), .B1(new_n1158), .B2(new_n916), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1159), .A2(new_n973), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n917), .A2(G330), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n1027), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1157), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n545), .A2(new_n661), .A3(new_n713), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n765), .A2(new_n767), .ZN(new_n1166));
  OAI211_X1 g0966(.A(G330), .B(new_n896), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n916), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1168), .A2(new_n1156), .A3(new_n893), .A4(new_n1151), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n773), .A2(G330), .A3(new_n896), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1170), .A2(new_n916), .B1(new_n917), .B2(G330), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1171), .B2(new_n1158), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n673), .A2(G330), .A3(new_n912), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n672), .A2(new_n978), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1161), .B1(new_n1148), .B2(new_n1155), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1164), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT122), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1162), .A2(new_n1175), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n672), .A2(new_n978), .A3(new_n1173), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1170), .A2(new_n916), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1161), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1158), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1181), .B1(new_n1185), .B2(new_n1169), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1176), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n1157), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n782), .B1(new_n1188), .B2(KEYINPUT122), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1163), .B1(new_n1180), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n973), .A2(new_n794), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n399), .B1(new_n867), .B2(G137), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n835), .A2(G150), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1193), .A2(KEYINPUT53), .B1(G159), .B2(new_n811), .ZN(new_n1194));
  INV_X1    g0994(.A(G125), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n826), .A2(new_n201), .B1(new_n815), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1192), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n830), .A2(G128), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(KEYINPUT53), .B2(new_n1193), .C1(new_n841), .C2(new_n874), .ZN(new_n1200));
  XOR2_X1   g1000(.A(KEYINPUT54), .B(G143), .Z(new_n1201));
  AOI211_X1 g1001(.A(new_n1198), .B(new_n1200), .C1(new_n832), .C2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n841), .A2(new_n597), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n832), .A2(G97), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n878), .A2(G68), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1204), .A2(new_n836), .A3(new_n1205), .A4(new_n1127), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n399), .B1(new_n1105), .B2(new_n815), .C1(new_n825), .C2(new_n207), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n829), .A2(new_n859), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1203), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n797), .B1(new_n1202), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n263), .A2(new_n890), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1191), .A2(new_n863), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1190), .A2(new_n1212), .ZN(G378));
  NAND2_X1  g1013(.A1(new_n275), .A2(new_n712), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n322), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n322), .A2(new_n1214), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1215), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n794), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n867), .A2(G132), .B1(G137), .B2(new_n832), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G150), .A2(new_n811), .B1(new_n835), .B2(new_n1201), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n1195), .C2(new_n829), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G128), .B2(new_n842), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n345), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G41), .B(new_n1231), .C1(G124), .C2(new_n851), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n1229), .B2(new_n1228), .C1(new_n816), .C2(new_n826), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1097), .A2(new_n847), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G41), .B1(new_n842), .B2(G107), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G68), .A2(new_n811), .B1(new_n851), .B2(G283), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n460), .C2(new_n826), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1234), .B(new_n1237), .C1(G116), .C2(new_n830), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n457), .B1(new_n835), .B2(G77), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n206), .C2(new_n825), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT58), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n345), .B1(new_n412), .B2(new_n413), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n222), .B1(new_n1243), .B2(G41), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1233), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n797), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n890), .A2(new_n201), .ZN(new_n1248));
  AND4_X1   g1048(.A1(new_n863), .A2(new_n1224), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1222), .B1(new_n963), .B2(G330), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n962), .A2(new_n918), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n941), .A2(KEYINPUT112), .A3(new_n942), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT112), .B1(new_n941), .B2(new_n942), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n927), .B1(new_n468), .B2(new_n483), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n956), .B1(new_n1255), .B2(KEYINPUT38), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(KEYINPUT40), .A3(new_n917), .ZN(new_n1257));
  AND4_X1   g1057(.A1(G330), .A2(new_n1251), .A3(new_n1257), .A4(new_n1222), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n977), .B1(new_n1250), .B2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(new_n1257), .A3(G330), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1223), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n968), .B1(new_n1262), .B2(new_n975), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1251), .A2(new_n1257), .A3(new_n1222), .A4(G330), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1261), .A2(new_n967), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1259), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1249), .B1(new_n1266), .B2(new_n1026), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1187), .A2(new_n1186), .A3(new_n1157), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1268), .A2(new_n1174), .B1(new_n1259), .B2(new_n1265), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n781), .B1(new_n1269), .B2(KEYINPUT57), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1174), .B1(new_n1162), .B2(new_n1175), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1266), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT57), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1267), .B1(new_n1270), .B2(new_n1274), .ZN(G375));
  NAND2_X1  g1075(.A1(new_n1172), .A2(new_n1026), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n916), .A2(new_n391), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n834), .A2(new_n206), .B1(new_n826), .B2(new_n202), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1278), .B(new_n1098), .C1(G303), .C2(new_n851), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n867), .A2(G116), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n832), .A2(G107), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n841), .A2(new_n859), .B1(new_n1105), .B2(new_n829), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1282), .A2(new_n285), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .A4(new_n1283), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(G132), .A2(new_n830), .B1(new_n867), .B2(new_n1201), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n841), .B2(new_n1058), .ZN(new_n1286));
  XOR2_X1   g1086(.A(new_n1286), .B(KEYINPUT123), .Z(new_n1287));
  AOI22_X1  g1087(.A1(G159), .A2(new_n835), .B1(new_n851), .B2(G128), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n826), .A2(new_n460), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n454), .B(new_n1289), .C1(G50), .C2(new_n811), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n847), .A2(new_n1087), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1284), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n797), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n890), .A2(new_n326), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1277), .A2(new_n1294), .A3(new_n863), .A4(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1276), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1185), .A2(new_n1181), .A3(new_n1169), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1175), .A3(new_n1044), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(G381));
  INV_X1    g1101(.A(new_n1267), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n782), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1269), .A2(KEYINPUT57), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1302), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1212), .ZN(new_n1306));
  AOI211_X1 g1106(.A(new_n1306), .B(new_n1163), .C1(new_n1180), .C2(new_n1189), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1047), .A2(new_n1070), .A3(new_n1119), .A4(new_n1143), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1075), .A2(new_n793), .A3(new_n865), .A4(new_n1112), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(G384), .A2(G381), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1305), .A2(new_n1307), .A3(new_n1310), .A4(new_n1311), .ZN(G407));
  NAND2_X1  g1112(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n705), .A2(G343), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n705), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(KEYINPUT124), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(G407), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT125), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1318), .A2(KEYINPUT125), .A3(G407), .A4(new_n1319), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(G409));
  NAND3_X1  g1124(.A1(new_n1271), .A2(new_n1044), .A3(new_n1266), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1325), .A2(new_n1267), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1326), .A2(new_n1190), .A3(new_n1212), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1327), .B(new_n1315), .C1(new_n1305), .C2(new_n1307), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT126), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT60), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1330), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1172), .A2(new_n1174), .A3(new_n1330), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1329), .B1(new_n1335), .B2(new_n781), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1299), .B1(new_n1186), .B2(new_n1330), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1337), .A2(new_n1338), .A3(new_n1329), .A4(new_n781), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1298), .B1(new_n1336), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n909), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1337), .A2(new_n781), .A3(new_n1338), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(KEYINPUT126), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n1339), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1345), .A2(G384), .A3(new_n1298), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1314), .A2(G2897), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1342), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1347), .ZN(new_n1349));
  AOI21_X1  g1149(.A(G384), .B1(new_n1345), .B2(new_n1298), .ZN(new_n1350));
  AOI211_X1 g1150(.A(new_n909), .B(new_n1297), .C1(new_n1344), .C2(new_n1339), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1328), .A2(new_n1348), .A3(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(KEYINPUT63), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1314), .B1(new_n1307), .B2(new_n1326), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G375), .A2(G378), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1355), .A2(new_n1356), .A3(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1354), .A2(new_n1358), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1355), .A2(new_n1356), .A3(new_n1357), .A4(KEYINPUT63), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(G393), .A2(G396), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1309), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1308), .ZN(new_n1364));
  AOI22_X1  g1164(.A1(new_n1047), .A2(new_n1070), .B1(new_n1119), .B2(new_n1143), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1363), .B1(new_n1364), .B2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1365), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1367), .A2(new_n1362), .A3(new_n1308), .ZN(new_n1368));
  AND2_X1   g1168(.A1(new_n1366), .A2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT61), .ZN(new_n1370));
  AND3_X1   g1170(.A1(new_n1360), .A2(new_n1369), .A3(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1359), .A2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1342), .A2(new_n1346), .ZN(new_n1373));
  OAI21_X1  g1173(.A(KEYINPUT62), .B1(new_n1328), .B2(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT62), .ZN(new_n1375));
  NAND4_X1  g1175(.A1(new_n1355), .A2(new_n1356), .A3(new_n1357), .A4(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1374), .A2(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1353), .A2(new_n1370), .ZN(new_n1378));
  AND3_X1   g1178(.A1(new_n1366), .A2(new_n1368), .A3(KEYINPUT127), .ZN(new_n1379));
  AOI21_X1  g1179(.A(KEYINPUT127), .B1(new_n1366), .B2(new_n1368), .ZN(new_n1380));
  OAI22_X1  g1180(.A1(new_n1377), .A2(new_n1378), .B1(new_n1379), .B2(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1372), .A2(new_n1381), .ZN(G405));
  NOR2_X1   g1182(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1313), .A2(new_n1357), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1384), .A2(new_n1355), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1373), .A2(new_n1313), .A3(new_n1357), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1385), .A2(new_n1386), .ZN(new_n1387));
  XNOR2_X1  g1187(.A(new_n1383), .B(new_n1387), .ZN(G402));
endmodule


