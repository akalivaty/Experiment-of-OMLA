//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT69), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT70), .Z(G217));
  NOR4_X1   g028(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT71), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n461), .B(new_n462), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(G2106), .B2(new_n456), .ZN(G319));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n471), .C1(new_n466), .C2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n477), .A2(KEYINPUT72), .A3(G137), .A4(new_n471), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n477), .A2(G2105), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT74), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR3_X1    g060(.A1(new_n468), .A2(KEYINPUT73), .A3(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT73), .B1(new_n468), .B2(G2105), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  INV_X1    g064(.A(G100), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n490), .A2(new_n471), .A3(KEYINPUT75), .ZN(new_n491));
  AOI21_X1  g066(.A(KEYINPUT75), .B1(new_n490), .B2(new_n471), .ZN(new_n492));
  OAI221_X1 g067(.A(G2104), .B1(G112), .B2(new_n471), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n485), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n466), .B2(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n497), .B(new_n500), .C1(new_n467), .C2(new_n466), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n471), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n482), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n503), .A2(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT77), .B1(new_n510), .B2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n509), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G50), .A3(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n521), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n520), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT78), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n520), .A2(new_n524), .A3(new_n527), .A4(KEYINPUT78), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(G166));
  NAND2_X1  g107(.A1(new_n526), .A2(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n525), .A2(KEYINPUT79), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT79), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n521), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n534), .A2(G51), .A3(G543), .A4(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n515), .A2(new_n516), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n540), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n533), .A2(new_n537), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n521), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n534), .A2(G543), .A3(new_n536), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n540), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n548), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n544), .A2(new_n554), .B1(new_n546), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n540), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n550), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND4_X1  g139(.A1(new_n534), .A2(G53), .A3(G543), .A4(new_n536), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  XOR2_X1   g142(.A(KEYINPUT80), .B(G65), .Z(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n517), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n526), .B2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  NAND2_X1  g146(.A1(G168), .A2(KEYINPUT81), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n542), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n526), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n540), .B2(G74), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n534), .A2(G49), .A3(G543), .A4(new_n536), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n582));
  NAND2_X1  g157(.A1(G48), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n525), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n521), .A2(KEYINPUT82), .A3(G48), .A4(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n515), .A2(G61), .A3(new_n516), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n550), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  NOR3_X1   g166(.A1(new_n517), .A2(new_n591), .A3(new_n525), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(G305));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n544), .A2(new_n595), .B1(new_n546), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT83), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n540), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n550), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G54), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n546), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n544), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT84), .B(G66), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n515), .A2(new_n516), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G79), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n510), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT85), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n612), .B(new_n616), .C1(new_n613), .C2(new_n510), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n615), .A2(G651), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT86), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n610), .A2(new_n621), .A3(new_n618), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n603), .B1(new_n623), .B2(new_n602), .ZN(G284));
  AOI21_X1  g199(.A(new_n603), .B1(new_n623), .B2(new_n602), .ZN(G321));
  NOR2_X1   g200(.A1(G299), .A2(G868), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(new_n575), .B2(G868), .ZN(G297));
  AOI21_X1  g202(.A(new_n626), .B1(new_n575), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n623), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n477), .A2(new_n472), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(G111), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n639), .A2(KEYINPUT87), .B1(new_n640), .B2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(KEYINPUT87), .B2(new_n639), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n486), .A2(new_n487), .ZN(new_n643));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  INV_X1    g219(.A(G123), .ZN(new_n645));
  OAI221_X1 g220(.A(new_n642), .B1(new_n643), .B2(new_n644), .C1(new_n483), .C2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(G2096), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n638), .A2(new_n647), .A3(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT89), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2427), .B(G2430), .Z(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT88), .B(KEYINPUT14), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT90), .ZN(new_n658));
  INV_X1    g233(.A(G1341), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2451), .B(G2454), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XOR2_X1   g239(.A(G2443), .B(G2446), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT18), .Z(new_n677));
  INV_X1    g252(.A(new_n674), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n675), .B1(new_n678), .B2(new_n672), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT91), .B(KEYINPUT17), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n672), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n679), .B1(new_n682), .B2(new_n678), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n678), .A3(new_n675), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n677), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT92), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1956), .B(G2474), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n690), .B1(new_n692), .B2(new_n694), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n692), .A2(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n696), .B(new_n699), .C1(new_n689), .C2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n706), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(G229));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G33), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n488), .A2(G139), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT97), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n714));
  NAND3_X1  g289(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(G115), .A2(G2104), .ZN(new_n718));
  INV_X1    g293(.A(G127), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n468), .B2(new_n719), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n716), .A2(new_n717), .B1(G2105), .B2(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n711), .B1(new_n722), .B2(new_n710), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G2072), .Z(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT26), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n727), .A2(new_n728), .B1(G105), .B2(new_n472), .ZN(new_n729));
  INV_X1    g304(.A(G141), .ZN(new_n730));
  INV_X1    g305(.A(G129), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n729), .B1(new_n643), .B2(new_n730), .C1(new_n483), .C2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(new_n710), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n710), .B2(G32), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  INV_X1    g317(.A(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n743), .B2(KEYINPUT24), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(KEYINPUT24), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n480), .B2(new_n710), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n724), .B(new_n741), .C1(new_n742), .C2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT99), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n710), .A2(G26), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT28), .Z(new_n751));
  OR2_X1    g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n753));
  INV_X1    g328(.A(G140), .ZN(new_n754));
  INV_X1    g329(.A(G128), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n753), .B1(new_n643), .B2(new_n754), .C1(new_n483), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n751), .B1(new_n756), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G16), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G19), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n559), .B2(new_n760), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(new_n659), .ZN(new_n763));
  NOR2_X1   g338(.A1(G168), .A2(new_n760), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n760), .B2(G21), .ZN(new_n765));
  INV_X1    g340(.A(G1966), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n763), .B1(new_n767), .B2(KEYINPUT100), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n759), .B(new_n768), .C1(KEYINPUT100), .C2(new_n767), .ZN(new_n769));
  INV_X1    g344(.A(G28), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT30), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n770), .B2(KEYINPUT30), .ZN(new_n772));
  OR2_X1    g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  NAND2_X1  g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n710), .A2(G27), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n710), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n775), .B1(new_n777), .B2(G2078), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(G2078), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n646), .B2(new_n710), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n778), .B(new_n780), .C1(new_n742), .C2(new_n746), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n710), .A2(G35), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n710), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT29), .Z(new_n784));
  INV_X1    g359(.A(G2090), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n781), .B1(new_n766), .B2(new_n765), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n760), .A2(G5), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G171), .B2(new_n760), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT101), .Z(new_n789));
  INV_X1    g364(.A(G1961), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n739), .A2(new_n740), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n749), .A2(new_n769), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n760), .A2(G4), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n623), .B2(new_n760), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(G1348), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n760), .A2(G20), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT23), .Z(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G299), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G1956), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n784), .B2(new_n785), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n795), .A2(G1348), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n789), .A2(new_n790), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n747), .A2(new_n748), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n793), .A2(new_n796), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n760), .A2(G6), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G305), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT94), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT32), .B(G1981), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n760), .A2(G22), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G166), .B2(new_n760), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G1971), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n760), .A2(G23), .ZN(new_n817));
  INV_X1    g392(.A(G288), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n760), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT33), .B(G1976), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n819), .B(new_n820), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n814), .A2(G1971), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n812), .A2(new_n816), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT34), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n760), .A2(G24), .ZN(new_n827));
  INV_X1    g402(.A(G290), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n760), .ZN(new_n829));
  INV_X1    g404(.A(G1986), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n710), .A2(G25), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n484), .A2(G119), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n488), .A2(G131), .ZN(new_n834));
  OR2_X1    g409(.A1(G95), .A2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n832), .B1(new_n838), .B2(new_n710), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT35), .B(G1991), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT93), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n839), .B(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n825), .A2(new_n826), .A3(new_n831), .A4(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n807), .A2(new_n845), .A3(new_n846), .ZN(G311));
  NAND3_X1  g422(.A1(new_n807), .A2(new_n845), .A3(new_n846), .ZN(G150));
  NAND2_X1  g423(.A1(new_n623), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  INV_X1    g425(.A(G93), .ZN(new_n851));
  INV_X1    g426(.A(G55), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n544), .A2(new_n851), .B1(new_n546), .B2(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n540), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n550), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n559), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n850), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n859));
  AOI21_X1  g434(.A(G860), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n856), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(G145));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n868));
  INV_X1    g443(.A(new_n501), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n500), .B1(new_n477), .B2(new_n497), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n499), .A2(KEYINPUT103), .A3(new_n501), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n507), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n722), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n488), .A2(G142), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n471), .A2(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(G130), .B2(new_n484), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n636), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n874), .B(new_n880), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n736), .B(new_n756), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n838), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n874), .B(new_n880), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n882), .B(new_n837), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n494), .B(new_n646), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n480), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n884), .A2(new_n890), .A3(new_n887), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n864), .A2(G868), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n631), .B(new_n857), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n619), .B(G299), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n902), .B(KEYINPUT41), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n900), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G290), .B(G305), .ZN(new_n908));
  XNOR2_X1  g483(.A(G166), .B(new_n818), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n903), .B(KEYINPUT105), .C1(new_n901), .C2(new_n905), .ZN(new_n913));
  INV_X1    g488(.A(new_n911), .ZN(new_n914));
  INV_X1    g489(.A(new_n908), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n915), .A2(new_n909), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n909), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n907), .A2(new_n912), .A3(new_n913), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n912), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n904), .A2(new_n906), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(KEYINPUT105), .A3(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n897), .B(new_n899), .C1(new_n923), .C2(new_n602), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n602), .B1(new_n919), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT106), .B1(new_n925), .B2(new_n898), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(G295));
  NOR2_X1   g502(.A1(new_n925), .A2(new_n898), .ZN(G331));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  NAND2_X1  g504(.A1(G301), .A2(G168), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT107), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  NAND3_X1  g507(.A1(G301), .A2(new_n932), .A3(G168), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n931), .B(new_n933), .C1(new_n575), .C2(G301), .ZN(new_n934));
  INV_X1    g509(.A(new_n857), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G286), .A2(G171), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n937), .A2(new_n857), .A3(new_n933), .A4(new_n931), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n905), .ZN(new_n940));
  INV_X1    g515(.A(new_n902), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n910), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n910), .B1(new_n940), .B2(new_n942), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(G37), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n943), .A2(new_n944), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(KEYINPUT108), .A3(new_n893), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n893), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n953), .B2(new_n945), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n929), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n945), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n949), .A2(new_n951), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n953), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n957), .A2(KEYINPUT43), .B1(new_n958), .B2(new_n946), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n955), .B1(new_n929), .B2(new_n959), .ZN(G397));
  XNOR2_X1  g535(.A(new_n756), .B(new_n758), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n737), .B(new_n961), .C1(new_n962), .C2(G1996), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n873), .B2(G1384), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT110), .B(G40), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n473), .A2(new_n479), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(KEYINPUT111), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(KEYINPUT111), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n963), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n962), .B1(new_n971), .B2(G1996), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT127), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n978), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n736), .B(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n984), .A2(new_n838), .A3(new_n840), .A4(new_n961), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n756), .A2(G2067), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n971), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n971), .A2(G1986), .A3(G290), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(KEYINPUT48), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n838), .A2(new_n840), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n838), .A2(new_n840), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n984), .A2(new_n961), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n972), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(KEYINPUT48), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n987), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n982), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n980), .B1(new_n979), .B2(new_n981), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n873), .A2(G1384), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n473), .A2(new_n479), .A3(new_n966), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1976), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(G288), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1002), .B(new_n1004), .C1(new_n1003), .C2(G288), .ZN(new_n1005));
  INV_X1    g580(.A(G1981), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n590), .A2(new_n1006), .A3(new_n593), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT117), .B(G86), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n526), .A2(new_n1008), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n590), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(KEYINPUT49), .B(new_n1007), .C1(new_n1010), .C2(new_n1006), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1006), .B1(new_n590), .B2(new_n1009), .ZN(new_n1013));
  NOR4_X1   g588(.A1(new_n589), .A2(new_n586), .A3(new_n592), .A4(G1981), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1015), .A3(new_n1002), .ZN(new_n1016));
  INV_X1    g591(.A(new_n507), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n499), .A2(KEYINPUT103), .A3(new_n501), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT103), .B1(new_n499), .B2(new_n501), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1001), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1022), .B(G8), .C1(new_n1003), .C2(G288), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1023), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT116), .B1(new_n1023), .B2(KEYINPUT52), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1005), .B(new_n1016), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1000), .A2(KEYINPUT45), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1021), .B1(new_n503), .B2(new_n507), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n967), .B1(new_n1028), .B2(new_n964), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1971), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n873), .B2(G1384), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n1017), .B2(new_n502), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n967), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT113), .B(G2090), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1030), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(KEYINPUT114), .A3(new_n1036), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n999), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(KEYINPUT55), .ZN(new_n1043));
  OR3_X1    g618(.A1(G166), .A2(new_n999), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1042), .A2(KEYINPUT55), .ZN(new_n1045));
  OAI22_X1  g620(.A1(G166), .A2(new_n999), .B1(new_n1045), .B2(new_n1043), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1026), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1000), .A2(new_n1031), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1036), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1001), .B1(new_n1028), .B2(KEYINPUT50), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1052), .B2(new_n1030), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(new_n1046), .A3(new_n1044), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT45), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1055));
  INV_X1    g630(.A(new_n964), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1021), .B(new_n1056), .C1(new_n503), .C2(new_n507), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1001), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n766), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n473), .A2(new_n742), .A3(new_n479), .A4(new_n966), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT50), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n999), .B(G286), .C1(new_n1059), .C2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1048), .A2(KEYINPUT119), .A3(new_n1054), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1030), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n1040), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(G8), .A3(new_n1047), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1016), .A2(new_n1005), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1025), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1023), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1070), .A2(new_n1074), .A3(new_n1054), .A4(new_n1065), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT63), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1066), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1080), .A2(new_n1048), .A3(KEYINPUT63), .A4(new_n1065), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n800), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT56), .B(G2072), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1027), .A2(new_n1029), .A3(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1086));
  NAND2_X1  g661(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1083), .A2(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n622), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n621), .B1(new_n610), .B2(new_n618), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1035), .A2(G1348), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1000), .A2(new_n758), .A3(new_n1001), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1083), .A2(new_n1086), .A3(new_n1087), .A4(new_n1085), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1088), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1092), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT60), .B1(new_n1097), .B2(new_n1094), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1027), .A2(new_n983), .A3(new_n1029), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1027), .A2(KEYINPUT120), .A3(new_n983), .A4(new_n1029), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  NAND2_X1  g678(.A1(new_n1022), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n559), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1105), .A2(new_n559), .A3(new_n1107), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1098), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1095), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n1088), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(KEYINPUT61), .A3(new_n1095), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1092), .A2(new_n623), .A3(new_n1119), .A4(new_n1093), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1114), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1096), .B1(new_n1111), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n1123));
  OR4_X1    g698(.A1(new_n1123), .A2(new_n1055), .A3(new_n1058), .A4(G2078), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1125), .B2(G2078), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1124), .B(new_n1126), .C1(G1961), .C2(new_n1035), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G171), .ZN(new_n1128));
  INV_X1    g703(.A(G40), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1123), .A2(new_n1129), .A3(G2078), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1027), .A2(new_n965), .A3(G160), .A4(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1126), .B(new_n1131), .C1(G1961), .C2(new_n1035), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1128), .B1(G171), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1134));
  OR2_X1    g709(.A1(new_n1127), .A2(G171), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1132), .B2(G171), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1133), .A2(new_n1134), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n967), .B1(new_n1033), .B2(new_n1056), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT45), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n873), .B2(G1384), .ZN(new_n1141));
  AOI21_X1  g716(.A(G1966), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1060), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n542), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1059), .A2(new_n1064), .A3(G168), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(G8), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT51), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT51), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n1149), .A3(G8), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1122), .A2(new_n1138), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1070), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1016), .A2(new_n1003), .A3(new_n818), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1007), .B(KEYINPUT118), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1156), .A2(new_n1074), .B1(new_n1002), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1082), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1128), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1048), .A2(new_n1162), .A3(new_n1054), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT122), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1163), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT124), .B1(new_n1153), .B2(KEYINPUT62), .ZN(new_n1170));
  AND4_X1   g745(.A1(KEYINPUT124), .A2(new_n1165), .A3(new_n1166), .A4(KEYINPUT62), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT125), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1169), .B(new_n1174), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1161), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n971), .A2(new_n830), .A3(new_n828), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n988), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT112), .Z(new_n1179));
  INV_X1    g754(.A(new_n992), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n971), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n998), .B1(new_n1176), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g757(.A(G319), .ZN(new_n1184));
  NOR3_X1   g758(.A1(G229), .A2(new_n1184), .A3(G227), .ZN(new_n1185));
  NAND3_X1  g759(.A1(new_n895), .A2(new_n1185), .A3(new_n670), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n1186), .A2(new_n959), .ZN(G308));
  NAND2_X1  g761(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n958), .A2(new_n946), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g764(.A1(new_n1190), .A2(new_n670), .A3(new_n895), .A4(new_n1185), .ZN(G225));
endmodule


