//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  AND2_X1   g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(G197gat), .B(G204gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n209), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT64), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n221), .A2(G169gat), .A3(G176gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G169gat), .ZN(new_n225));
  INV_X1    g024(.A(G176gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT23), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n219), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n229), .A2(new_n232), .A3(new_n233), .A4(new_n217), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n220), .A2(new_n228), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n238), .A2(new_n239), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n238), .B2(new_n239), .ZN(new_n241));
  INV_X1    g040(.A(new_n218), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n221), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT25), .B1(new_n244), .B2(new_n223), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n223), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(KEYINPUT23), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n243), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n237), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT27), .B(G183gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n231), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n254), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257));
  OR3_X1    g056(.A1(new_n256), .A2(new_n223), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT26), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n248), .A2(new_n259), .A3(new_n249), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n257), .B1(new_n256), .B2(new_n223), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n253), .A2(new_n263), .A3(new_n231), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n255), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n252), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G226gat), .A2(G233gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT72), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n245), .B1(new_n242), .B2(new_n241), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n250), .A2(new_n271), .B1(new_n235), .B2(new_n236), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n255), .A2(new_n262), .A3(new_n264), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n252), .A2(KEYINPUT73), .A3(new_n265), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT29), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n267), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n216), .B(new_n269), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  AOI21_X1  g080(.A(new_n267), .B1(new_n274), .B2(new_n275), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n268), .B1(new_n266), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n215), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n286), .A2(KEYINPUT30), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n278), .A2(new_n285), .A3(new_n288), .A4(new_n281), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n278), .A2(new_n285), .ZN(new_n291));
  INV_X1    g090(.A(new_n281), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT74), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n294));
  AOI211_X1 g093(.A(new_n294), .B(new_n281), .C1(new_n278), .C2(new_n285), .ZN(new_n295));
  OAI22_X1  g094(.A1(new_n287), .A2(new_n290), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n298), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(KEYINPUT68), .ZN(new_n301));
  INV_X1    g100(.A(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G113gat), .ZN(new_n303));
  INV_X1    g102(.A(G113gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G120gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT1), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n305), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310));
  AND4_X1   g109(.A1(KEYINPUT69), .A2(new_n309), .A3(new_n300), .A4(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT69), .B1(new_n306), .B2(new_n300), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n315));
  INV_X1    g114(.A(G141gat), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n321), .A3(new_n319), .ZN(new_n322));
  INV_X1    g121(.A(new_n314), .ZN(new_n323));
  NOR2_X1   g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G155gat), .B(G162gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n329), .B(new_n315), .C1(new_n330), .C2(new_n321), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n326), .A2(new_n331), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n309), .A2(new_n300), .A3(new_n310), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n306), .A2(KEYINPUT69), .A3(new_n300), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(new_n339), .A3(new_n308), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n297), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n313), .B2(new_n332), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n326), .A2(new_n331), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n313), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT4), .A4(new_n308), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n346), .A2(new_n350), .A3(new_n342), .A4(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n350), .A2(new_n297), .A3(new_n342), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n313), .B2(new_n332), .ZN(new_n355));
  INV_X1    g154(.A(new_n345), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n334), .A2(new_n339), .A3(new_n308), .A4(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n344), .A2(new_n352), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G1gat), .B(G29gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT0), .ZN(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT81), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT6), .B1(new_n359), .B2(new_n363), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n313), .A2(new_n332), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n339), .A2(new_n308), .B1(new_n331), .B2(new_n326), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n343), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n368), .A3(KEYINPUT5), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n358), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n372));
  INV_X1    g171(.A(new_n363), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n364), .A2(new_n365), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n363), .B1(new_n369), .B2(new_n370), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT6), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n375), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n202), .B1(new_n296), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n313), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n272), .B2(new_n273), .ZN(new_n384));
  AND2_X1   g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n252), .A2(new_n313), .A3(new_n265), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT32), .ZN(new_n388));
  XOR2_X1   g187(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G15gat), .B(G43gat), .Z(new_n392));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n388), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n387), .B(KEYINPUT32), .C1(new_n390), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT34), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(KEYINPUT71), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(KEYINPUT71), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n397), .A3(new_n401), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n395), .A2(new_n397), .A3(new_n401), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n401), .B1(new_n395), .B2(new_n397), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT31), .B(G50gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT78), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n349), .A2(new_n283), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT80), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n349), .A2(new_n417), .A3(new_n283), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n215), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT29), .B1(new_n210), .B2(new_n214), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n332), .B1(new_n420), .B2(KEYINPUT3), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n414), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(KEYINPUT79), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(new_n332), .C1(new_n420), .C2(KEYINPUT3), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n415), .A2(new_n215), .ZN(new_n426));
  AND4_X1   g225(.A1(new_n414), .A2(new_n423), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(G22gat), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n418), .A2(new_n215), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n417), .B1(new_n349), .B2(new_n283), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n421), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n414), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n425), .A2(new_n414), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n421), .A2(KEYINPUT79), .B1(new_n415), .B2(new_n215), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G22gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G78gat), .B(G106gat), .ZN(new_n439));
  AND4_X1   g238(.A1(new_n413), .A2(new_n428), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n431), .A2(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT78), .B1(new_n441), .B2(new_n437), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n442), .B2(new_n428), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n412), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n439), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(new_n413), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n441), .A2(new_n437), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n428), .A3(new_n439), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n411), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n407), .A2(new_n410), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT35), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n291), .A2(new_n292), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n294), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n291), .A2(KEYINPUT74), .A3(new_n292), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n375), .A2(new_n379), .A3(new_n380), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n286), .A2(KEYINPUT30), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n289), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n456), .A2(KEYINPUT84), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n382), .A2(new_n451), .A3(new_n452), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n410), .A2(new_n407), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n450), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n365), .B1(KEYINPUT77), .B2(new_n376), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n376), .A2(KEYINPUT77), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n377), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n456), .A2(new_n467), .A3(new_n459), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT35), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT82), .B(KEYINPUT37), .Z(new_n471));
  NAND3_X1  g270(.A1(new_n278), .A2(new_n285), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n292), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n278), .B2(new_n285), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT38), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n215), .B(new_n269), .C1(new_n276), .C2(new_n277), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n216), .B1(new_n282), .B2(new_n284), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(KEYINPUT37), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n472), .A2(new_n479), .A3(new_n480), .A4(new_n292), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n381), .A2(new_n476), .A3(new_n481), .A4(new_n286), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT40), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT39), .B1(new_n341), .B2(new_n343), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n355), .A2(new_n350), .A3(new_n357), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n343), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n343), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n363), .B1(new_n487), .B2(KEYINPUT39), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n483), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(new_n364), .A3(new_n374), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n486), .A2(new_n488), .A3(new_n483), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n296), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n482), .A2(new_n463), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n410), .A2(new_n407), .A3(KEYINPUT36), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT36), .B1(new_n410), .B2(new_n407), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n444), .A2(new_n450), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n468), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n470), .A2(KEYINPUT85), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT85), .B1(new_n470), .B2(new_n500), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT87), .B(G29gat), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G36gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n508));
  OR3_X1    g307(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n505), .A2(new_n507), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT86), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n514), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n509), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n508), .B1(new_n517), .B2(new_n507), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n503), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT88), .A3(new_n512), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n524), .A3(G1gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT16), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G8gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n520), .B2(new_n512), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n535), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n533), .B(new_n534), .C1(new_n538), .C2(new_n532), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT90), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT18), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(KEYINPUT90), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n522), .A2(new_n532), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n533), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(new_n534), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G197gat), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT11), .B(G169gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT12), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n541), .A2(new_n556), .A3(new_n543), .A4(new_n548), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n501), .A2(new_n502), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G64gat), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G57gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n564), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT93), .ZN(new_n571));
  OR2_X1    g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n568), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n572), .B2(new_n568), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n570), .B(new_n571), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n568), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT93), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n569), .B1(new_n581), .B2(new_n574), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n583), .A2(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n584), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT20), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n584), .B(new_n585), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n532), .B1(KEYINPUT21), .B2(new_n583), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n590), .A2(new_n593), .A3(new_n597), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n599), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n562), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n602), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n561), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(G85gat), .ZN(new_n614));
  INV_X1    g413(.A(G92gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT8), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G99gat), .B(G106gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT97), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n619), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n617), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n538), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n522), .A2(new_n625), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G190gat), .B(G218gat), .Z(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n630), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n626), .A2(new_n635), .A3(new_n628), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n631), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n634), .B1(new_n631), .B2(new_n636), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n610), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n618), .B1(new_n623), .B2(KEYINPUT98), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n620), .A2(new_n644), .A3(new_n617), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n583), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(KEYINPUT93), .A3(new_n579), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n648), .A2(new_n621), .A3(new_n624), .A4(new_n577), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT99), .B(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n625), .A2(new_n583), .A3(KEYINPUT10), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n642), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n641), .B1(new_n646), .B2(new_n649), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  AOI21_X1  g457(.A(KEYINPUT100), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n655), .B2(new_n658), .ZN(new_n660));
  INV_X1    g459(.A(new_n658), .ZN(new_n661));
  OAI211_X1 g460(.A(KEYINPUT100), .B(new_n661), .C1(new_n653), .C2(new_n654), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n640), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n560), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n467), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT101), .B(G1gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1324gat));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND4_X1  g469(.A1(new_n560), .A2(new_n296), .A3(new_n665), .A4(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n296), .ZN(new_n672));
  OAI21_X1  g471(.A(G8gat), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n671), .ZN(new_n674));
  MUX2_X1   g473(.A(new_n671), .B(new_n674), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g474(.A(G15gat), .B1(new_n666), .B2(new_n497), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n560), .A2(new_n462), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n664), .A2(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n470), .A2(new_n500), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT85), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n470), .A2(KEYINPUT85), .A3(new_n500), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n682), .A2(new_n498), .A3(new_n683), .A4(new_n558), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n664), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT43), .B(G22gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  INV_X1    g486(.A(new_n467), .ZN(new_n688));
  INV_X1    g487(.A(new_n506), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n610), .A2(new_n639), .A3(new_n663), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n560), .A2(new_n688), .A3(new_n689), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n605), .A2(new_n609), .A3(KEYINPUT103), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT103), .B1(new_n605), .B2(new_n609), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n558), .A3(new_n663), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n639), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT44), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n410), .A2(new_n407), .A3(KEYINPUT36), .ZN(new_n702));
  INV_X1    g501(.A(new_n496), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n499), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n701), .B1(new_n704), .B2(new_n494), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n500), .A2(KEYINPUT104), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n470), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n639), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n698), .B1(new_n700), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(new_n688), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n694), .B1(new_n711), .B2(new_n689), .ZN(G1328gat));
  AOI21_X1  g511(.A(G36gat), .B1(KEYINPUT106), .B2(KEYINPUT46), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n560), .A2(new_n296), .A3(new_n691), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n710), .A2(new_n296), .ZN(new_n717));
  INV_X1    g516(.A(G36gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n690), .A2(G43gat), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n677), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n560), .A2(KEYINPUT107), .A3(new_n462), .A4(new_n721), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n497), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n710), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(G43gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n725), .B(KEYINPUT47), .C1(new_n727), .C2(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1330gat));
  NOR2_X1   g532(.A1(new_n690), .A2(G50gat), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n463), .B(new_n698), .C1(new_n700), .C2(new_n709), .ZN(new_n736));
  INV_X1    g535(.A(G50gat), .ZN(new_n737));
  OAI221_X1 g536(.A(KEYINPUT48), .B1(new_n684), .B2(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n560), .A2(new_n734), .A3(KEYINPUT108), .A4(new_n498), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n684), .B2(new_n735), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n736), .B2(new_n737), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n739), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n698), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n501), .A2(new_n502), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n639), .ZN(new_n751));
  INV_X1    g550(.A(new_n639), .ZN(new_n752));
  INV_X1    g551(.A(new_n708), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n704), .A2(new_n701), .A3(new_n494), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n500), .A2(KEYINPUT104), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI211_X1 g555(.A(new_n752), .B(new_n753), .C1(new_n756), .C2(new_n470), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n498), .B(new_n748), .C1(new_n751), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n743), .B1(new_n758), .B2(G50gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n759), .A2(KEYINPUT109), .A3(KEYINPUT48), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n738), .B1(new_n747), .B2(new_n760), .ZN(G1331gat));
  NOR4_X1   g560(.A1(new_n610), .A2(new_n558), .A3(new_n639), .A4(new_n663), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n707), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n467), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n563), .ZN(G1332gat));
  AND2_X1   g564(.A1(new_n707), .A2(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT110), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n296), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT49), .B(G64gat), .Z(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(G1333gat));
  INV_X1    g573(.A(G71gat), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n766), .A2(KEYINPUT111), .A3(new_n462), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT111), .B1(new_n766), .B2(new_n462), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n767), .A2(new_n726), .A3(new_n769), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G71gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1334gat));
  NAND2_X1  g582(.A1(new_n770), .A2(new_n498), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g584(.A1(new_n610), .A2(new_n559), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT112), .ZN(new_n787));
  INV_X1    g586(.A(new_n663), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n700), .B2(new_n709), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n688), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n707), .A2(new_n639), .A3(new_n787), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n707), .A2(KEYINPUT51), .A3(new_n639), .A4(new_n787), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(KEYINPUT113), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n792), .A2(new_n797), .A3(new_n793), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n788), .A2(new_n688), .A3(new_n614), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT114), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n614), .A2(new_n791), .B1(new_n799), .B2(new_n801), .ZN(G1336gat));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n794), .A2(new_n803), .A3(new_n795), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n296), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(G92gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n792), .A2(KEYINPUT115), .A3(new_n793), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n615), .B1(new_n790), .B2(new_n296), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT52), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n799), .A2(G92gat), .A3(new_n805), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n809), .A2(KEYINPUT52), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(G1337gat));
  NAND2_X1  g612(.A1(new_n790), .A2(new_n726), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G99gat), .ZN(new_n815));
  INV_X1    g614(.A(new_n462), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n663), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(G99gat), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n815), .B1(new_n799), .B2(new_n819), .ZN(G1338gat));
  NAND2_X1  g619(.A1(new_n790), .A2(new_n498), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G106gat), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n463), .A2(G106gat), .A3(new_n663), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n804), .A2(new_n807), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT53), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n796), .A2(new_n798), .A3(new_n824), .ZN(new_n827));
  XOR2_X1   g626(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n828));
  NAND3_X1  g627(.A1(new_n822), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n826), .A2(new_n829), .ZN(G1339gat));
  AND3_X1   g629(.A1(new_n651), .A2(new_n642), .A3(new_n652), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n831), .A2(new_n653), .A3(new_n832), .ZN(new_n833));
  AOI211_X1 g632(.A(KEYINPUT54), .B(new_n642), .C1(new_n651), .C2(new_n652), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(new_n658), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n651), .A2(new_n652), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n832), .A3(new_n641), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT117), .B1(new_n838), .B2(new_n661), .ZN(new_n839));
  OAI211_X1 g638(.A(KEYINPUT55), .B(new_n833), .C1(new_n836), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n655), .A2(new_n658), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(KEYINPUT118), .A3(new_n841), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n833), .B1(new_n836), .B2(new_n839), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n558), .A2(new_n844), .A3(new_n845), .A4(new_n848), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n538), .A2(new_n532), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n534), .B1(new_n850), .B2(new_n533), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n545), .A2(new_n547), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n553), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n788), .A2(new_n557), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n639), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n639), .A2(new_n557), .A3(new_n853), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n844), .A2(new_n848), .ZN(new_n857));
  INV_X1    g656(.A(new_n845), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n697), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n640), .A2(new_n559), .A3(new_n663), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n498), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n296), .A2(new_n467), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n816), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n559), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n467), .B1(new_n860), .B2(new_n861), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(new_n451), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n672), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n558), .A2(new_n304), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT120), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n867), .B1(new_n872), .B2(new_n874), .ZN(G1340gat));
  NOR3_X1   g674(.A1(new_n864), .A2(new_n302), .A3(new_n818), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n872), .A2(new_n663), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n302), .ZN(G1341gat));
  OAI21_X1  g677(.A(G127gat), .B1(new_n866), .B2(new_n697), .ZN(new_n879));
  INV_X1    g678(.A(new_n610), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n298), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n872), .B2(new_n881), .ZN(G1342gat));
  NOR2_X1   g681(.A1(new_n752), .A2(G134gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n872), .A2(KEYINPUT56), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n866), .B2(new_n752), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT56), .B1(new_n872), .B2(new_n884), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(G1343gat));
  NAND2_X1  g687(.A1(new_n497), .A2(new_n863), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n463), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n842), .B1(new_n555), .B2(new_n557), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n831), .A2(new_n653), .A3(new_n832), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n835), .B1(new_n834), .B2(new_n658), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n838), .A2(KEYINPUT117), .A3(new_n661), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n847), .B1(new_n897), .B2(KEYINPUT121), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n899), .B(new_n894), .C1(new_n896), .C2(new_n895), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n893), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT55), .B1(new_n846), .B2(new_n899), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(KEYINPUT122), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n892), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n854), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n854), .A3(KEYINPUT123), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n752), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n859), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n880), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n861), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n891), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n860), .A2(new_n861), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n498), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n890), .ZN(new_n917));
  AOI211_X1 g716(.A(new_n559), .B(new_n889), .C1(new_n914), .C2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT124), .B1(new_n918), .B2(new_n316), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n726), .A2(new_n463), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n868), .A2(new_n672), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n316), .A3(new_n558), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n918), .B2(new_n316), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n919), .A2(new_n923), .A3(KEYINPUT58), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT58), .ZN(new_n925));
  OAI221_X1 g724(.A(new_n922), .B1(KEYINPUT124), .B2(new_n925), .C1(new_n918), .C2(new_n316), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1344gat));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n317), .A3(new_n788), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n889), .B1(new_n914), .B2(new_n917), .ZN(new_n929));
  AOI211_X1 g728(.A(KEYINPUT59), .B(new_n317), .C1(new_n929), .C2(new_n788), .ZN(new_n930));
  XNOR2_X1  g729(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n890), .B(new_n498), .C1(new_n912), .C2(new_n913), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT57), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n889), .A2(new_n663), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(G148gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n928), .B1(new_n930), .B2(new_n936), .ZN(G1345gat));
  INV_X1    g736(.A(G155gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n938), .A3(new_n880), .ZN(new_n939));
  AOI211_X1 g738(.A(new_n697), .B(new_n889), .C1(new_n914), .C2(new_n917), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n938), .ZN(G1346gat));
  AOI21_X1  g740(.A(G162gat), .B1(new_n921), .B2(new_n639), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n639), .A2(G162gat), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n929), .B2(new_n943), .ZN(G1347gat));
  NAND2_X1  g743(.A1(new_n296), .A2(new_n467), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n816), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n862), .A2(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n947), .A2(new_n225), .A3(new_n559), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n688), .B1(new_n860), .B2(new_n861), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(new_n296), .A3(new_n451), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n558), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n225), .B2(new_n951), .ZN(G1348gat));
  NOR3_X1   g751(.A1(new_n947), .A2(new_n226), .A3(new_n663), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n788), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n226), .B2(new_n954), .ZN(G1349gat));
  OR2_X1    g754(.A1(new_n947), .A2(new_n697), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n880), .A2(new_n253), .ZN(new_n957));
  AOI22_X1  g756(.A1(new_n956), .A2(G183gat), .B1(new_n950), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g758(.A1(new_n950), .A2(new_n231), .A3(new_n639), .ZN(new_n960));
  OAI21_X1  g759(.A(G190gat), .B1(new_n947), .B2(new_n752), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n961), .A2(KEYINPUT61), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n961), .A2(KEYINPUT61), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1351gat));
  AND2_X1   g763(.A1(new_n949), .A2(new_n920), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n296), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  XOR2_X1   g766(.A(KEYINPUT126), .B(G197gat), .Z(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n558), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n726), .A2(new_n945), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n932), .A2(new_n933), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(new_n559), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n972), .B2(new_n968), .ZN(G1352gat));
  NOR2_X1   g772(.A1(new_n805), .A2(G204gat), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n975), .B(KEYINPUT62), .Z(new_n976));
  OAI21_X1  g775(.A(G204gat), .B1(new_n971), .B2(new_n663), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1353gat));
  NOR3_X1   g777(.A1(new_n966), .A2(G211gat), .A3(new_n610), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n979), .B(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(G211gat), .B1(new_n971), .B2(new_n610), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n982), .A2(KEYINPUT63), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(KEYINPUT63), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(G1354gat));
  OAI21_X1  g784(.A(G218gat), .B1(new_n971), .B2(new_n752), .ZN(new_n986));
  OR3_X1    g785(.A1(new_n966), .A2(G218gat), .A3(new_n752), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1355gat));
endmodule


