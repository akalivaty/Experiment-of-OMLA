

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X2 U547 ( .A(KEYINPUT64), .B(n516), .Z(n856) );
  NAND2_X1 U548 ( .A1(n786), .A2(n679), .ZN(n728) );
  XNOR2_X1 U549 ( .A(n765), .B(n764), .ZN(n766) );
  INV_X1 U550 ( .A(KEYINPUT26), .ZN(n686) );
  INV_X1 U551 ( .A(n728), .ZN(n705) );
  AND2_X1 U552 ( .A1(n736), .A2(n735), .ZN(n737) );
  OR2_X1 U553 ( .A1(n725), .A2(n724), .ZN(n755) );
  INV_X1 U554 ( .A(KEYINPUT97), .ZN(n764) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n786) );
  NOR2_X1 U556 ( .A1(G651), .A2(n639), .ZN(n638) );
  NOR2_X1 U557 ( .A1(G651), .A2(G543), .ZN(n635) );
  OR2_X1 U558 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U559 ( .A(n521), .B(KEYINPUT83), .ZN(G164) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n512) );
  XOR2_X2 U561 ( .A(KEYINPUT17), .B(n512), .Z(n860) );
  NAND2_X1 U562 ( .A1(G138), .A2(n860), .ZN(n514) );
  INV_X1 U563 ( .A(G2105), .ZN(n515) );
  NOR2_X1 U564 ( .A1(G2104), .A2(n515), .ZN(n855) );
  NAND2_X1 U565 ( .A1(G126), .A2(n855), .ZN(n513) );
  NAND2_X1 U566 ( .A1(n514), .A2(n513), .ZN(n520) );
  AND2_X1 U567 ( .A1(n515), .A2(G2104), .ZN(n859) );
  NAND2_X1 U568 ( .A1(G102), .A2(n859), .ZN(n518) );
  NAND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  NAND2_X1 U570 ( .A1(G114), .A2(n856), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n518), .A2(n517), .ZN(n519) );
  INV_X1 U572 ( .A(G651), .ZN(n525) );
  NOR2_X1 U573 ( .A1(G543), .A2(n525), .ZN(n522) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n522), .Z(n643) );
  NAND2_X1 U575 ( .A1(G60), .A2(n643), .ZN(n524) );
  NAND2_X1 U576 ( .A1(G85), .A2(n635), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n524), .A2(n523), .ZN(n529) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  NOR2_X1 U579 ( .A1(n639), .A2(n525), .ZN(n631) );
  NAND2_X1 U580 ( .A1(G72), .A2(n631), .ZN(n527) );
  NAND2_X1 U581 ( .A1(G47), .A2(n638), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  OR2_X1 U583 ( .A1(n529), .A2(n528), .ZN(G290) );
  XNOR2_X1 U584 ( .A(G2435), .B(G2443), .ZN(n539) );
  XOR2_X1 U585 ( .A(G2454), .B(G2430), .Z(n531) );
  XNOR2_X1 U586 ( .A(G2446), .B(KEYINPUT101), .ZN(n530) );
  XNOR2_X1 U587 ( .A(n531), .B(n530), .ZN(n535) );
  XOR2_X1 U588 ( .A(G2451), .B(G2427), .Z(n533) );
  XNOR2_X1 U589 ( .A(G1341), .B(G1348), .ZN(n532) );
  XNOR2_X1 U590 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U591 ( .A(n535), .B(n534), .Z(n537) );
  XNOR2_X1 U592 ( .A(KEYINPUT102), .B(G2438), .ZN(n536) );
  XNOR2_X1 U593 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U594 ( .A(n539), .B(n538), .ZN(n540) );
  AND2_X1 U595 ( .A1(n540), .A2(G14), .ZN(G401) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U597 ( .A1(G123), .A2(n855), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n541), .B(KEYINPUT18), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n859), .A2(G99), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G135), .A2(n860), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G111), .A2(n856), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n957) );
  XNOR2_X1 U605 ( .A(n957), .B(G2096), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n548), .B(KEYINPUT75), .ZN(n549) );
  OR2_X1 U607 ( .A1(G2100), .A2(n549), .ZN(G156) );
  INV_X1 U608 ( .A(G132), .ZN(G219) );
  INV_X1 U609 ( .A(G82), .ZN(G220) );
  NAND2_X1 U610 ( .A1(G75), .A2(n631), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G88), .A2(n635), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G50), .A2(n638), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n552), .B(KEYINPUT78), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n643), .A2(G62), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U617 ( .A1(n556), .A2(n555), .ZN(G166) );
  NAND2_X1 U618 ( .A1(n638), .A2(G52), .ZN(n557) );
  XNOR2_X1 U619 ( .A(KEYINPUT65), .B(n557), .ZN(n566) );
  NAND2_X1 U620 ( .A1(n635), .A2(G90), .ZN(n558) );
  XNOR2_X1 U621 ( .A(n558), .B(KEYINPUT66), .ZN(n560) );
  NAND2_X1 U622 ( .A1(G77), .A2(n631), .ZN(n559) );
  NAND2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  XNOR2_X1 U625 ( .A(n562), .B(KEYINPUT67), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G64), .A2(n643), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U628 ( .A1(n566), .A2(n565), .ZN(G171) );
  NAND2_X1 U629 ( .A1(n635), .A2(G89), .ZN(n567) );
  XNOR2_X1 U630 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G76), .A2(n631), .ZN(n568) );
  NAND2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT5), .ZN(n576) );
  XNOR2_X1 U634 ( .A(KEYINPUT6), .B(KEYINPUT73), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G63), .A2(n643), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G51), .A2(n638), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT7), .B(n577), .ZN(G168) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U642 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U644 ( .A(G223), .ZN(n822) );
  NAND2_X1 U645 ( .A1(n822), .A2(G567), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  NAND2_X1 U647 ( .A1(n643), .A2(G56), .ZN(n580) );
  XNOR2_X1 U648 ( .A(KEYINPUT14), .B(n580), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n635), .A2(G81), .ZN(n581) );
  XNOR2_X1 U650 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G68), .A2(n631), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U653 ( .A(KEYINPUT13), .B(n584), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT71), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n638), .A2(G43), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n987) );
  INV_X1 U658 ( .A(G860), .ZN(n612) );
  OR2_X1 U659 ( .A1(n987), .A2(n612), .ZN(G153) );
  INV_X1 U660 ( .A(G171), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U662 ( .A1(n638), .A2(G54), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G66), .A2(n643), .ZN(n591) );
  NAND2_X1 U664 ( .A1(G92), .A2(n635), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n631), .A2(G79), .ZN(n592) );
  XOR2_X1 U667 ( .A(KEYINPUT72), .B(n592), .Z(n593) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U670 ( .A(KEYINPUT15), .B(n597), .Z(n1000) );
  INV_X1 U671 ( .A(G868), .ZN(n609) );
  NAND2_X1 U672 ( .A1(n1000), .A2(n609), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U674 ( .A1(n643), .A2(G65), .ZN(n600) );
  XNOR2_X1 U675 ( .A(n600), .B(KEYINPUT68), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G53), .A2(n638), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT69), .B(n603), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n631), .A2(G78), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G91), .A2(n635), .ZN(n604) );
  AND2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(G299) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n608), .B(KEYINPUT74), .ZN(n611) );
  NOR2_X1 U685 ( .A1(n609), .A2(G286), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n612), .A2(G559), .ZN(n613) );
  INV_X1 U688 ( .A(n1000), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n613), .A2(n618), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n614), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U691 ( .A1(G868), .A2(n987), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(G868), .ZN(n615) );
  NOR2_X1 U693 ( .A1(G559), .A2(n615), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G559), .A2(n618), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n987), .B(n619), .ZN(n654) );
  NOR2_X1 U697 ( .A1(n654), .A2(G860), .ZN(n628) );
  NAND2_X1 U698 ( .A1(G80), .A2(n631), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G93), .A2(n635), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n643), .A2(G67), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n622), .B(KEYINPUT76), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G55), .A2(n638), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U705 ( .A(KEYINPUT77), .B(n625), .Z(n626) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n651) );
  XNOR2_X1 U707 ( .A(n628), .B(n651), .ZN(G145) );
  NAND2_X1 U708 ( .A1(G61), .A2(n643), .ZN(n630) );
  NAND2_X1 U709 ( .A1(G48), .A2(n638), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G73), .A2(n631), .ZN(n632) );
  XOR2_X1 U712 ( .A(KEYINPUT2), .B(n632), .Z(n633) );
  NOR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n635), .A2(G86), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U716 ( .A1(G49), .A2(n638), .ZN(n641) );
  NAND2_X1 U717 ( .A1(G87), .A2(n639), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G651), .A2(G74), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(G288) );
  NOR2_X1 U722 ( .A1(G868), .A2(n651), .ZN(n646) );
  XOR2_X1 U723 ( .A(n646), .B(KEYINPUT80), .Z(n657) );
  INV_X1 U724 ( .A(G299), .ZN(n988) );
  XNOR2_X1 U725 ( .A(n988), .B(G305), .ZN(n647) );
  XNOR2_X1 U726 ( .A(n647), .B(G290), .ZN(n650) );
  XOR2_X1 U727 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n648) );
  XNOR2_X1 U728 ( .A(G288), .B(n648), .ZN(n649) );
  XOR2_X1 U729 ( .A(n650), .B(n649), .Z(n653) );
  XNOR2_X1 U730 ( .A(G166), .B(n651), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n874) );
  XOR2_X1 U732 ( .A(n874), .B(n654), .Z(n655) );
  NAND2_X1 U733 ( .A1(G868), .A2(n655), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2078), .A2(G2084), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n658), .B(KEYINPUT81), .ZN(n659) );
  XNOR2_X1 U737 ( .A(KEYINPUT20), .B(n659), .ZN(n660) );
  NAND2_X1 U738 ( .A1(n660), .A2(G2090), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(KEYINPUT82), .ZN(n662) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XOR2_X1 U742 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U744 ( .A1(G108), .A2(G120), .ZN(n664) );
  NOR2_X1 U745 ( .A1(G237), .A2(n664), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G69), .A2(n665), .ZN(n827) );
  NAND2_X1 U747 ( .A1(n827), .A2(G567), .ZN(n670) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U750 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U751 ( .A1(G96), .A2(n668), .ZN(n828) );
  NAND2_X1 U752 ( .A1(n828), .A2(G2106), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n670), .A2(n669), .ZN(n829) );
  NAND2_X1 U754 ( .A1(G483), .A2(G661), .ZN(n671) );
  NOR2_X1 U755 ( .A1(n829), .A2(n671), .ZN(n826) );
  NAND2_X1 U756 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U757 ( .A1(n860), .A2(G137), .ZN(n674) );
  NAND2_X1 U758 ( .A1(G101), .A2(n859), .ZN(n672) );
  XOR2_X1 U759 ( .A(KEYINPUT23), .B(n672), .Z(n673) );
  NAND2_X1 U760 ( .A1(n674), .A2(n673), .ZN(n678) );
  NAND2_X1 U761 ( .A1(G125), .A2(n855), .ZN(n676) );
  NAND2_X1 U762 ( .A1(G113), .A2(n856), .ZN(n675) );
  NAND2_X1 U763 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U764 ( .A1(n678), .A2(n677), .ZN(G160) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n785) );
  INV_X1 U767 ( .A(n785), .ZN(n679) );
  NAND2_X1 U768 ( .A1(G8), .A2(n728), .ZN(n760) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n680) );
  XOR2_X1 U770 ( .A(n680), .B(KEYINPUT24), .Z(n681) );
  NOR2_X1 U771 ( .A1(n760), .A2(n681), .ZN(n767) );
  NAND2_X1 U772 ( .A1(n705), .A2(G2072), .ZN(n682) );
  XNOR2_X1 U773 ( .A(n682), .B(KEYINPUT27), .ZN(n684) );
  INV_X1 U774 ( .A(G1956), .ZN(n903) );
  NOR2_X1 U775 ( .A1(n903), .A2(n705), .ZN(n683) );
  NOR2_X1 U776 ( .A1(n684), .A2(n683), .ZN(n698) );
  OR2_X1 U777 ( .A1(n698), .A2(n988), .ZN(n685) );
  XNOR2_X1 U778 ( .A(n685), .B(KEYINPUT28), .ZN(n702) );
  INV_X1 U779 ( .A(G1996), .ZN(n932) );
  NOR2_X1 U780 ( .A1(n728), .A2(n932), .ZN(n687) );
  XNOR2_X1 U781 ( .A(n687), .B(n686), .ZN(n689) );
  NAND2_X1 U782 ( .A1(n728), .A2(G1341), .ZN(n688) );
  NAND2_X1 U783 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U784 ( .A1(n987), .A2(n690), .ZN(n694) );
  NAND2_X1 U785 ( .A1(G1348), .A2(n728), .ZN(n692) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n705), .ZN(n691) );
  NAND2_X1 U787 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U788 ( .A1(n1000), .A2(n695), .ZN(n693) );
  OR2_X1 U789 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n1000), .A2(n695), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n988), .A2(n698), .ZN(n699) );
  NAND2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U795 ( .A(KEYINPUT29), .B(n703), .Z(n710) );
  XOR2_X1 U796 ( .A(G1961), .B(KEYINPUT90), .Z(n915) );
  NAND2_X1 U797 ( .A1(n915), .A2(n728), .ZN(n707) );
  XOR2_X1 U798 ( .A(G2078), .B(KEYINPUT25), .Z(n704) );
  XNOR2_X1 U799 ( .A(KEYINPUT91), .B(n704), .ZN(n931) );
  NAND2_X1 U800 ( .A1(n705), .A2(n931), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n714) );
  NAND2_X1 U802 ( .A1(G171), .A2(n714), .ZN(n708) );
  XNOR2_X1 U803 ( .A(n708), .B(KEYINPUT92), .ZN(n709) );
  NAND2_X1 U804 ( .A1(n710), .A2(n709), .ZN(n719) );
  NOR2_X1 U805 ( .A1(G2084), .A2(n728), .ZN(n723) );
  NOR2_X1 U806 ( .A1(G1966), .A2(n760), .ZN(n720) );
  NOR2_X1 U807 ( .A1(n723), .A2(n720), .ZN(n711) );
  NAND2_X1 U808 ( .A1(G8), .A2(n711), .ZN(n712) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n712), .ZN(n713) );
  NOR2_X1 U810 ( .A1(G168), .A2(n713), .ZN(n716) );
  NOR2_X1 U811 ( .A1(G171), .A2(n714), .ZN(n715) );
  NOR2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U813 ( .A(KEYINPUT31), .B(n717), .Z(n718) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n727) );
  INV_X1 U815 ( .A(n727), .ZN(n721) );
  NOR2_X1 U816 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U817 ( .A(n722), .B(KEYINPUT93), .ZN(n725) );
  AND2_X1 U818 ( .A1(G8), .A2(n723), .ZN(n724) );
  AND2_X1 U819 ( .A1(G286), .A2(G8), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n736) );
  INV_X1 U821 ( .A(G8), .ZN(n734) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n760), .ZN(n730) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n731), .A2(G303), .ZN(n732) );
  XNOR2_X1 U826 ( .A(n732), .B(KEYINPUT94), .ZN(n733) );
  OR2_X1 U827 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U828 ( .A(n737), .B(KEYINPUT32), .ZN(n756) );
  INV_X1 U829 ( .A(KEYINPUT33), .ZN(n743) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n996) );
  INV_X1 U831 ( .A(n760), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n996), .A2(n738), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n743), .A2(n739), .ZN(n741) );
  AND2_X1 U834 ( .A1(n756), .A2(n741), .ZN(n740) );
  NAND2_X1 U835 ( .A1(n755), .A2(n740), .ZN(n747) );
  INV_X1 U836 ( .A(n741), .ZN(n745) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n742) );
  NOR2_X1 U839 ( .A1(n749), .A2(n742), .ZN(n997) );
  AND2_X1 U840 ( .A1(n997), .A2(n743), .ZN(n744) );
  OR2_X1 U841 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U842 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U843 ( .A(n748), .B(KEYINPUT95), .ZN(n753) );
  XNOR2_X1 U844 ( .A(G1981), .B(G305), .ZN(n992) );
  NAND2_X1 U845 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U846 ( .A1(n760), .A2(n750), .ZN(n751) );
  NOR2_X1 U847 ( .A1(n992), .A2(n751), .ZN(n752) );
  NAND2_X1 U848 ( .A1(n753), .A2(n752), .ZN(n763) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n754) );
  NAND2_X1 U850 ( .A1(G8), .A2(n754), .ZN(n758) );
  NAND2_X1 U851 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U852 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U853 ( .A(n759), .B(KEYINPUT96), .ZN(n761) );
  NAND2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n765) );
  NOR2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n801) );
  NAND2_X1 U857 ( .A1(n856), .A2(G107), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G95), .A2(n859), .ZN(n769) );
  NAND2_X1 U859 ( .A1(G131), .A2(n860), .ZN(n768) );
  NAND2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U861 ( .A1(G119), .A2(n855), .ZN(n770) );
  XNOR2_X1 U862 ( .A(KEYINPUT87), .B(n770), .ZN(n771) );
  NOR2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U865 ( .A(n775), .B(KEYINPUT88), .ZN(n848) );
  NAND2_X1 U866 ( .A1(G1991), .A2(n848), .ZN(n784) );
  NAND2_X1 U867 ( .A1(G129), .A2(n855), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G141), .A2(n860), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G105), .A2(n859), .ZN(n778) );
  XOR2_X1 U871 ( .A(KEYINPUT38), .B(n778), .Z(n779) );
  NOR2_X1 U872 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G117), .A2(n856), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n866) );
  NAND2_X1 U875 ( .A1(G1996), .A2(n866), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n956) );
  NOR2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n816) );
  NAND2_X1 U878 ( .A1(n956), .A2(n816), .ZN(n787) );
  XNOR2_X1 U879 ( .A(n787), .B(KEYINPUT89), .ZN(n808) );
  INV_X1 U880 ( .A(n808), .ZN(n799) );
  NAND2_X1 U881 ( .A1(G104), .A2(n859), .ZN(n789) );
  NAND2_X1 U882 ( .A1(G140), .A2(n860), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U884 ( .A(KEYINPUT34), .B(n790), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G128), .A2(n855), .ZN(n792) );
  NAND2_X1 U886 ( .A1(G116), .A2(n856), .ZN(n791) );
  NAND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U888 ( .A(n793), .B(KEYINPUT35), .Z(n794) );
  NOR2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U890 ( .A(KEYINPUT36), .B(n796), .Z(n797) );
  XNOR2_X1 U891 ( .A(KEYINPUT85), .B(n797), .ZN(n852) );
  XNOR2_X1 U892 ( .A(KEYINPUT37), .B(G2067), .ZN(n805) );
  NOR2_X1 U893 ( .A1(n852), .A2(n805), .ZN(n798) );
  XNOR2_X1 U894 ( .A(n798), .B(KEYINPUT86), .ZN(n961) );
  NAND2_X1 U895 ( .A1(n816), .A2(n961), .ZN(n812) );
  NAND2_X1 U896 ( .A1(n799), .A2(n812), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n804) );
  XNOR2_X1 U898 ( .A(KEYINPUT84), .B(G1986), .ZN(n802) );
  XNOR2_X1 U899 ( .A(n802), .B(G290), .ZN(n1007) );
  NAND2_X1 U900 ( .A1(n816), .A2(n1007), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n819) );
  NAND2_X1 U902 ( .A1(n805), .A2(n852), .ZN(n976) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n866), .ZN(n965) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U905 ( .A1(n848), .A2(G1991), .ZN(n958) );
  NOR2_X1 U906 ( .A1(n806), .A2(n958), .ZN(n807) );
  NOR2_X1 U907 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U908 ( .A(n809), .B(KEYINPUT98), .ZN(n810) );
  NOR2_X1 U909 ( .A1(n965), .A2(n810), .ZN(n811) );
  XNOR2_X1 U910 ( .A(n811), .B(KEYINPUT39), .ZN(n813) );
  NAND2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n976), .A2(n814), .ZN(n815) );
  NAND2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U914 ( .A(KEYINPUT99), .B(n817), .Z(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n821) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n821), .B(n820), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U920 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n824) );
  XOR2_X1 U922 ( .A(KEYINPUT103), .B(n824), .Z(n825) );
  NAND2_X1 U923 ( .A1(n826), .A2(n825), .ZN(G188) );
  XOR2_X1 U924 ( .A(G96), .B(KEYINPUT104), .Z(G221) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  INV_X1 U927 ( .A(G108), .ZN(G238) );
  INV_X1 U928 ( .A(G69), .ZN(G235) );
  NOR2_X1 U929 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  INV_X1 U931 ( .A(n829), .ZN(G319) );
  NAND2_X1 U932 ( .A1(G124), .A2(n855), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n830), .B(KEYINPUT44), .ZN(n831) );
  XNOR2_X1 U934 ( .A(n831), .B(KEYINPUT106), .ZN(n833) );
  NAND2_X1 U935 ( .A1(G100), .A2(n859), .ZN(n832) );
  NAND2_X1 U936 ( .A1(n833), .A2(n832), .ZN(n837) );
  NAND2_X1 U937 ( .A1(G136), .A2(n860), .ZN(n835) );
  NAND2_X1 U938 ( .A1(G112), .A2(n856), .ZN(n834) );
  NAND2_X1 U939 ( .A1(n835), .A2(n834), .ZN(n836) );
  NOR2_X1 U940 ( .A1(n837), .A2(n836), .ZN(G162) );
  XOR2_X1 U941 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n839) );
  XNOR2_X1 U942 ( .A(G164), .B(G160), .ZN(n838) );
  XNOR2_X1 U943 ( .A(n839), .B(n838), .ZN(n851) );
  NAND2_X1 U944 ( .A1(G103), .A2(n859), .ZN(n841) );
  NAND2_X1 U945 ( .A1(G139), .A2(n860), .ZN(n840) );
  NAND2_X1 U946 ( .A1(n841), .A2(n840), .ZN(n847) );
  NAND2_X1 U947 ( .A1(n855), .A2(G127), .ZN(n842) );
  XOR2_X1 U948 ( .A(KEYINPUT107), .B(n842), .Z(n844) );
  NAND2_X1 U949 ( .A1(G115), .A2(n856), .ZN(n843) );
  NAND2_X1 U950 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U951 ( .A(KEYINPUT47), .B(n845), .Z(n846) );
  NOR2_X1 U952 ( .A1(n847), .A2(n846), .ZN(n970) );
  XNOR2_X1 U953 ( .A(n848), .B(n970), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n849), .B(n957), .ZN(n850) );
  XNOR2_X1 U955 ( .A(n851), .B(n850), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n852), .B(KEYINPUT108), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n870) );
  NAND2_X1 U958 ( .A1(G130), .A2(n855), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G118), .A2(n856), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G106), .A2(n859), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G142), .A2(n860), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(n863), .B(KEYINPUT45), .Z(n864) );
  NOR2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U967 ( .A(G162), .B(n868), .Z(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n871) );
  NOR2_X1 U969 ( .A1(G37), .A2(n871), .ZN(G395) );
  XNOR2_X1 U970 ( .A(G286), .B(KEYINPUT109), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n1000), .B(G171), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n876) );
  XNOR2_X1 U973 ( .A(n987), .B(n874), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n877) );
  NOR2_X1 U975 ( .A1(G37), .A2(n877), .ZN(G397) );
  XOR2_X1 U976 ( .A(G1976), .B(G1971), .Z(n879) );
  XNOR2_X1 U977 ( .A(G1981), .B(G1966), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U979 ( .A(n880), .B(G2474), .Z(n882) );
  XNOR2_X1 U980 ( .A(G1996), .B(G1991), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n886) );
  XOR2_X1 U982 ( .A(KEYINPUT41), .B(G1986), .Z(n884) );
  XNOR2_X1 U983 ( .A(G1956), .B(G1961), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(G229) );
  XOR2_X1 U986 ( .A(KEYINPUT105), .B(G2078), .Z(n888) );
  XNOR2_X1 U987 ( .A(G2090), .B(G2072), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(n889), .B(G2100), .Z(n891) );
  XNOR2_X1 U990 ( .A(G2067), .B(G2084), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U992 ( .A(G2096), .B(KEYINPUT43), .Z(n893) );
  XNOR2_X1 U993 ( .A(G2678), .B(KEYINPUT42), .ZN(n892) );
  XNOR2_X1 U994 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(n895), .B(n894), .Z(G227) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n896), .B(KEYINPUT110), .ZN(n897) );
  NAND2_X1 U998 ( .A1(G319), .A2(n897), .ZN(n898) );
  NOR2_X1 U999 ( .A1(G401), .A2(n898), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n899) );
  XOR2_X1 U1001 ( .A(KEYINPUT49), .B(n899), .Z(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1004 ( .A(KEYINPUT59), .B(G1348), .ZN(n902) );
  XNOR2_X1 U1005 ( .A(n902), .B(G4), .ZN(n909) );
  XOR2_X1 U1006 ( .A(G1341), .B(G19), .Z(n905) );
  XNOR2_X1 U1007 ( .A(n903), .B(G20), .ZN(n904) );
  NAND2_X1 U1008 ( .A1(n905), .A2(n904), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(G6), .B(G1981), .ZN(n906) );
  NOR2_X1 U1010 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(n910), .B(KEYINPUT60), .ZN(n911) );
  XNOR2_X1 U1013 ( .A(n911), .B(KEYINPUT123), .ZN(n914) );
  XOR2_X1 U1014 ( .A(G1966), .B(G21), .Z(n912) );
  XNOR2_X1 U1015 ( .A(KEYINPUT124), .B(n912), .ZN(n913) );
  NAND2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n917) );
  XOR2_X1 U1017 ( .A(n915), .B(G5), .Z(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(KEYINPUT125), .B(n918), .ZN(n926) );
  XOR2_X1 U1020 ( .A(G1986), .B(G24), .Z(n922) );
  XNOR2_X1 U1021 ( .A(G1971), .B(G22), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(G23), .B(G1976), .ZN(n919) );
  NOR2_X1 U1023 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1025 ( .A(KEYINPUT126), .B(n923), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(KEYINPUT58), .B(n924), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1028 ( .A(KEYINPUT61), .B(n927), .Z(n928) );
  NOR2_X1 U1029 ( .A1(G16), .A2(n928), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT127), .B(n929), .ZN(n986) );
  XNOR2_X1 U1031 ( .A(KEYINPUT115), .B(G2090), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(n930), .B(G35), .ZN(n950) );
  XNOR2_X1 U1033 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n945) );
  XNOR2_X1 U1034 ( .A(n931), .B(G27), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(KEYINPUT116), .B(G32), .ZN(n933) );
  XNOR2_X1 U1036 ( .A(n933), .B(n932), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(n936), .B(KEYINPUT117), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(G1991), .B(G25), .ZN(n938) );
  XNOR2_X1 U1040 ( .A(G26), .B(G2067), .ZN(n937) );
  NOR2_X1 U1041 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1043 ( .A(G2072), .B(G33), .Z(n941) );
  NAND2_X1 U1044 ( .A1(G28), .A2(n941), .ZN(n942) );
  NOR2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(n945), .B(n944), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(G2084), .B(G34), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(KEYINPUT54), .B(n946), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n952) );
  XOR2_X1 U1051 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n951) );
  XNOR2_X1 U1052 ( .A(n952), .B(n951), .ZN(n953) );
  OR2_X1 U1053 ( .A1(G29), .A2(n953), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(G11), .A2(n954), .ZN(n984) );
  XOR2_X1 U1055 ( .A(KEYINPUT52), .B(KEYINPUT113), .Z(n979) );
  XOR2_X1 U1056 ( .A(G160), .B(G2084), .Z(n955) );
  NOR2_X1 U1057 ( .A1(n956), .A2(n955), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(KEYINPUT111), .B(n959), .ZN(n960) );
  NOR2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n968) );
  XOR2_X1 U1062 ( .A(G2090), .B(G162), .Z(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(n966), .B(KEYINPUT51), .ZN(n967) );
  NOR2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1066 ( .A(KEYINPUT112), .B(n969), .Z(n975) );
  XOR2_X1 U1067 ( .A(G2072), .B(n970), .Z(n972) );
  XOR2_X1 U1068 ( .A(G164), .B(G2078), .Z(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1070 ( .A(KEYINPUT50), .B(n973), .Z(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n979), .B(n978), .ZN(n980) );
  OR2_X1 U1074 ( .A1(KEYINPUT55), .A2(n980), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n981), .A2(G29), .ZN(n982) );
  XOR2_X1 U1076 ( .A(KEYINPUT114), .B(n982), .Z(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n1016) );
  XOR2_X1 U1079 ( .A(G16), .B(KEYINPUT56), .Z(n1014) );
  XOR2_X1 U1080 ( .A(n987), .B(G1341), .Z(n990) );
  XNOR2_X1 U1081 ( .A(n988), .B(G1956), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n1011) );
  XOR2_X1 U1083 ( .A(G168), .B(G1966), .Z(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1085 ( .A(KEYINPUT120), .B(n993), .Z(n994) );
  XNOR2_X1 U1086 ( .A(KEYINPUT57), .B(n994), .ZN(n1009) );
  INV_X1 U1087 ( .A(G1971), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(G166), .A2(n995), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1000), .B(G1348), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(G1961), .B(KEYINPUT121), .Z(n1001) );
  XNOR2_X1 U1093 ( .A(G301), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT122), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(n1017), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

