//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n617, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n467), .ZN(new_n468));
  XOR2_X1   g043(.A(new_n468), .B(KEYINPUT66), .Z(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(new_n466), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n473), .A2(G2105), .B1(G101), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n476), .B(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n464), .A2(new_n466), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n479), .A2(new_n467), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n467), .A2(G112), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n479), .A2(G2105), .A3(new_n481), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n479), .A2(new_n489), .A3(G2105), .A4(new_n481), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n486), .B1(new_n491), .B2(G124), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n464), .A3(new_n466), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n494), .A2(new_n464), .A3(new_n466), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n496), .A2(KEYINPUT71), .A3(KEYINPUT4), .A4(new_n498), .ZN(new_n502));
  XOR2_X1   g077(.A(KEYINPUT72), .B(KEYINPUT4), .Z(new_n503));
  OR2_X1    g078(.A1(new_n503), .A2(new_n495), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(G114), .A2(G2104), .ZN(new_n506));
  INV_X1    g081(.A(G126), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n471), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G2105), .B1(G102), .B2(new_n474), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT74), .B(G88), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(new_n517), .B1(G50), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT75), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT73), .A2(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT6), .ZN(new_n521));
  OR3_X1    g096(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n519), .B1(new_n518), .B2(new_n521), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n522), .A2(new_n529), .A3(new_n525), .A4(new_n526), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(G166));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n520), .B(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n516), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  INV_X1    g113(.A(G51), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT77), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n521), .A2(KEYINPUT77), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(new_n542), .A3(G543), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n536), .B(new_n538), .C1(new_n539), .C2(new_n543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(KEYINPUT78), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(KEYINPUT78), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G168));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n513), .A2(new_n515), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G651), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n533), .A2(new_n516), .ZN(new_n554));
  INV_X1    g129(.A(G52), .ZN(new_n555));
  OAI221_X1 g130(.A(new_n552), .B1(new_n553), .B2(new_n554), .C1(new_n543), .C2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  AOI22_X1  g132(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT79), .Z(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  INV_X1    g135(.A(new_n543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G43), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n521), .A2(new_n549), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G81), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n560), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT80), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT81), .ZN(G188));
  INV_X1    g149(.A(KEYINPUT82), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(KEYINPUT82), .A2(KEYINPUT9), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n561), .A2(G53), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n549), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n563), .A2(G91), .B1(new_n582), .B2(G651), .ZN(new_n583));
  INV_X1    g158(.A(G53), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n575), .B(new_n576), .C1(new_n543), .C2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n579), .A2(new_n583), .A3(new_n585), .ZN(G299));
  INV_X1    g161(.A(G168), .ZN(G286));
  INV_X1    g162(.A(G166), .ZN(G303));
  NAND4_X1  g163(.A1(new_n541), .A2(new_n542), .A3(G49), .A4(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n563), .A2(G87), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  NAND3_X1  g167(.A1(new_n533), .A2(G48), .A3(G543), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT83), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n595), .A2(new_n524), .B1(new_n554), .B2(new_n596), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n594), .A2(new_n597), .ZN(G305));
  AND2_X1   g173(.A1(new_n561), .A2(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n600), .A2(new_n524), .B1(new_n554), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n563), .A2(G92), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT10), .Z(new_n607));
  NAND2_X1  g182(.A1(new_n561), .A2(G54), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(new_n524), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G868), .ZN(G284));
  XOR2_X1   g188(.A(G284), .B(KEYINPUT84), .Z(G321));
  MUX2_X1   g189(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g190(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g191(.A(KEYINPUT85), .B(G559), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n612), .B1(G860), .B2(new_n618), .ZN(G148));
  NAND2_X1  g194(.A1(new_n612), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(KEYINPUT86), .B1(new_n467), .B2(G111), .ZN(new_n627));
  OR3_X1    g202(.A1(new_n467), .A2(KEYINPUT86), .A3(G111), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n625), .ZN(new_n629));
  NAND4_X1  g204(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G135), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n482), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n491), .B2(G123), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2096), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2100), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT88), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  XOR2_X1   g220(.A(G2443), .B(G2446), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT89), .B(KEYINPUT16), .Z(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G14), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT90), .Z(G401));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT17), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2084), .B(G2090), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT91), .ZN(new_n660));
  XOR2_X1   g235(.A(G2067), .B(G2678), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT92), .ZN(new_n663));
  INV_X1    g238(.A(new_n661), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n656), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  AOI21_X1  g241(.A(new_n660), .B1(new_n657), .B2(new_n664), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n656), .B2(new_n664), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT94), .ZN(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n674), .A2(new_n675), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(new_n679), .ZN(new_n683));
  OR3_X1    g258(.A1(new_n676), .A2(new_n682), .A3(new_n679), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT95), .B(G1981), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n689), .B(new_n692), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(KEYINPUT28), .ZN(new_n695));
  INV_X1    g270(.A(G26), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G29), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(G29), .ZN(new_n698));
  INV_X1    g273(.A(G140), .ZN(new_n699));
  OAI21_X1  g274(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n467), .A2(G116), .ZN(new_n701));
  OAI22_X1  g276(.A1(new_n482), .A2(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n491), .B2(G128), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT98), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n698), .B1(new_n705), .B2(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n697), .B1(new_n706), .B2(new_n695), .ZN(new_n707));
  INV_X1    g282(.A(G2067), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT106), .B(KEYINPUT30), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G28), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n474), .A2(G103), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT25), .Z(new_n714));
  INV_X1    g289(.A(G139), .ZN(new_n715));
  INV_X1    g290(.A(G127), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n471), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G115), .B2(G2104), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n714), .B1(new_n715), .B2(new_n482), .C1(new_n718), .C2(new_n467), .ZN(new_n719));
  MUX2_X1   g294(.A(G33), .B(new_n719), .S(G29), .Z(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(G2072), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n712), .B(new_n721), .C1(G29), .C2(new_n633), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n723), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT105), .B(G1966), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n709), .A2(new_n722), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G34), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT99), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(G34), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(new_n732), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT100), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n738), .B(new_n739), .C1(G160), .C2(G29), .ZN(new_n740));
  NOR2_X1   g315(.A1(G29), .A2(G35), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G162), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT108), .B(KEYINPUT29), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n740), .A2(G2084), .B1(new_n744), .B2(G2090), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n740), .A2(G2084), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT101), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n723), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n612), .B2(new_n723), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(G1348), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT101), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n740), .A2(new_n751), .A3(G2084), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n749), .A2(G1348), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n747), .A2(new_n750), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n729), .A2(G27), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G164), .B2(new_n729), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2078), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n728), .A2(new_n745), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n725), .A2(new_n726), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT107), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n744), .A2(G2090), .ZN(new_n761));
  INV_X1    g336(.A(G1961), .ZN(new_n762));
  NOR2_X1   g337(.A1(G171), .A2(new_n723), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G5), .B2(new_n723), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n761), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(G299), .A2(G16), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n723), .A2(KEYINPUT23), .A3(G20), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n769));
  INV_X1    g344(.A(G20), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(G16), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n758), .A2(new_n760), .A3(new_n766), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n723), .A2(G23), .ZN(new_n776));
  INV_X1    g351(.A(G288), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n723), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT33), .B(G1976), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT97), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n778), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G6), .A2(G16), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n594), .A2(new_n597), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G16), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT32), .B(G1981), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(G166), .A2(G16), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G16), .B2(G22), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n788), .A2(G1971), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(G1971), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n781), .B(new_n786), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT34), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n788), .B(G1971), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT34), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n793), .A2(new_n794), .A3(new_n781), .A4(new_n786), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n723), .A2(G24), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n603), .B2(new_n723), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(new_n686), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n729), .A2(G25), .ZN(new_n799));
  INV_X1    g374(.A(new_n482), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n491), .A2(G119), .B1(G131), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(G95), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT96), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n729), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT35), .B(G1991), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n806), .B(new_n807), .Z(new_n808));
  NAND4_X1  g383(.A1(new_n792), .A2(new_n795), .A3(new_n798), .A4(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n729), .A2(G32), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n491), .A2(G129), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT102), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n491), .A2(KEYINPUT102), .A3(G129), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT104), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n800), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n819));
  NAND3_X1  g394(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT103), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT26), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT102), .B1(new_n491), .B2(G129), .ZN(new_n824));
  INV_X1    g399(.A(G129), .ZN(new_n825));
  AOI211_X1 g400(.A(new_n814), .B(new_n825), .C1(new_n488), .C2(new_n490), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n819), .B(new_n822), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT104), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n812), .B1(new_n830), .B2(new_n729), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT27), .B(G1996), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n775), .A2(new_n811), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(G16), .A2(G19), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n566), .B2(G16), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(G1341), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n720), .A2(G2072), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT31), .B(G11), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n834), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(G311));
  NAND2_X1  g416(.A1(new_n840), .A2(KEYINPUT109), .ZN(new_n842));
  INV_X1    g417(.A(new_n839), .ZN(new_n843));
  NOR4_X1   g418(.A1(new_n775), .A2(new_n811), .A3(new_n843), .A4(new_n833), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT109), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n837), .A4(new_n838), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(new_n846), .ZN(G150));
  AOI22_X1  g422(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n848), .A2(new_n524), .B1(new_n554), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n561), .B2(G55), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n612), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n851), .B(KEYINPUT110), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n565), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n851), .B(KEYINPUT110), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n566), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n854), .B1(new_n863), .B2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT111), .Z(G145));
  INV_X1    g440(.A(KEYINPUT114), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n703), .B(KEYINPUT98), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n823), .A2(new_n828), .A3(G164), .ZN(new_n868));
  AOI21_X1  g443(.A(G164), .B1(new_n823), .B2(new_n828), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n829), .A2(new_n510), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n823), .A2(new_n828), .A3(G164), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n705), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT112), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n719), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n870), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n870), .B2(new_n873), .ZN(new_n878));
  INV_X1    g453(.A(new_n636), .ZN(new_n879));
  OR2_X1    g454(.A1(G106), .A2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n880), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n881));
  INV_X1    g456(.A(G142), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n482), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n491), .B2(G130), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n805), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n801), .A2(new_n804), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n884), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT113), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n886), .B2(new_n888), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n879), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n636), .A3(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n877), .A2(new_n878), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n893), .A2(new_n895), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n868), .A2(new_n869), .A3(new_n867), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n705), .B1(new_n871), .B2(new_n872), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n875), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n870), .A2(new_n873), .A3(new_n876), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n866), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(G160), .B(new_n633), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(G162), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n896), .B1(new_n877), .B2(new_n878), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT114), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n901), .A2(new_n898), .A3(new_n902), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT115), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n913), .B1(new_n912), .B2(new_n866), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n917), .B2(new_n908), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT115), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n914), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(new_n920), .A3(KEYINPUT40), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT40), .B1(new_n916), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(G395));
  XNOR2_X1  g498(.A(new_n862), .B(new_n620), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n611), .B(G299), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT116), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n925), .B(KEYINPUT41), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n931));
  XNOR2_X1  g506(.A(G166), .B(G288), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(G290), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(new_n783), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n927), .A2(new_n935), .A3(new_n929), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n931), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n931), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(G868), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(G868), .B2(new_n851), .ZN(G295));
  OAI21_X1  g515(.A(new_n939), .B1(G868), .B2(new_n851), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT117), .ZN(new_n942));
  XNOR2_X1  g517(.A(G168), .B(G171), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n943), .A2(new_n862), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n862), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n928), .ZN(new_n947));
  INV_X1    g522(.A(new_n925), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n933), .B(G305), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n942), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G37), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n934), .A2(KEYINPUT117), .A3(new_n949), .A4(new_n947), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT118), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT44), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n956), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n958), .B(new_n961), .ZN(G397));
  AOI21_X1  g537(.A(G1384), .B1(new_n505), .B2(new_n509), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT45), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n469), .A2(G40), .A3(new_n475), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT119), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n966), .B(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n830), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n705), .B(new_n708), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n829), .A2(G1996), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n887), .A2(new_n807), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n807), .B2(new_n887), .ZN(new_n977));
  NAND2_X1  g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(G290), .A2(G1986), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n969), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT61), .ZN(new_n984));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n510), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n963), .A2(KEYINPUT45), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT56), .B(G2072), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n988), .A2(new_n965), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n992));
  XNOR2_X1  g567(.A(G299), .B(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n963), .A2(new_n994), .ZN(new_n995));
  AOI211_X1 g570(.A(KEYINPUT50), .B(G1384), .C1(new_n505), .C2(new_n509), .ZN(new_n996));
  INV_X1    g571(.A(new_n965), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n991), .B(new_n993), .C1(new_n998), .C2(G1956), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n963), .A2(new_n994), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n965), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n773), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n993), .B1(new_n1004), .B2(new_n991), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n984), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT123), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT123), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(new_n984), .C1(new_n1000), .C2(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n988), .A2(new_n965), .A3(new_n989), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n963), .A2(new_n965), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT58), .B(G1341), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n1011), .A2(G1996), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n566), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT59), .ZN(new_n1017));
  INV_X1    g592(.A(G1348), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1003), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1012), .A2(G2067), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n611), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n612), .B(new_n1020), .C1(new_n1003), .C2(new_n1018), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT60), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n993), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n995), .A2(new_n996), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1956), .B1(new_n1026), .B2(new_n965), .ZN(new_n1027));
  INV_X1    g602(.A(new_n991), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT61), .A3(new_n999), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n611), .A2(KEYINPUT60), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1019), .A2(new_n1021), .A3(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1024), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1010), .A2(new_n1017), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT124), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1005), .B1(new_n999), .B2(new_n1022), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1035), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1038));
  AOI211_X1 g613(.A(new_n987), .B(G1384), .C1(new_n505), .C2(new_n509), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n964), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n726), .B1(new_n1040), .B2(new_n965), .ZN(new_n1041));
  NOR4_X1   g616(.A1(new_n995), .A2(new_n996), .A3(G2084), .A4(new_n997), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(KEYINPUT125), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G286), .A2(G8), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(KEYINPUT125), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n964), .A2(new_n1039), .A3(new_n997), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1050), .A2(new_n726), .B1(new_n1003), .B2(G2084), .ZN(new_n1051));
  OAI211_X1 g626(.A(G8), .B(new_n1045), .C1(new_n1051), .C2(G286), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1043), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G286), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G305), .A2(G1981), .ZN(new_n1057));
  OR3_X1    g632(.A1(new_n594), .A2(G1981), .A3(new_n597), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT49), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1013), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1057), .A2(KEYINPUT49), .A3(new_n1058), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n777), .A2(G1976), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1012), .A2(G8), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n1069));
  INV_X1    g644(.A(G1976), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G288), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1012), .A2(G8), .A3(new_n1066), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1071), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1073), .A2(KEYINPUT52), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT121), .B1(new_n1073), .B2(KEYINPUT52), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1065), .B(new_n1072), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1050), .A2(G1971), .B1(new_n1003), .B2(G2090), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G8), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n528), .A2(KEYINPUT55), .A3(G8), .A4(new_n530), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(G166), .B2(new_n1062), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1080), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1079), .A3(G8), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1078), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  OR3_X1    g667(.A1(new_n1011), .A2(new_n1092), .A3(G2078), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1003), .A2(new_n762), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1011), .B2(G2078), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1093), .A2(G301), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1056), .B(new_n1091), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1037), .A2(new_n1038), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1056), .A2(KEYINPUT62), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1097), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1053), .A2(new_n1106), .A3(new_n1055), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1104), .A2(new_n1091), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1091), .A2(G168), .A3(new_n1054), .A4(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1078), .A2(new_n1089), .A3(new_n1054), .A4(new_n1090), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1109), .B(new_n1110), .C1(new_n1113), .C2(G286), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1090), .A2(new_n1077), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1065), .A2(new_n1070), .A3(new_n777), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1058), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1116), .B1(new_n1063), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1108), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n983), .B1(new_n1103), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT46), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n969), .B2(G1996), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n972), .A2(new_n830), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n968), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n968), .A2(KEYINPUT46), .A3(new_n970), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT126), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT47), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n977), .A2(new_n969), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n968), .A2(new_n980), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT48), .ZN(new_n1132));
  INV_X1    g707(.A(new_n974), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n1133), .A2(new_n975), .B1(G2067), .B2(new_n705), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1130), .A2(new_n1132), .B1(new_n968), .B2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1121), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1102), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1108), .A2(new_n1119), .A3(new_n1115), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n982), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT127), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1138), .A2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g723(.A(new_n919), .B1(new_n918), .B2(new_n914), .ZN(new_n1150));
  AND4_X1   g724(.A1(new_n919), .A2(new_n909), .A3(new_n910), .A4(new_n914), .ZN(new_n1151));
  OAI211_X1 g725(.A(new_n671), .B(new_n693), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g726(.A(G401), .ZN(new_n1153));
  NAND3_X1  g727(.A1(new_n961), .A2(G319), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1154), .ZN(G308));
  AOI21_X1  g729(.A(G227), .B1(new_n916), .B2(new_n920), .ZN(new_n1156));
  AOI211_X1 g730(.A(new_n461), .B(G401), .C1(new_n960), .C2(new_n956), .ZN(new_n1157));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n693), .A3(new_n1157), .ZN(G225));
endmodule


