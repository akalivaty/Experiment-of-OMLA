//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  OR2_X1    g001(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n204));
  AOI21_X1  g003(.A(G36gat), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  AND3_X1   g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  OR3_X1    g006(.A1(new_n205), .A2(KEYINPUT15), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT15), .B1(new_n205), .B2(new_n207), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n209), .B2(new_n210), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT17), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(G1gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216));
  AOI21_X1  g015(.A(G8gat), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT16), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n214), .B1(new_n218), .B2(G1gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n217), .B(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n213), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n221), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n212), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n202), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n222), .A2(KEYINPUT18), .A3(new_n226), .A4(new_n224), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n221), .B(new_n212), .Z(new_n230));
  XOR2_X1   g029(.A(new_n226), .B(KEYINPUT13), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G113gat), .B(G141gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(G169gat), .B(G197gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT12), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n239), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G78gat), .B(G106gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G22gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(G197gat), .A2(G204gat), .ZN(new_n247));
  AND2_X1   g046(.A1(G197gat), .A2(G204gat), .ZN(new_n248));
  AND2_X1   g047(.A1(G211gat), .A2(G218gat), .ZN(new_n249));
  OAI22_X1  g048(.A1(new_n247), .A2(new_n248), .B1(new_n249), .B2(KEYINPUT22), .ZN(new_n250));
  XOR2_X1   g049(.A(G211gat), .B(G218gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT74), .ZN(new_n253));
  NAND2_X1  g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT2), .ZN(new_n255));
  INV_X1    g054(.A(G141gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G148gat), .ZN(new_n257));
  INV_X1    g056(.A(G148gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(G141gat), .ZN(new_n259));
  OAI211_X1 g058(.A(KEYINPUT79), .B(new_n255), .C1(new_n257), .C2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G155gat), .B(G162gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT79), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n258), .A2(G141gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n256), .A2(G148gat), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(new_n261), .A3(new_n255), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT3), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n263), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT29), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n263), .A2(new_n268), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT3), .B1(new_n252), .B2(new_n271), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n273), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(G228gat), .A3(G233gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n252), .A2(KEYINPUT83), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n250), .A2(KEYINPUT83), .A3(new_n251), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n271), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n269), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n274), .ZN(new_n283));
  NAND2_X1  g082(.A1(G228gat), .A2(G233gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n273), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT31), .B(G50gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n278), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(new_n278), .B2(new_n285), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n246), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(new_n245), .A3(new_n288), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G71gat), .B(G99gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT72), .ZN(new_n296));
  INV_X1    g095(.A(G15gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G43gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT27), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(G183gat), .ZN(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(G183gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(KEYINPUT65), .A3(KEYINPUT27), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n304), .ZN(new_n311));
  NAND2_X1  g110(.A1(KEYINPUT66), .A2(KEYINPUT27), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n307), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n302), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT67), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n316), .B(new_n302), .C1(new_n309), .C2(new_n313), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT27), .B(G183gat), .Z(new_n318));
  NOR3_X1   g117(.A1(new_n318), .A2(new_n302), .A3(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n315), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n324), .A2(KEYINPUT26), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n331));
  NOR2_X1   g130(.A1(G127gat), .A2(G134gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G113gat), .B(G120gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(KEYINPUT1), .ZN(new_n335));
  NAND2_X1  g134(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n338));
  OAI21_X1  g137(.A(G127gat), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n342));
  NAND2_X1  g141(.A1(G127gat), .A2(G134gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n344), .B2(new_n332), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT69), .B1(new_n346), .B2(G120gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT69), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(G113gat), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT70), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G113gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n354), .A3(G120gat), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n345), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n331), .B1(new_n341), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT1), .B1(new_n333), .B2(new_n343), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n352), .A2(new_n354), .A3(G120gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n347), .A2(new_n350), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n339), .B(new_n333), .C1(KEYINPUT1), .C2(new_n334), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT71), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT64), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n364), .A2(new_n365), .B1(G169gat), .B2(G176gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(G169gat), .B2(G176gat), .ZN(new_n372));
  INV_X1    g171(.A(G169gat), .ZN(new_n373));
  INV_X1    g172(.A(G176gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT23), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n368), .A2(new_n370), .A3(new_n372), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n307), .A2(new_n306), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n377), .A2(KEYINPUT24), .A3(new_n326), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n367), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n365), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n370), .A2(new_n380), .A3(new_n322), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n375), .A2(new_n372), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(KEYINPUT24), .A3(new_n326), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n366), .A4(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n330), .A2(new_n357), .A3(new_n363), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n357), .A2(new_n363), .ZN(new_n388));
  INV_X1    g187(.A(new_n329), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n319), .B1(new_n314), .B2(KEYINPUT67), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n317), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n388), .B1(new_n391), .B2(new_n385), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n301), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n387), .A2(new_n392), .A3(new_n394), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT34), .B1(new_n395), .B2(KEYINPUT73), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n387), .A2(new_n392), .A3(new_n394), .A4(new_n400), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n394), .B1(new_n387), .B2(new_n392), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n300), .B1(new_n406), .B2(KEYINPUT33), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n403), .A3(new_n402), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n396), .A2(KEYINPUT32), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n405), .B2(new_n408), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n294), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n271), .B1(new_n391), .B2(new_n385), .ZN(new_n415));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n416), .B(KEYINPUT75), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n330), .A2(new_n386), .ZN(new_n419));
  INV_X1    g218(.A(new_n416), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n415), .A2(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n253), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT76), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n385), .B1(new_n321), .B2(new_n329), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n418), .B1(new_n424), .B2(KEYINPUT29), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(new_n420), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n253), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n415), .A2(new_n416), .B1(new_n419), .B2(new_n417), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT77), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n431), .A3(new_n422), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n416), .B1(new_n424), .B2(KEYINPUT29), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n417), .B1(new_n391), .B2(new_n385), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n422), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT77), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n423), .A2(new_n429), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT5), .ZN(new_n443));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT80), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n361), .A2(new_n362), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(new_n274), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n361), .A2(new_n362), .B1(new_n263), .B2(new_n268), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n274), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n361), .A2(new_n362), .A3(new_n263), .A4(new_n268), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n446), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n443), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n357), .A2(KEYINPUT4), .A3(new_n275), .A4(new_n363), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n447), .A3(new_n270), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n458), .A2(new_n460), .A3(new_n462), .A4(new_n445), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n453), .A2(new_n459), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n357), .A2(new_n275), .A3(new_n363), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(new_n459), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n462), .A2(new_n443), .A3(new_n445), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n457), .A2(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G1gat), .B(G29gat), .Z(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G57gat), .B(G85gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT6), .B1(new_n468), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n456), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n455), .B1(new_n454), .B2(new_n446), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT5), .B(new_n463), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n467), .A2(new_n466), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n473), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(KEYINPUT6), .A3(new_n473), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n441), .A2(new_n442), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n428), .B1(new_n427), .B2(new_n253), .ZN(new_n486));
  AOI211_X1 g285(.A(KEYINPUT76), .B(new_n422), .C1(new_n425), .C2(new_n426), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n431), .B1(new_n430), .B2(new_n422), .ZN(new_n488));
  AND4_X1   g287(.A1(new_n431), .A2(new_n433), .A3(new_n422), .A4(new_n434), .ZN(new_n489));
  OAI22_X1  g288(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n440), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n423), .A2(new_n429), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n432), .A2(new_n436), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT30), .A4(new_n440), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n485), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n492), .A2(new_n485), .A3(new_n495), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n414), .B(new_n484), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n492), .A2(new_n495), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT30), .B1(new_n437), .B2(new_n440), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n414), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT85), .B1(new_n468), .B2(new_n474), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n480), .A2(new_n505), .A3(new_n473), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n475), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT35), .B1(new_n507), .B2(new_n483), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n499), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n484), .B1(new_n497), .B2(new_n496), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n291), .A2(new_n293), .A3(KEYINPUT84), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT84), .B1(new_n291), .B2(new_n293), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n465), .A2(new_n459), .ZN(new_n516));
  INV_X1    g315(.A(new_n464), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n462), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT39), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n446), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n474), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT39), .B1(new_n454), .B2(new_n446), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n518), .B2(new_n446), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n521), .A2(KEYINPUT40), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT40), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n445), .B1(new_n466), .B2(new_n462), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n473), .B1(new_n526), .B2(new_n519), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n518), .A2(new_n446), .ZN(new_n528));
  INV_X1    g327(.A(new_n522), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n525), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n504), .A2(new_n506), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n500), .B2(new_n501), .ZN(new_n535));
  INV_X1    g334(.A(new_n294), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(new_n430), .B2(new_n253), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n427), .A2(new_n422), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT38), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n491), .B(new_n540), .C1(new_n490), .C2(KEYINPUT37), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n541), .A2(new_n483), .A3(new_n441), .A4(new_n507), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT38), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n440), .B1(new_n437), .B2(new_n537), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n490), .A2(KEYINPUT37), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n535), .B(new_n536), .C1(new_n542), .C2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n412), .B2(new_n413), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n405), .A2(new_n408), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n409), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(KEYINPUT36), .A3(new_n411), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n515), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n243), .B1(new_n510), .B2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G155gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(KEYINPUT89), .A2(G57gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(G64gat), .ZN(new_n567));
  INV_X1    g366(.A(G64gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(KEYINPUT89), .A3(G57gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n567), .A2(new_n569), .B1(new_n563), .B2(new_n562), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(KEYINPUT91), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n572));
  INV_X1    g371(.A(new_n570), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(new_n564), .ZN(new_n574));
  XOR2_X1   g373(.A(G71gat), .B(G78gat), .Z(new_n575));
  XNOR2_X1  g374(.A(G57gat), .B(G64gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT88), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n563), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n577), .B2(new_n576), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n571), .A2(new_n574), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(KEYINPUT21), .ZN(new_n581));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n581), .B(new_n582), .Z(new_n583));
  INV_X1    g382(.A(G127gat), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n223), .B1(KEYINPUT21), .B2(new_n580), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n584), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n587), .B1(new_n585), .B2(new_n588), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n560), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n589), .A3(new_n559), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT92), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n599));
  XOR2_X1   g398(.A(G134gat), .B(G162gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT95), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n604), .B(new_n605), .Z(new_n606));
  XOR2_X1   g405(.A(G99gat), .B(G106gat), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n606), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT94), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n607), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n613), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n213), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n615), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n621), .A2(new_n212), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G190gat), .B(G218gat), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n603), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n601), .A2(KEYINPUT95), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n625), .A2(new_n627), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n595), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n608), .B1(new_n606), .B2(new_n612), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n614), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n580), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n636), .B(new_n637), .C1(new_n621), .C2(new_n580), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n580), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT98), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n636), .B1(new_n621), .B2(new_n580), .ZN(new_n644));
  INV_X1    g443(.A(new_n641), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n640), .A2(new_n647), .A3(new_n641), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n643), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n646), .B2(KEYINPUT97), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(KEYINPUT97), .B2(new_n646), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n645), .B1(new_n640), .B2(KEYINPUT96), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(KEYINPUT96), .B2(new_n640), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n633), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n555), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n482), .A2(new_n483), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  INV_X1    g465(.A(new_n502), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(G8gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(KEYINPUT42), .B2(new_n671), .ZN(G1325gat));
  NAND2_X1  g472(.A1(new_n553), .A2(KEYINPUT99), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n549), .A2(new_n552), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n297), .B1(new_n662), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n412), .A2(new_n413), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(G15gat), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n678), .B1(new_n662), .B2(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT100), .Z(G1326gat));
  NAND2_X1  g482(.A1(new_n662), .A2(new_n514), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  AOI22_X1  g486(.A1(KEYINPUT35), .A2(new_n498), .B1(new_n503), .B2(new_n508), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n515), .A2(new_n547), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT102), .B1(new_n689), .B2(new_n677), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n549), .A2(new_n552), .A3(new_n675), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n675), .B1(new_n549), .B2(new_n552), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n515), .A4(new_n547), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n688), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n687), .B1(new_n696), .B2(new_n632), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n510), .A2(new_n554), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(KEYINPUT44), .A3(new_n631), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n243), .A2(new_n595), .A3(new_n660), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G29gat), .B1(new_n702), .B2(new_n663), .ZN(new_n703));
  INV_X1    g502(.A(new_n595), .ZN(new_n704));
  INV_X1    g503(.A(new_n660), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n631), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT101), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n555), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n206), .A3(new_n664), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n703), .A2(KEYINPUT103), .A3(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1328gat));
  OAI21_X1  g515(.A(G36gat), .B1(new_n702), .B2(new_n502), .ZN(new_n717));
  AOI21_X1  g516(.A(G36gat), .B1(KEYINPUT104), .B2(KEYINPUT46), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n709), .A2(new_n667), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(new_n721), .ZN(G1329gat));
  NAND4_X1  g521(.A1(new_n697), .A2(new_n677), .A3(new_n699), .A4(new_n701), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n299), .B1(new_n723), .B2(KEYINPUT105), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(KEYINPUT105), .B2(new_n723), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n299), .A3(new_n679), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(KEYINPUT47), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(G43gat), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n726), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(KEYINPUT47), .B2(new_n729), .ZN(G1330gat));
  OAI21_X1  g529(.A(G50gat), .B1(new_n702), .B2(new_n536), .ZN(new_n731));
  INV_X1    g530(.A(new_n514), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n708), .A2(G50gat), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n700), .A2(new_n514), .A3(new_n701), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n736), .B2(G50gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(KEYINPUT48), .B2(new_n737), .ZN(G1331gat));
  INV_X1    g537(.A(new_n696), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n633), .A2(new_n242), .A3(new_n705), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n664), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT106), .B(G57gat), .Z(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1332gat));
  INV_X1    g543(.A(new_n741), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n502), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  AND2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n746), .B2(new_n747), .ZN(G1333gat));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n745), .B2(new_n680), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n741), .A2(G71gat), .A3(new_n677), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(KEYINPUT107), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(KEYINPUT107), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT50), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n758), .B(new_n752), .C1(new_n754), .C2(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1334gat));
  NAND2_X1  g559(.A1(new_n741), .A2(new_n514), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g561(.A1(new_n595), .A2(new_n242), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n705), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n700), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n663), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n690), .A2(new_n695), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n632), .B1(new_n768), .B2(new_n510), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT51), .B1(new_n769), .B2(new_n763), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NOR4_X1   g570(.A1(new_n696), .A2(new_n771), .A3(new_n632), .A4(new_n764), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n773), .A2(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(KEYINPUT108), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n660), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n664), .A2(new_n610), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n767), .B1(new_n776), .B2(new_n777), .ZN(G1336gat));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n769), .A2(new_n763), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n771), .ZN(new_n783));
  INV_X1    g582(.A(new_n772), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n502), .A2(new_n705), .A3(G92gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT109), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n781), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n779), .A2(new_n780), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n700), .A2(new_n667), .A3(new_n765), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G92gat), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n789), .B1(new_n788), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n766), .B2(new_n693), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n680), .A2(G99gat), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n776), .B2(new_n796), .ZN(G1338gat));
  NOR3_X1   g596(.A1(new_n536), .A2(new_n705), .A3(G106gat), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n770), .B2(new_n772), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n697), .A2(new_n514), .A3(new_n699), .A4(new_n765), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G106gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT111), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n805), .A3(G106gat), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT112), .B(new_n798), .C1(new_n770), .C2(new_n772), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n801), .A2(new_n804), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT53), .ZN(new_n809));
  OAI21_X1  g608(.A(G106gat), .B1(new_n766), .B2(new_n536), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n811), .A3(new_n799), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n812), .ZN(G1339gat));
  NOR3_X1   g612(.A1(new_n633), .A2(new_n242), .A3(new_n660), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n638), .A2(new_n645), .A3(new_n639), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n647), .B1(new_n640), .B2(new_n641), .ZN(new_n818));
  AOI211_X1 g617(.A(KEYINPUT98), .B(new_n645), .C1(new_n638), .C2(new_n639), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n820), .A2(new_n821), .A3(new_n653), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n820), .B2(new_n653), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n816), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT55), .B(new_n816), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n233), .A2(new_n239), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n230), .A2(new_n231), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n225), .A2(new_n227), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(KEYINPUT114), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n225), .A2(new_n832), .A3(new_n227), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n238), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n826), .A2(new_n659), .A3(new_n827), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n595), .B1(new_n836), .B2(new_n631), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n631), .B1(new_n835), .B2(new_n660), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n653), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT113), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n821), .A3(new_n653), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n242), .B1(new_n843), .B2(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n659), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n814), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n514), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n848), .A2(new_n664), .A3(new_n502), .A4(new_n679), .ZN(new_n849));
  OAI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n243), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n847), .A2(new_n663), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n503), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n242), .A2(new_n352), .A3(new_n354), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n849), .B2(new_n705), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n660), .A2(new_n349), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT115), .Z(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n852), .B2(new_n857), .ZN(G1341gat));
  INV_X1    g657(.A(new_n852), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n584), .A3(new_n595), .ZN(new_n860));
  OAI21_X1  g659(.A(G127gat), .B1(new_n849), .B2(new_n704), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1342gat));
  OR4_X1    g661(.A1(new_n338), .A2(new_n852), .A3(new_n337), .A4(new_n632), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n849), .B2(new_n632), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n677), .A2(new_n663), .A3(new_n667), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT116), .B(new_n870), .C1(new_n847), .C2(new_n536), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n835), .B1(new_n843), .B2(KEYINPUT55), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n631), .B1(new_n872), .B2(new_n845), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n846), .A2(new_n873), .A3(new_n704), .ZN(new_n874));
  INV_X1    g673(.A(new_n814), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(KEYINPUT57), .A3(new_n514), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n294), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT116), .B1(new_n879), .B2(new_n870), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n242), .B(new_n869), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n868), .B1(new_n881), .B2(G141gat), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n677), .A2(new_n536), .A3(new_n667), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n851), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(G141gat), .A3(new_n243), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n881), .B2(G141gat), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n882), .A2(new_n886), .A3(KEYINPUT58), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  AOI221_X4 g687(.A(new_n885), .B1(new_n868), .B2(new_n888), .C1(new_n881), .C2(G141gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n887), .A2(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n879), .A2(KEYINPUT57), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n870), .A3(new_n514), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n892), .A2(new_n660), .A3(new_n869), .A4(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n891), .B1(new_n894), .B2(G148gat), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n660), .B(new_n869), .C1(new_n878), .C2(new_n880), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n258), .A2(KEYINPUT59), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n851), .A2(new_n258), .A3(new_n660), .A4(new_n883), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT118), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n896), .A2(new_n897), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n902), .B(new_n899), .C1(new_n903), .C2(new_n895), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1345gat));
  OAI21_X1  g704(.A(new_n869), .B1(new_n878), .B2(new_n880), .ZN(new_n906));
  OAI21_X1  g705(.A(G155gat), .B1(new_n906), .B2(new_n704), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n704), .A2(G155gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n884), .B2(new_n908), .ZN(G1346gat));
  INV_X1    g708(.A(G162gat), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n906), .A2(new_n910), .A3(new_n632), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n851), .A2(new_n631), .A3(new_n883), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(G1347gat));
  NAND2_X1  g712(.A1(new_n667), .A2(new_n663), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n680), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n848), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(new_n373), .A3(new_n243), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n876), .A2(new_n663), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n502), .B1(new_n918), .B2(KEYINPUT119), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n664), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n414), .A3(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n919), .A2(KEYINPUT120), .A3(new_n920), .A4(new_n414), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n242), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n917), .B1(new_n925), .B2(new_n373), .ZN(G1348gat));
  NAND4_X1  g725(.A1(new_n923), .A2(new_n374), .A3(new_n660), .A4(new_n924), .ZN(new_n927));
  OAI21_X1  g726(.A(G176gat), .B1(new_n916), .B2(new_n705), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(KEYINPUT121), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n848), .A2(new_n595), .A3(new_n915), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n307), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n848), .A2(KEYINPUT122), .A3(new_n595), .A4(new_n915), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n704), .A2(new_n318), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n938), .B(new_n939), .C1(new_n921), .C2(new_n940), .ZN(new_n941));
  OR2_X1    g740(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n941), .B(new_n942), .ZN(G1350gat));
  NAND4_X1  g742(.A1(new_n923), .A2(new_n306), .A3(new_n631), .A4(new_n924), .ZN(new_n944));
  OAI21_X1  g743(.A(G190gat), .B1(new_n916), .B2(new_n632), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1351gat));
  NOR2_X1   g746(.A1(new_n677), .A2(new_n536), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n919), .A2(new_n948), .A3(new_n920), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n919), .A2(new_n951), .A3(new_n920), .A4(new_n948), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n243), .A2(G197gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n892), .A2(new_n893), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n677), .A2(new_n914), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n242), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G197gat), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n954), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n955), .B1(new_n954), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(G1352gat));
  NOR3_X1   g761(.A1(new_n949), .A2(G204gat), .A3(new_n705), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n956), .A2(new_n957), .ZN(new_n967));
  OAI21_X1  g766(.A(G204gat), .B1(new_n967), .B2(new_n705), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(G1353gat));
  NAND3_X1  g768(.A1(new_n956), .A2(new_n595), .A3(new_n957), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n950), .A2(new_n952), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n704), .A2(G211gat), .ZN(new_n974));
  OAI22_X1  g773(.A1(new_n971), .A2(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  INV_X1    g774(.A(new_n967), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n631), .A2(G218gat), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT127), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n979), .B1(new_n976), .B2(KEYINPUT126), .ZN(new_n980));
  INV_X1    g779(.A(G218gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n950), .A2(new_n631), .A3(new_n952), .ZN(new_n982));
  AOI22_X1  g781(.A1(new_n977), .A2(new_n980), .B1(new_n981), .B2(new_n982), .ZN(G1355gat));
endmodule


