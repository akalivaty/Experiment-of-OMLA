

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n371, n372, n373, n375, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815;

  BUF_X1 U374 ( .A(n720), .Z(n356) );
  XNOR2_X1 U375 ( .A(n695), .B(n359), .ZN(n358) );
  INV_X1 U376 ( .A(KEYINPUT2), .ZN(n359) );
  XNOR2_X1 U377 ( .A(n354), .B(n353), .ZN(n423) );
  INV_X1 U378 ( .A(n663), .ZN(n353) );
  XOR2_X1 U379 ( .A(G116), .B(G107), .Z(n562) );
  XOR2_X1 U380 ( .A(G146), .B(G125), .Z(n534) );
  XNOR2_X1 U381 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n527) );
  XNOR2_X1 U382 ( .A(G140), .B(G110), .ZN(n430) );
  OR2_X2 U383 ( .A1(n693), .A2(n457), .ZN(n456) );
  XNOR2_X1 U384 ( .A(G119), .B(G128), .ZN(n431) );
  NOR2_X1 U385 ( .A1(n689), .A2(KEYINPUT2), .ZN(n690) );
  NOR2_X2 U386 ( .A1(n710), .A2(n814), .ZN(n354) );
  XNOR2_X2 U387 ( .A(n542), .B(n541), .ZN(n578) );
  XNOR2_X2 U388 ( .A(n355), .B(n623), .ZN(n737) );
  NAND2_X1 U389 ( .A1(n372), .A2(n362), .ZN(n355) );
  XNOR2_X2 U390 ( .A(n652), .B(KEYINPUT6), .ZN(n420) );
  XNOR2_X2 U391 ( .A(n790), .B(n538), .ZN(n731) );
  NAND2_X1 U392 ( .A1(n436), .A2(n366), .ZN(n361) );
  NOR2_X2 U393 ( .A1(n585), .A2(n584), .ZN(n371) );
  NAND2_X1 U394 ( .A1(n357), .A2(n373), .ZN(n372) );
  NAND2_X1 U395 ( .A1(n378), .A2(n377), .ZN(n357) );
  NOR2_X2 U396 ( .A1(G953), .A2(n788), .ZN(n789) );
  NAND2_X1 U397 ( .A1(n358), .A2(n785), .ZN(n787) );
  XNOR2_X2 U398 ( .A(n361), .B(n544), .ZN(n585) );
  XNOR2_X2 U399 ( .A(n371), .B(KEYINPUT0), .ZN(n607) );
  XNOR2_X2 U400 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X2 U401 ( .A(n356), .B(n721), .ZN(n722) );
  XNOR2_X2 U402 ( .A(n731), .B(n730), .ZN(n732) );
  NAND2_X1 U403 ( .A1(n375), .A2(n379), .ZN(n362) );
  NAND2_X1 U404 ( .A1(n661), .A2(n685), .ZN(n750) );
  XNOR2_X1 U405 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n533) );
  NAND2_X1 U406 ( .A1(G234), .A2(G237), .ZN(n499) );
  INV_X1 U407 ( .A(G237), .ZN(n539) );
  OR2_X1 U408 ( .A1(n720), .A2(n397), .ZN(n396) );
  INV_X2 U409 ( .A(G953), .ZN(n531) );
  AND2_X1 U410 ( .A1(n465), .A2(n414), .ZN(n363) );
  AND2_X1 U411 ( .A1(n465), .A2(n413), .ZN(n364) );
  AND2_X1 U412 ( .A1(n465), .A2(n697), .ZN(n365) );
  NOR2_X1 U413 ( .A1(n748), .A2(n622), .ZN(n375) );
  OR2_X1 U414 ( .A1(n676), .A2(n674), .ZN(n661) );
  NAND2_X2 U415 ( .A1(n399), .A2(n396), .ZN(n652) );
  AND2_X1 U416 ( .A1(n697), .A2(n367), .ZN(n413) );
  NAND2_X1 U417 ( .A1(n696), .A2(KEYINPUT2), .ZN(n697) );
  AND2_X1 U418 ( .A1(n672), .A2(n388), .ZN(n387) );
  NAND2_X1 U419 ( .A1(n744), .A2(n368), .ZN(n388) );
  NOR2_X2 U420 ( .A1(n649), .A2(n585), .ZN(n744) );
  XNOR2_X1 U421 ( .A(n681), .B(KEYINPUT110), .ZN(n813) );
  NOR2_X1 U422 ( .A1(n399), .A2(KEYINPUT30), .ZN(n393) );
  AND2_X1 U423 ( .A1(n395), .A2(n653), .ZN(n394) );
  NAND2_X1 U424 ( .A1(n396), .A2(n366), .ZN(n395) );
  NOR2_X1 U425 ( .A1(n725), .A2(G902), .ZN(n473) );
  NAND2_X1 U426 ( .A1(n367), .A2(n398), .ZN(n397) );
  INV_X1 U427 ( .A(KEYINPUT89), .ZN(n405) );
  INV_X1 U428 ( .A(KEYINPUT83), .ZN(n386) );
  INV_X1 U429 ( .A(KEYINPUT47), .ZN(n369) );
  INV_X1 U430 ( .A(KEYINPUT34), .ZN(n620) );
  NOR2_X2 U431 ( .A1(G953), .A2(G237), .ZN(n549) );
  INV_X1 U432 ( .A(KEYINPUT35), .ZN(n623) );
  INV_X1 U433 ( .A(G902), .ZN(n398) );
  INV_X1 U434 ( .A(KEYINPUT48), .ZN(n445) );
  BUF_X1 U435 ( .A(G475), .Z(n711) );
  INV_X1 U436 ( .A(KEYINPUT8), .ZN(n492) );
  XNOR2_X2 U437 ( .A(G146), .B(G125), .ZN(n433) );
  XNOR2_X1 U438 ( .A(G137), .B(G134), .ZN(n482) );
  AND2_X1 U439 ( .A1(n697), .A2(n711), .ZN(n412) );
  XNOR2_X1 U440 ( .A(n403), .B(n445), .ZN(n684) );
  XNOR2_X1 U441 ( .A(n380), .B(KEYINPUT31), .ZN(n634) );
  NAND2_X1 U442 ( .A1(n387), .A2(n385), .ZN(n407) );
  INV_X1 U443 ( .A(n769), .ZN(n381) );
  OR2_X1 U444 ( .A1(n671), .A2(n670), .ZN(n672) );
  AND2_X1 U445 ( .A1(n594), .A2(n595), .ZN(n410) );
  XNOR2_X1 U446 ( .A(n682), .B(n405), .ZN(n404) );
  XNOR2_X1 U447 ( .A(n813), .B(n386), .ZN(n385) );
  AND2_X1 U448 ( .A1(n628), .A2(n595), .ZN(n409) );
  NOR2_X1 U449 ( .A1(n619), .A2(n620), .ZN(n379) );
  INV_X1 U450 ( .A(n619), .ZN(n377) );
  INV_X1 U451 ( .A(n607), .ZN(n619) );
  XNOR2_X1 U452 ( .A(n408), .B(KEYINPUT107), .ZN(n616) );
  AND2_X1 U453 ( .A1(n750), .A2(n369), .ZN(n368) );
  AND2_X1 U454 ( .A1(n411), .A2(n620), .ZN(n373) );
  NAND2_X1 U455 ( .A1(n399), .A2(n390), .ZN(n389) );
  NOR2_X1 U456 ( .A1(n394), .A2(n393), .ZN(n392) );
  INV_X1 U457 ( .A(n622), .ZN(n411) );
  AND2_X1 U458 ( .A1(n396), .A2(n391), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n383), .B(n515), .ZN(n382) );
  XNOR2_X1 U460 ( .A(n432), .B(n428), .ZN(n725) );
  XNOR2_X1 U461 ( .A(n518), .B(n384), .ZN(n383) );
  NOR2_X1 U462 ( .A1(n651), .A2(n653), .ZN(n391) );
  XNOR2_X1 U463 ( .A(n526), .B(n525), .ZN(n790) );
  XNOR2_X1 U464 ( .A(n551), .B(n523), .ZN(n526) );
  XNOR2_X1 U465 ( .A(n498), .B(n497), .ZN(n505) );
  INV_X1 U466 ( .A(n651), .ZN(n366) );
  XNOR2_X1 U467 ( .A(n433), .B(KEYINPUT10), .ZN(n546) );
  NAND2_X1 U468 ( .A1(n719), .A2(G902), .ZN(n400) );
  XNOR2_X1 U469 ( .A(G134), .B(G122), .ZN(n558) );
  XNOR2_X1 U470 ( .A(G113), .B(KEYINPUT5), .ZN(n487) );
  XOR2_X1 U471 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n559) );
  XNOR2_X1 U472 ( .A(G131), .B(G116), .ZN(n488) );
  XOR2_X1 U473 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n497) );
  INV_X1 U474 ( .A(n719), .ZN(n367) );
  XOR2_X1 U475 ( .A(G110), .B(KEYINPUT16), .Z(n523) );
  XNOR2_X2 U476 ( .A(G104), .B(KEYINPUT96), .ZN(n516) );
  XNOR2_X2 U477 ( .A(G110), .B(G107), .ZN(n517) );
  XNOR2_X1 U478 ( .A(KEYINPUT84), .B(KEYINPUT23), .ZN(n494) );
  XNOR2_X1 U479 ( .A(KEYINPUT3), .B(G119), .ZN(n524) );
  XNOR2_X1 U480 ( .A(G137), .B(KEYINPUT24), .ZN(n495) );
  INV_X2 U481 ( .A(G140), .ZN(n513) );
  NOR2_X1 U482 ( .A1(n684), .A2(KEYINPUT87), .ZN(n441) );
  NAND2_X2 U483 ( .A1(n794), .A2(n805), .ZN(n694) );
  XNOR2_X2 U484 ( .A(n425), .B(n421), .ZN(n794) );
  NOR2_X2 U485 ( .A1(n438), .A2(n441), .ZN(n805) );
  INV_X1 U486 ( .A(n748), .ZN(n378) );
  NOR2_X1 U487 ( .A1(n739), .A2(n634), .ZN(n636) );
  NAND2_X1 U488 ( .A1(n381), .A2(n607), .ZN(n380) );
  NAND2_X1 U489 ( .A1(n698), .A2(n520), .ZN(n480) );
  XNOR2_X2 U490 ( .A(n519), .B(n382), .ZN(n698) );
  INV_X1 U491 ( .A(n514), .ZN(n384) );
  XNOR2_X2 U492 ( .A(n801), .B(n484), .ZN(n519) );
  XNOR2_X2 U493 ( .A(n530), .B(n483), .ZN(n801) );
  NAND2_X1 U494 ( .A1(n392), .A2(n389), .ZN(n656) );
  AND2_X2 U495 ( .A1(n401), .A2(n400), .ZN(n399) );
  NAND2_X1 U496 ( .A1(n720), .A2(n719), .ZN(n401) );
  NAND2_X1 U497 ( .A1(n402), .A2(n439), .ZN(n438) );
  NAND2_X1 U498 ( .A1(n684), .A2(n418), .ZN(n402) );
  NAND2_X1 U499 ( .A1(n447), .A2(n423), .ZN(n403) );
  NAND2_X1 U500 ( .A1(n406), .A2(n404), .ZN(n448) );
  NAND2_X1 U501 ( .A1(n449), .A2(n627), .ZN(n682) );
  XNOR2_X1 U502 ( .A(n407), .B(KEYINPUT75), .ZN(n406) );
  INV_X1 U503 ( .A(n652), .ZN(n602) );
  NAND2_X1 U504 ( .A1(n420), .A2(n417), .ZN(n408) );
  NAND2_X1 U505 ( .A1(n594), .A2(n409), .ZN(n630) );
  NAND2_X1 U506 ( .A1(n410), .A2(n592), .ZN(n631) );
  AND2_X1 U507 ( .A1(n465), .A2(n412), .ZN(n715) );
  AND2_X1 U508 ( .A1(n697), .A2(G210), .ZN(n414) );
  NAND2_X1 U509 ( .A1(n437), .A2(n521), .ZN(n649) );
  NOR2_X2 U510 ( .A1(n416), .A2(n463), .ZN(n462) );
  NOR2_X2 U511 ( .A1(n415), .A2(KEYINPUT64), .ZN(n458) );
  NOR2_X1 U512 ( .A1(n693), .A2(n692), .ZN(n415) );
  NOR2_X1 U513 ( .A1(n689), .A2(KEYINPUT2), .ZN(n416) );
  NOR2_X2 U514 ( .A1(n694), .A2(KEYINPUT85), .ZN(n689) );
  XNOR2_X1 U515 ( .A(n448), .B(KEYINPUT71), .ZN(n447) );
  NAND2_X1 U516 ( .A1(KEYINPUT85), .A2(KEYINPUT64), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n683), .A2(KEYINPUT87), .ZN(n440) );
  NAND2_X1 U518 ( .A1(n477), .A2(n398), .ZN(n476) );
  XNOR2_X1 U519 ( .A(n473), .B(n471), .ZN(n426) );
  XNOR2_X1 U520 ( .A(n472), .B(KEYINPUT25), .ZN(n471) );
  NAND2_X1 U521 ( .A1(n505), .A2(G217), .ZN(n472) );
  INV_X1 U522 ( .A(n426), .ZN(n595) );
  XOR2_X1 U523 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n548) );
  XNOR2_X1 U524 ( .A(G143), .B(KEYINPUT11), .ZN(n547) );
  NAND2_X1 U525 ( .A1(n464), .A2(KEYINPUT64), .ZN(n463) );
  INV_X1 U526 ( .A(KEYINPUT33), .ZN(n452) );
  NOR2_X1 U527 ( .A1(n815), .A2(n440), .ZN(n439) );
  INV_X1 U528 ( .A(KEYINPUT41), .ZN(n647) );
  INV_X1 U529 ( .A(n578), .ZN(n436) );
  XNOR2_X1 U530 ( .A(n496), .B(n429), .ZN(n428) );
  XNOR2_X1 U531 ( .A(n434), .B(n546), .ZN(n432) );
  XNOR2_X1 U532 ( .A(n431), .B(n430), .ZN(n429) );
  XOR2_X1 U533 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n566) );
  XNOR2_X1 U534 ( .A(n451), .B(n450), .ZN(n449) );
  INV_X1 U535 ( .A(KEYINPUT36), .ZN(n450) );
  XNOR2_X1 U536 ( .A(n630), .B(n629), .ZN(n709) );
  AND2_X1 U537 ( .A1(n595), .A2(n419), .ZN(n417) );
  AND2_X1 U538 ( .A1(n683), .A2(KEYINPUT87), .ZN(n418) );
  AND2_X1 U539 ( .A1(n673), .A2(n764), .ZN(n419) );
  INV_X1 U540 ( .A(KEYINPUT1), .ZN(n470) );
  XNOR2_X1 U541 ( .A(KEYINPUT86), .B(KEYINPUT45), .ZN(n421) );
  XNOR2_X1 U542 ( .A(n618), .B(n454), .ZN(n444) );
  XNOR2_X2 U543 ( .A(n422), .B(KEYINPUT76), .ZN(n618) );
  NAND2_X1 U544 ( .A1(n573), .A2(n654), .ZN(n422) );
  XNOR2_X2 U545 ( .A(n600), .B(n599), .ZN(n654) );
  NAND2_X1 U546 ( .A1(n469), .A2(n467), .ZN(n573) );
  XNOR2_X2 U547 ( .A(n677), .B(KEYINPUT38), .ZN(n753) );
  XNOR2_X2 U548 ( .A(n522), .B(G122), .ZN(n551) );
  XNOR2_X2 U549 ( .A(n646), .B(KEYINPUT111), .ZN(n751) );
  AND2_X2 U550 ( .A1(n475), .A2(n470), .ZN(n468) );
  NAND2_X1 U551 ( .A1(n460), .A2(n424), .ZN(n465) );
  NAND2_X1 U552 ( .A1(n458), .A2(n459), .ZN(n424) );
  NAND2_X1 U553 ( .A1(n442), .A2(n443), .ZN(n425) );
  NAND2_X1 U554 ( .A1(n565), .A2(G221), .ZN(n434) );
  NAND2_X1 U555 ( .A1(n426), .A2(n764), .ZN(n600) );
  AND2_X1 U556 ( .A1(n595), .A2(n427), .ZN(n765) );
  INV_X1 U557 ( .A(n764), .ZN(n427) );
  XNOR2_X2 U558 ( .A(n493), .B(n492), .ZN(n565) );
  XNOR2_X1 U559 ( .A(n511), .B(n510), .ZN(n437) );
  XNOR2_X1 U560 ( .A(n633), .B(n474), .ZN(n442) );
  AND2_X1 U561 ( .A1(n644), .A2(n645), .ZN(n443) );
  NAND2_X1 U562 ( .A1(n444), .A2(n420), .ZN(n453) );
  NAND2_X1 U563 ( .A1(n616), .A2(n615), .ZN(n451) );
  XNOR2_X2 U564 ( .A(n453), .B(n452), .ZN(n748) );
  INV_X1 U565 ( .A(KEYINPUT106), .ZN(n454) );
  NAND2_X1 U566 ( .A1(n455), .A2(n464), .ZN(n459) );
  INV_X1 U567 ( .A(n690), .ZN(n455) );
  INV_X1 U568 ( .A(n456), .ZN(n461) );
  NOR2_X1 U569 ( .A1(n462), .A2(n461), .ZN(n460) );
  INV_X1 U570 ( .A(n691), .ZN(n464) );
  XNOR2_X2 U571 ( .A(KEYINPUT66), .B(G101), .ZN(n528) );
  OR2_X2 U572 ( .A1(n698), .A2(n476), .ZN(n475) );
  XNOR2_X2 U573 ( .A(G902), .B(KEYINPUT15), .ZN(n691) );
  NAND2_X1 U574 ( .A1(n466), .A2(KEYINPUT1), .ZN(n469) );
  NAND2_X1 U575 ( .A1(n478), .A2(n475), .ZN(n466) );
  NAND2_X1 U576 ( .A1(n478), .A2(n475), .ZN(n521) );
  NAND2_X1 U577 ( .A1(n468), .A2(n478), .ZN(n467) );
  INV_X1 U578 ( .A(KEYINPUT73), .ZN(n474) );
  INV_X1 U579 ( .A(n520), .ZN(n477) );
  AND2_X2 U580 ( .A1(n480), .A2(n479), .ZN(n478) );
  NAND2_X1 U581 ( .A1(n520), .A2(G902), .ZN(n479) );
  BUF_X1 U582 ( .A(n573), .Z(n627) );
  XNOR2_X2 U583 ( .A(G143), .B(G128), .ZN(n560) );
  XNOR2_X2 U584 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n481) );
  XNOR2_X2 U585 ( .A(n560), .B(n481), .ZN(n530) );
  XNOR2_X1 U586 ( .A(n482), .B(KEYINPUT70), .ZN(n483) );
  XNOR2_X1 U587 ( .A(n528), .B(G146), .ZN(n484) );
  NAND2_X1 U588 ( .A1(G210), .A2(n549), .ZN(n485) );
  XNOR2_X1 U589 ( .A(n485), .B(KEYINPUT99), .ZN(n486) );
  XNOR2_X1 U590 ( .A(n524), .B(n486), .ZN(n490) );
  XNOR2_X1 U591 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U592 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U593 ( .A(n519), .B(n491), .ZN(n720) );
  INV_X1 U594 ( .A(G472), .ZN(n719) );
  INV_X1 U595 ( .A(n652), .ZN(n509) );
  NAND2_X1 U596 ( .A1(n531), .A2(G234), .ZN(n493) );
  XNOR2_X1 U597 ( .A(n495), .B(n494), .ZN(n496) );
  NAND2_X1 U598 ( .A1(n691), .A2(G234), .ZN(n498) );
  XNOR2_X1 U599 ( .A(n499), .B(KEYINPUT14), .ZN(n500) );
  NAND2_X1 U600 ( .A1(G952), .A2(n500), .ZN(n780) );
  NOR2_X1 U601 ( .A1(G953), .A2(n780), .ZN(n582) );
  AND2_X1 U602 ( .A1(G902), .A2(n500), .ZN(n501) );
  NAND2_X1 U603 ( .A1(n501), .A2(G953), .ZN(n580) );
  NOR2_X1 U604 ( .A1(n580), .A2(G900), .ZN(n502) );
  OR2_X1 U605 ( .A1(n582), .A2(n502), .ZN(n504) );
  INV_X1 U606 ( .A(KEYINPUT81), .ZN(n503) );
  XNOR2_X1 U607 ( .A(n504), .B(n503), .ZN(n673) );
  NAND2_X1 U608 ( .A1(n505), .A2(G221), .ZN(n508) );
  INV_X1 U609 ( .A(KEYINPUT98), .ZN(n506) );
  XNOR2_X1 U610 ( .A(n506), .B(KEYINPUT21), .ZN(n507) );
  XNOR2_X1 U611 ( .A(n508), .B(n507), .ZN(n764) );
  NAND2_X1 U612 ( .A1(n509), .A2(n417), .ZN(n511) );
  INV_X1 U613 ( .A(KEYINPUT28), .ZN(n510) );
  NAND2_X1 U614 ( .A1(n531), .A2(G227), .ZN(n512) );
  XNOR2_X1 U615 ( .A(n512), .B(KEYINPUT77), .ZN(n515) );
  XNOR2_X1 U616 ( .A(n513), .B(G131), .ZN(n545) );
  INV_X1 U617 ( .A(n545), .ZN(n514) );
  XNOR2_X1 U618 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U619 ( .A(G469), .B(KEYINPUT72), .ZN(n520) );
  XNOR2_X2 U620 ( .A(G113), .B(G104), .ZN(n522) );
  XNOR2_X1 U621 ( .A(n524), .B(n562), .ZN(n525) );
  XNOR2_X1 U622 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U623 ( .A(n530), .B(n529), .ZN(n537) );
  NAND2_X1 U624 ( .A1(n531), .A2(G224), .ZN(n532) );
  XNOR2_X1 U625 ( .A(n533), .B(n532), .ZN(n535) );
  XNOR2_X1 U626 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U627 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U628 ( .A1(n731), .A2(n691), .ZN(n542) );
  NAND2_X1 U629 ( .A1(n398), .A2(n539), .ZN(n543) );
  NAND2_X1 U630 ( .A1(n543), .A2(G210), .ZN(n540) );
  XNOR2_X1 U631 ( .A(n540), .B(KEYINPUT80), .ZN(n541) );
  AND2_X1 U632 ( .A1(n543), .A2(G214), .ZN(n651) );
  INV_X1 U633 ( .A(KEYINPUT19), .ZN(n544) );
  XNOR2_X1 U634 ( .A(n546), .B(n545), .ZN(n803) );
  XNOR2_X1 U635 ( .A(n548), .B(n547), .ZN(n553) );
  NAND2_X1 U636 ( .A1(G214), .A2(n549), .ZN(n550) );
  XNOR2_X1 U637 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U638 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U639 ( .A(n803), .B(n554), .ZN(n713) );
  OR2_X1 U640 ( .A1(n713), .A2(G902), .ZN(n557) );
  XNOR2_X1 U641 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n555) );
  XNOR2_X1 U642 ( .A(n555), .B(G475), .ZN(n556) );
  XNOR2_X1 U643 ( .A(n557), .B(n556), .ZN(n676) );
  XNOR2_X1 U644 ( .A(n559), .B(n558), .ZN(n564) );
  BUF_X1 U645 ( .A(n560), .Z(n561) );
  XNOR2_X1 U646 ( .A(n561), .B(n562), .ZN(n563) );
  XNOR2_X1 U647 ( .A(n564), .B(n563), .ZN(n569) );
  AND2_X1 U648 ( .A1(n565), .A2(G217), .ZN(n567) );
  XNOR2_X1 U649 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U650 ( .A(n569), .B(n568), .ZN(n705) );
  NAND2_X1 U651 ( .A1(n705), .A2(n398), .ZN(n570) );
  XNOR2_X1 U652 ( .A(n570), .B(G478), .ZN(n674) );
  INV_X1 U653 ( .A(n661), .ZN(n609) );
  NAND2_X1 U654 ( .A1(n744), .A2(n609), .ZN(n572) );
  XNOR2_X1 U655 ( .A(G146), .B(KEYINPUT116), .ZN(n571) );
  XNOR2_X1 U656 ( .A(n572), .B(n571), .ZN(G48) );
  NOR2_X1 U657 ( .A1(n661), .A2(n651), .ZN(n614) );
  NAND2_X1 U658 ( .A1(n616), .A2(n614), .ZN(n574) );
  NOR2_X1 U659 ( .A1(n574), .A2(n627), .ZN(n577) );
  XOR2_X1 U660 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n575) );
  XOR2_X1 U661 ( .A(n575), .B(KEYINPUT108), .Z(n576) );
  XNOR2_X1 U662 ( .A(n577), .B(n576), .ZN(n579) );
  BUF_X2 U663 ( .A(n578), .Z(n677) );
  NAND2_X1 U664 ( .A1(n579), .A2(n677), .ZN(n683) );
  XNOR2_X1 U665 ( .A(n683), .B(G140), .ZN(G42) );
  NOR2_X1 U666 ( .A1(n580), .A2(G898), .ZN(n581) );
  OR2_X1 U667 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U668 ( .A(n583), .B(KEYINPUT95), .ZN(n584) );
  INV_X1 U669 ( .A(n674), .ZN(n586) );
  AND2_X1 U670 ( .A1(n586), .A2(n676), .ZN(n755) );
  NAND2_X1 U671 ( .A1(n755), .A2(n764), .ZN(n587) );
  XNOR2_X1 U672 ( .A(n587), .B(KEYINPUT105), .ZN(n588) );
  NAND2_X1 U673 ( .A1(n607), .A2(n588), .ZN(n591) );
  INV_X1 U674 ( .A(KEYINPUT74), .ZN(n589) );
  XNOR2_X1 U675 ( .A(n589), .B(KEYINPUT22), .ZN(n590) );
  XNOR2_X1 U676 ( .A(n591), .B(n590), .ZN(n594) );
  INV_X1 U677 ( .A(n627), .ZN(n762) );
  AND2_X1 U678 ( .A1(n652), .A2(n762), .ZN(n592) );
  XNOR2_X1 U679 ( .A(G110), .B(KEYINPUT114), .ZN(n593) );
  XNOR2_X1 U680 ( .A(n631), .B(n593), .ZN(G12) );
  INV_X1 U681 ( .A(n594), .ZN(n598) );
  NOR2_X1 U682 ( .A1(n420), .A2(n595), .ZN(n596) );
  NAND2_X1 U683 ( .A1(n596), .A2(n762), .ZN(n597) );
  NOR2_X1 U684 ( .A1(n598), .A2(n597), .ZN(n637) );
  XOR2_X1 U685 ( .A(G101), .B(n637), .Z(G3) );
  INV_X1 U686 ( .A(KEYINPUT68), .ZN(n599) );
  BUF_X1 U687 ( .A(n618), .Z(n601) );
  INV_X1 U688 ( .A(n601), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n603), .A2(n602), .ZN(n769) );
  NAND2_X1 U690 ( .A1(n634), .A2(n609), .ZN(n604) );
  XNOR2_X1 U691 ( .A(n604), .B(G113), .ZN(G15) );
  XNOR2_X1 U692 ( .A(G104), .B(KEYINPUT113), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n521), .A2(n652), .ZN(n605) );
  INV_X1 U694 ( .A(n654), .ZN(n761) );
  NOR2_X1 U695 ( .A1(n605), .A2(n761), .ZN(n606) );
  NAND2_X1 U696 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U697 ( .A(KEYINPUT100), .B(n608), .Z(n739) );
  NAND2_X1 U698 ( .A1(n739), .A2(n609), .ZN(n610) );
  XOR2_X1 U699 ( .A(n611), .B(n610), .Z(G6) );
  XNOR2_X1 U700 ( .A(G116), .B(KEYINPUT117), .ZN(n613) );
  NAND2_X1 U701 ( .A1(n676), .A2(n674), .ZN(n685) );
  INV_X1 U702 ( .A(n685), .ZN(n743) );
  NAND2_X1 U703 ( .A1(n634), .A2(n743), .ZN(n612) );
  XOR2_X1 U704 ( .A(n613), .B(n612), .Z(G18) );
  AND2_X1 U705 ( .A1(n614), .A2(n436), .ZN(n615) );
  XOR2_X1 U706 ( .A(G125), .B(KEYINPUT37), .Z(n617) );
  XNOR2_X1 U707 ( .A(n682), .B(n617), .ZN(G27) );
  INV_X1 U708 ( .A(n676), .ZN(n621) );
  NAND2_X1 U709 ( .A1(n621), .A2(n674), .ZN(n622) );
  NOR2_X2 U710 ( .A1(n737), .A2(KEYINPUT44), .ZN(n625) );
  INV_X1 U711 ( .A(KEYINPUT67), .ZN(n624) );
  XNOR2_X1 U712 ( .A(n625), .B(n624), .ZN(n632) );
  XNOR2_X1 U713 ( .A(n420), .B(KEYINPUT79), .ZN(n626) );
  AND2_X1 U714 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U715 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n629) );
  AND2_X1 U716 ( .A1(n709), .A2(n631), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n632), .A2(n642), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n737), .A2(KEYINPUT44), .ZN(n640) );
  INV_X1 U719 ( .A(n750), .ZN(n635) );
  NOR2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U723 ( .A(n641), .B(KEYINPUT91), .ZN(n645) );
  INV_X1 U724 ( .A(n642), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n643), .A2(KEYINPUT44), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n753), .A2(n366), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n751), .A2(n755), .ZN(n648) );
  XNOR2_X2 U728 ( .A(n648), .B(n647), .ZN(n781) );
  NOR2_X1 U729 ( .A1(n781), .A2(n649), .ZN(n650) );
  XNOR2_X1 U730 ( .A(n650), .B(KEYINPUT42), .ZN(n710) );
  INV_X1 U731 ( .A(KEYINPUT30), .ZN(n653) );
  AND2_X1 U732 ( .A1(n521), .A2(n654), .ZN(n655) );
  AND2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n680) );
  AND2_X1 U734 ( .A1(n753), .A2(n673), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n680), .A2(n657), .ZN(n660) );
  INV_X1 U736 ( .A(KEYINPUT90), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n658), .B(KEYINPUT39), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n660), .B(n659), .ZN(n686) );
  NOR2_X1 U739 ( .A1(n686), .A2(n661), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n662), .B(KEYINPUT40), .ZN(n814) );
  XOR2_X1 U741 ( .A(KEYINPUT88), .B(KEYINPUT46), .Z(n663) );
  AND2_X1 U742 ( .A1(n750), .A2(KEYINPUT82), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n744), .A2(n664), .ZN(n667) );
  INV_X1 U744 ( .A(KEYINPUT82), .ZN(n665) );
  OR2_X1 U745 ( .A1(n665), .A2(KEYINPUT47), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n665), .A2(KEYINPUT47), .ZN(n668) );
  NOR2_X1 U748 ( .A1(n750), .A2(n668), .ZN(n669) );
  AND2_X1 U749 ( .A1(n744), .A2(n669), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n674), .A2(n673), .ZN(n675) );
  OR2_X1 U751 ( .A1(n676), .A2(n675), .ZN(n678) );
  NOR2_X1 U752 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U753 ( .A1(n680), .A2(n679), .ZN(n681) );
  OR2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n688) );
  INV_X1 U755 ( .A(KEYINPUT112), .ZN(n687) );
  XNOR2_X1 U756 ( .A(n688), .B(n687), .ZN(n815) );
  NOR2_X2 U757 ( .A1(n694), .A2(n691), .ZN(n693) );
  INV_X1 U758 ( .A(KEYINPUT85), .ZN(n692) );
  BUF_X1 U759 ( .A(n694), .Z(n695) );
  INV_X1 U760 ( .A(n695), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n365), .A2(G469), .ZN(n702) );
  BUF_X1 U762 ( .A(n698), .Z(n699) );
  XOR2_X1 U763 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n700) );
  XNOR2_X1 U764 ( .A(n699), .B(n700), .ZN(n701) );
  XNOR2_X1 U765 ( .A(n702), .B(n701), .ZN(n704) );
  INV_X1 U766 ( .A(G952), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n703), .A2(G953), .ZN(n733) );
  INV_X1 U768 ( .A(n733), .ZN(n727) );
  NOR2_X1 U769 ( .A1(n704), .A2(n727), .ZN(G54) );
  NAND2_X1 U770 ( .A1(n365), .A2(G478), .ZN(n707) );
  XNOR2_X1 U771 ( .A(n705), .B(KEYINPUT125), .ZN(n706) );
  XNOR2_X1 U772 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U773 ( .A1(n708), .A2(n727), .ZN(G63) );
  XNOR2_X1 U774 ( .A(n709), .B(G119), .ZN(G21) );
  XOR2_X1 U775 ( .A(n710), .B(G137), .Z(G39) );
  XNOR2_X1 U776 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n712) );
  XNOR2_X1 U777 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U778 ( .A1(n716), .A2(n733), .ZN(n718) );
  INV_X1 U779 ( .A(KEYINPUT60), .ZN(n717) );
  XNOR2_X1 U780 ( .A(n718), .B(n717), .ZN(G60) );
  XNOR2_X1 U781 ( .A(KEYINPUT92), .B(KEYINPUT62), .ZN(n721) );
  XNOR2_X1 U782 ( .A(n364), .B(n722), .ZN(n723) );
  NAND2_X1 U783 ( .A1(n723), .A2(n733), .ZN(n724) );
  XNOR2_X1 U784 ( .A(n724), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U785 ( .A1(n365), .A2(G217), .ZN(n726) );
  XNOR2_X1 U786 ( .A(n726), .B(n725), .ZN(n728) );
  NOR2_X1 U787 ( .A1(n728), .A2(n727), .ZN(G66) );
  XNOR2_X1 U788 ( .A(KEYINPUT124), .B(KEYINPUT54), .ZN(n729) );
  XNOR2_X1 U789 ( .A(n729), .B(KEYINPUT55), .ZN(n730) );
  XNOR2_X1 U790 ( .A(n363), .B(n732), .ZN(n734) );
  NAND2_X1 U791 ( .A1(n734), .A2(n733), .ZN(n736) );
  INV_X1 U792 ( .A(KEYINPUT56), .ZN(n735) );
  XNOR2_X1 U793 ( .A(n736), .B(n735), .ZN(G51) );
  BUF_X1 U794 ( .A(n737), .Z(n738) );
  XOR2_X1 U795 ( .A(n738), .B(G122), .Z(G24) );
  XNOR2_X1 U796 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n741) );
  NAND2_X1 U797 ( .A1(n739), .A2(n743), .ZN(n740) );
  XOR2_X1 U798 ( .A(n741), .B(n740), .Z(n742) );
  XNOR2_X1 U799 ( .A(G107), .B(n742), .ZN(G9) );
  NAND2_X1 U800 ( .A1(n744), .A2(n743), .ZN(n746) );
  XOR2_X1 U801 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n745) );
  XNOR2_X1 U802 ( .A(n746), .B(n745), .ZN(n747) );
  XOR2_X1 U803 ( .A(G128), .B(n747), .Z(G30) );
  XNOR2_X1 U804 ( .A(KEYINPUT52), .B(KEYINPUT121), .ZN(n778) );
  BUF_X1 U805 ( .A(n748), .Z(n749) );
  INV_X1 U806 ( .A(n749), .ZN(n760) );
  NAND2_X1 U807 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U808 ( .A(n752), .B(KEYINPUT120), .ZN(n758) );
  NOR2_X1 U809 ( .A1(n366), .A2(n753), .ZN(n754) );
  XNOR2_X1 U810 ( .A(KEYINPUT119), .B(n754), .ZN(n756) );
  NAND2_X1 U811 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U812 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U813 ( .A1(n760), .A2(n759), .ZN(n776) );
  INV_X1 U814 ( .A(n781), .ZN(n774) );
  NAND2_X1 U815 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U816 ( .A(n763), .B(KEYINPUT50), .ZN(n768) );
  XOR2_X1 U817 ( .A(KEYINPUT49), .B(n765), .Z(n766) );
  NOR2_X1 U818 ( .A1(n602), .A2(n766), .ZN(n767) );
  NAND2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U820 ( .A1(n770), .A2(n769), .ZN(n772) );
  XOR2_X1 U821 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n771) );
  XNOR2_X1 U822 ( .A(n772), .B(n771), .ZN(n773) );
  NAND2_X1 U823 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U824 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U825 ( .A(n778), .B(n777), .ZN(n779) );
  NOR2_X1 U826 ( .A1(n780), .A2(n779), .ZN(n784) );
  NOR2_X1 U827 ( .A1(n749), .A2(n781), .ZN(n782) );
  XNOR2_X1 U828 ( .A(n782), .B(KEYINPUT122), .ZN(n783) );
  NOR2_X1 U829 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U830 ( .A(KEYINPUT123), .B(n787), .Z(n788) );
  XNOR2_X1 U831 ( .A(KEYINPUT53), .B(n789), .ZN(G75) );
  XOR2_X1 U832 ( .A(n790), .B(G101), .Z(n793) );
  INV_X1 U833 ( .A(G898), .ZN(n791) );
  NAND2_X1 U834 ( .A1(n791), .A2(G953), .ZN(n792) );
  NAND2_X1 U835 ( .A1(n793), .A2(n792), .ZN(n800) );
  NAND2_X1 U836 ( .A1(n794), .A2(n531), .ZN(n798) );
  NAND2_X1 U837 ( .A1(G953), .A2(G224), .ZN(n795) );
  XNOR2_X1 U838 ( .A(KEYINPUT61), .B(n795), .ZN(n796) );
  NAND2_X1 U839 ( .A1(n796), .A2(G898), .ZN(n797) );
  NAND2_X1 U840 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U841 ( .A(n800), .B(n799), .Z(G69) );
  BUF_X1 U842 ( .A(n801), .Z(n802) );
  XNOR2_X1 U843 ( .A(n803), .B(KEYINPUT126), .ZN(n804) );
  XOR2_X1 U844 ( .A(n802), .B(n804), .Z(n808) );
  XNOR2_X1 U845 ( .A(n805), .B(n808), .ZN(n806) );
  NOR2_X1 U846 ( .A1(n806), .A2(G953), .ZN(n807) );
  XNOR2_X1 U847 ( .A(n807), .B(KEYINPUT127), .ZN(n812) );
  XNOR2_X1 U848 ( .A(G227), .B(n808), .ZN(n809) );
  NAND2_X1 U849 ( .A1(n809), .A2(G900), .ZN(n810) );
  NAND2_X1 U850 ( .A1(n810), .A2(G953), .ZN(n811) );
  NAND2_X1 U851 ( .A1(n812), .A2(n811), .ZN(G72) );
  XNOR2_X1 U852 ( .A(G143), .B(n813), .ZN(G45) );
  XOR2_X1 U853 ( .A(G131), .B(n814), .Z(G33) );
  XOR2_X1 U854 ( .A(G134), .B(n815), .Z(G36) );
endmodule

