//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT92), .ZN(new_n209));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT89), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT90), .ZN(new_n213));
  OAI21_X1  g012(.A(G8gat), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n210), .B(KEYINPUT89), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  AOI21_X1  g015(.A(G1gat), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G8gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(KEYINPUT90), .A3(new_n218), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n214), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n214), .B2(new_n219), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n209), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n225));
  INV_X1    g024(.A(G29gat), .ZN(new_n226));
  INV_X1    g025(.A(G36gat), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n224), .A2(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G43gat), .B(G50gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(KEYINPUT15), .A3(new_n229), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n229), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT87), .B(G50gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(G43gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n225), .A2(KEYINPUT88), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n225), .A2(KEYINPUT88), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n224), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n230), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NOR3_X1   g038(.A1(new_n212), .A2(new_n213), .A3(G8gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n218), .B1(new_n215), .B2(KEYINPUT90), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n212), .A2(KEYINPUT16), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n240), .A2(new_n241), .B1(new_n242), .B2(G1gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n214), .A2(new_n217), .A3(new_n219), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(KEYINPUT92), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n222), .A2(new_n239), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT91), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n220), .B2(new_n221), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(KEYINPUT91), .A3(new_n244), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n239), .B(KEYINPUT17), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G229gat), .A2(G233gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT18), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n252), .B(KEYINPUT13), .Z(new_n256));
  INV_X1    g055(.A(new_n246), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n239), .B1(new_n222), .B2(new_n245), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n246), .A2(new_n251), .A3(KEYINPUT18), .A4(new_n252), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT93), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(KEYINPUT93), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT86), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n208), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n239), .ZN(new_n267));
  INV_X1    g066(.A(new_n245), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT92), .B1(new_n243), .B2(new_n244), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n246), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n271), .A2(new_n256), .B1(new_n253), .B2(new_n254), .ZN(new_n272));
  INV_X1    g071(.A(new_n262), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n261), .A2(KEYINPUT93), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT86), .A3(new_n207), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n266), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT97), .B(G85gat), .ZN(new_n279));
  INV_X1    g078(.A(G92gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G85gat), .A2(G92gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT7), .ZN(new_n283));
  INV_X1    g082(.A(G99gat), .ZN(new_n284));
  INV_X1    g083(.A(G106gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT8), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G99gat), .B(G106gat), .Z(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n288), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n290), .A2(new_n281), .A3(new_n283), .A4(new_n286), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n250), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n292), .ZN(new_n294));
  AND2_X1   g093(.A1(G232gat), .A2(G233gat), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n294), .A2(new_n239), .B1(KEYINPUT41), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G190gat), .B(G218gat), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n295), .A2(KEYINPUT41), .ZN(new_n303));
  XNOR2_X1  g102(.A(G134gat), .B(G162gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n297), .A2(new_n299), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n302), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n305), .B1(new_n302), .B2(new_n307), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G71gat), .A2(G78gat), .ZN(new_n312));
  OR2_X1    g111(.A1(G71gat), .A2(G78gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(G57gat), .B(G64gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT9), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT94), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n313), .A2(new_n312), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n319), .B(KEYINPUT94), .C1(new_n315), .C2(new_n314), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT95), .ZN(new_n322));
  INV_X1    g121(.A(G64gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(G57gat), .ZN(new_n324));
  INV_X1    g123(.A(G57gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(KEYINPUT95), .A3(G64gat), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n324), .B(new_n326), .C1(new_n325), .C2(G64gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(KEYINPUT96), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT96), .B1(new_n327), .B2(new_n328), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n321), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT21), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G231gat), .A2(G233gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(G127gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n268), .A2(new_n269), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n332), .A2(new_n333), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G127gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n336), .B(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n347));
  INV_X1    g146(.A(G155gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G183gat), .B(G211gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n342), .A2(new_n345), .A3(new_n351), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT98), .B1(new_n311), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(KEYINPUT98), .A3(new_n311), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n332), .A2(new_n292), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n327), .A2(KEYINPUT96), .A3(new_n328), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(new_n330), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n362), .A2(new_n321), .A3(new_n291), .A4(new_n289), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n365), .A3(new_n363), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT99), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n363), .A2(new_n365), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n360), .A2(KEYINPUT99), .A3(new_n363), .A4(new_n365), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G230gat), .A2(G233gat), .ZN(new_n372));
  MUX2_X1   g171(.A(new_n364), .B(new_n371), .S(new_n372), .Z(new_n373));
  XNOR2_X1  g172(.A(G120gat), .B(G148gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G176gat), .B(G204gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  XOR2_X1   g175(.A(new_n376), .B(KEYINPUT101), .Z(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n366), .A2(new_n367), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n370), .A2(new_n369), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT100), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT100), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n368), .A2(new_n382), .A3(new_n369), .A4(new_n370), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n383), .A3(new_n372), .ZN(new_n384));
  INV_X1    g183(.A(new_n376), .ZN(new_n385));
  INV_X1    g184(.A(new_n372), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n364), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n378), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n359), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(G197gat), .A2(G204gat), .ZN(new_n399));
  AND2_X1   g198(.A1(G197gat), .A2(G204gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G211gat), .B(G218gat), .Z(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G211gat), .B(G218gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G197gat), .B(G204gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n398), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G226gat), .ZN(new_n409));
  INV_X1    g208(.A(G233gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT67), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT27), .B(G183gat), .ZN(new_n413));
  INV_X1    g212(.A(G190gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n415), .A2(KEYINPUT28), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(KEYINPUT28), .ZN(new_n417));
  NOR2_X1   g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT26), .ZN(new_n419));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G169gat), .ZN(new_n422));
  INV_X1    g221(.A(G176gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n416), .A2(new_n417), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n418), .A2(KEYINPUT23), .ZN(new_n428));
  NAND2_X1  g227(.A1(G169gat), .A2(G176gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT23), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(G169gat), .B2(G176gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT64), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT24), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n420), .ZN(new_n435));
  NOR2_X1   g234(.A1(G183gat), .A2(G190gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT64), .B(KEYINPUT24), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n435), .B(new_n437), .C1(new_n438), .C2(new_n420), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n432), .B1(new_n439), .B2(KEYINPUT65), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n436), .B1(new_n434), .B2(new_n420), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n441), .B(new_n442), .C1(new_n420), .C2(new_n438), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT25), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n432), .ZN(new_n445));
  OR2_X1    g244(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(new_n420), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT25), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n437), .A2(new_n446), .A3(new_n420), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n427), .B1(new_n444), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT29), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n411), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n411), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n437), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT24), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT64), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n420), .B1(new_n434), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT65), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n443), .A3(new_n445), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n448), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n451), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n456), .B1(new_n464), .B2(new_n427), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n408), .B1(new_n455), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n453), .A2(new_n411), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT29), .B1(new_n464), .B2(new_n427), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n467), .B(new_n407), .C1(new_n468), .C2(new_n411), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n466), .A2(KEYINPUT72), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT72), .B1(new_n466), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n395), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n394), .A3(new_n469), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT73), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT30), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT30), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(KEYINPUT73), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT76), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480));
  NAND2_X1  g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT2), .ZN(new_n482));
  OR2_X1    g281(.A1(G141gat), .A2(G148gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(G141gat), .A2(G148gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(KEYINPUT74), .A3(new_n484), .ZN(new_n486));
  INV_X1    g285(.A(new_n481), .ZN(new_n487));
  NOR2_X1   g286(.A1(G155gat), .A2(G162gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(G141gat), .A2(G148gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(G141gat), .A2(G148gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G155gat), .B(G162gat), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n493), .B(new_n482), .C1(new_n494), .C2(KEYINPUT74), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G113gat), .ZN(new_n497));
  INV_X1    g296(.A(G120gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT1), .ZN(new_n500));
  NAND2_X1  g299(.A1(G113gat), .A2(G120gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(G127gat), .A2(G134gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(G127gat), .A2(G134gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(G113gat), .A2(G120gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(G113gat), .A2(G120gat), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT69), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT69), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n499), .A2(new_n510), .A3(new_n501), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n511), .A3(new_n500), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT68), .B(G127gat), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n504), .B1(new_n513), .B2(G134gat), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n506), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n490), .A2(new_n495), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT3), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n512), .A2(new_n514), .ZN(new_n521));
  INV_X1    g320(.A(new_n506), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT3), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n490), .A2(new_n495), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G225gat), .A2(G233gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n496), .A2(new_n515), .A3(KEYINPUT4), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n518), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT5), .ZN(new_n530));
  AND2_X1   g329(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n532));
  OAI21_X1  g331(.A(G134gat), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n504), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n499), .A2(new_n501), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT1), .B1(new_n536), .B2(KEYINPUT69), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n535), .B1(new_n537), .B2(new_n511), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n519), .B1(new_n538), .B2(new_n506), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n516), .ZN(new_n540));
  INV_X1    g339(.A(new_n527), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n530), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n526), .A2(new_n530), .A3(new_n527), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT4), .B1(new_n496), .B2(new_n515), .ZN(new_n544));
  INV_X1    g343(.A(new_n516), .ZN(new_n545));
  INV_X1    g344(.A(new_n517), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n529), .A2(new_n542), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G1gat), .B(G29gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT0), .ZN(new_n550));
  XNOR2_X1  g349(.A(G57gat), .B(G85gat), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n550), .B(new_n551), .Z(new_n552));
  OAI21_X1  g351(.A(new_n480), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n542), .A2(new_n529), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n543), .A2(new_n547), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n554), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n479), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n555), .ZN(new_n558));
  INV_X1    g357(.A(new_n552), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT6), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n548), .A2(new_n552), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT76), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(KEYINPUT6), .A3(new_n559), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n557), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n478), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n453), .A2(new_n515), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n464), .A2(new_n523), .A3(new_n427), .ZN(new_n567));
  INV_X1    g366(.A(G227gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(new_n410), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT32), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n574));
  XNOR2_X1  g373(.A(G15gat), .B(G43gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G99gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n577), .B1(new_n570), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n570), .B(KEYINPUT32), .C1(new_n578), .C2(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n583));
  INV_X1    g382(.A(new_n569), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT34), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n583), .A2(new_n587), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n580), .A2(new_n581), .B1(new_n586), .B2(new_n588), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT81), .ZN(new_n593));
  AND2_X1   g392(.A1(G228gat), .A2(G233gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n401), .A2(new_n402), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n404), .B1(new_n398), .B2(new_n405), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n454), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n597), .A2(new_n524), .B1(new_n495), .B2(new_n490), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n407), .B1(new_n525), .B2(new_n454), .ZN(new_n599));
  OAI211_X1 g398(.A(KEYINPUT77), .B(new_n594), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n525), .A2(new_n454), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n408), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT29), .B1(new_n403), .B2(new_n406), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n519), .B1(new_n603), .B2(KEYINPUT3), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n594), .A2(KEYINPUT77), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n594), .A2(KEYINPUT77), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n602), .A2(new_n604), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n600), .A2(new_n607), .A3(KEYINPUT78), .A4(G22gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G78gat), .B(G106gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT31), .B(G50gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n600), .A2(new_n607), .ZN(new_n614));
  INV_X1    g413(.A(G22gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT79), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n600), .A2(G22gat), .A3(new_n607), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT78), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT79), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n614), .A2(new_n621), .A3(new_n615), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n613), .A2(new_n617), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT80), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n614), .B2(new_n615), .ZN(new_n625));
  AOI211_X1 g424(.A(KEYINPUT79), .B(G22gat), .C1(new_n600), .C2(new_n607), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT80), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n627), .A2(new_n628), .A3(new_n613), .A4(new_n620), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n612), .B1(new_n616), .B2(new_n618), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n593), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AOI211_X1 g432(.A(KEYINPUT81), .B(new_n631), .C1(new_n624), .C2(new_n629), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n565), .B(new_n592), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT35), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT83), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n635), .A2(KEYINPUT83), .A3(KEYINPUT35), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT35), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n560), .A2(KEYINPUT82), .A3(new_n561), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n563), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT82), .B1(new_n560), .B2(new_n561), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n478), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n645), .B(new_n592), .C1(new_n633), .C2(new_n634), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n638), .A2(new_n639), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT84), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n633), .A2(new_n634), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n470), .A2(new_n471), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n466), .A2(new_n651), .A3(new_n469), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(KEYINPUT38), .A3(new_n395), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n395), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n651), .B1(new_n466), .B2(new_n469), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI22_X1  g456(.A1(new_n652), .A2(new_n654), .B1(new_n657), .B2(KEYINPUT38), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n473), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n547), .A2(new_n526), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n541), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n662), .B(KEYINPUT39), .C1(new_n541), .C2(new_n540), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n663), .B(new_n552), .C1(KEYINPUT39), .C2(new_n662), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n558), .A2(new_n559), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n478), .A2(new_n666), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n649), .A2(new_n660), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n582), .B(new_n589), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT36), .B1(new_n671), .B2(KEYINPUT71), .ZN(new_n672));
  OAI211_X1 g471(.A(KEYINPUT71), .B(KEYINPUT36), .C1(new_n590), .C2(new_n591), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n633), .A2(new_n634), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n564), .B2(new_n478), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n670), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n647), .A2(new_n648), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n648), .B1(new_n647), .B2(new_n678), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n278), .B(new_n391), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n635), .A2(KEYINPUT83), .A3(KEYINPUT35), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT83), .B1(new_n635), .B2(KEYINPUT35), .ZN(new_n685));
  INV_X1    g484(.A(new_n646), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n670), .A2(new_n675), .A3(new_n677), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT84), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n647), .A2(new_n648), .A3(new_n678), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n691), .A2(KEYINPUT102), .A3(new_n278), .A4(new_n391), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n564), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n478), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT16), .B(G8gat), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n698), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n696), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT103), .B1(new_n698), .B2(KEYINPUT42), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n701), .B(new_n702), .C1(new_n696), .C2(new_n697), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n699), .A2(new_n700), .A3(new_n703), .ZN(G1325gat));
  INV_X1    g503(.A(G15gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n693), .A2(new_n705), .A3(new_n592), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n675), .B1(new_n683), .B2(new_n692), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n705), .ZN(G1326gat));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n693), .B2(new_n676), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AOI211_X1 g511(.A(KEYINPUT104), .B(new_n649), .C1(new_n683), .C2(new_n692), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n709), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n709), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n711), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(new_n717), .ZN(G1327gat));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n691), .B2(new_n310), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n647), .A2(new_n678), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n647), .B2(new_n678), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n310), .A2(new_n719), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n355), .B(KEYINPUT105), .Z(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(new_n277), .A3(new_n390), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n564), .ZN(new_n732));
  OAI21_X1  g531(.A(G29gat), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n311), .A2(new_n355), .A3(new_n390), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n691), .A2(new_n278), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n564), .A2(new_n226), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n736), .A2(new_n734), .A3(new_n737), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n733), .A2(new_n738), .A3(new_n739), .ZN(G1328gat));
  INV_X1    g539(.A(new_n478), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n731), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n478), .A2(new_n227), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT46), .B1(new_n736), .B2(new_n743), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n743), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(G1329gat));
  OR2_X1    g545(.A1(new_n671), .A2(G43gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n736), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n675), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n749), .B(new_n730), .C1(new_n720), .C2(new_n726), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n748), .B1(new_n750), .B2(G43gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g551(.A1(new_n649), .A2(new_n233), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n736), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n676), .B(new_n730), .C1(new_n720), .C2(new_n726), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(new_n233), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g556(.A1(new_n722), .A2(new_n724), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n359), .A2(new_n278), .A3(new_n389), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n732), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n325), .ZN(G1332gat));
  NOR2_X1   g561(.A1(new_n760), .A2(new_n741), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(G1333gat));
  OAI21_X1  g566(.A(G71gat), .B1(new_n760), .B2(new_n675), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n671), .A2(G71gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n760), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g570(.A1(new_n760), .A2(new_n649), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g572(.A1(new_n278), .A2(new_n355), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n310), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n647), .B2(new_n678), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n776), .A2(KEYINPUT51), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT107), .B1(new_n777), .B2(new_n778), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n781), .A2(new_n389), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n783), .A2(new_n564), .A3(new_n279), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n774), .A2(new_n390), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n727), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n732), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n784), .B1(new_n788), .B2(new_n279), .ZN(G1336gat));
  OAI211_X1 g588(.A(new_n478), .B(new_n786), .C1(new_n720), .C2(new_n726), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G92gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n779), .A2(new_n390), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n478), .A2(new_n280), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT52), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n791), .B(new_n796), .C1(new_n792), .C2(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n787), .B2(new_n675), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n284), .A3(new_n592), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(G1338gat));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n676), .B(new_n786), .C1(new_n720), .C2(new_n726), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(G106gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n676), .A2(new_n285), .ZN(new_n805));
  AOI211_X1 g604(.A(new_n389), .B(new_n805), .C1(new_n777), .C2(new_n778), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n803), .B2(G106gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n804), .A2(new_n807), .A3(KEYINPUT53), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  AOI221_X4 g608(.A(new_n806), .B1(new_n802), .B2(new_n809), .C1(new_n803), .C2(G106gat), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n808), .A2(new_n810), .ZN(G1339gat));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n371), .A2(new_n812), .A3(new_n372), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n385), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(new_n386), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT54), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n814), .B1(new_n384), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n818), .A2(KEYINPUT55), .B1(new_n384), .B2(new_n387), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n384), .A2(new_n817), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n813), .A2(new_n385), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n266), .A2(new_n276), .A3(new_n819), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n264), .A2(new_n207), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n271), .A2(new_n256), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n252), .B1(new_n246), .B2(new_n251), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n206), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n390), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n310), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n826), .A2(new_n310), .A3(new_n829), .A4(new_n824), .ZN(new_n832));
  INV_X1    g631(.A(new_n819), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n728), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n357), .A2(new_n277), .A3(new_n358), .A4(new_n389), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n676), .B(new_n671), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n732), .A2(new_n478), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n278), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n390), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n729), .ZN(new_n844));
  INV_X1    g643(.A(new_n355), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n513), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n844), .A2(new_n513), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT109), .Z(G1342gat));
  AOI21_X1  g647(.A(new_n311), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n839), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT110), .ZN(new_n851));
  NOR2_X1   g650(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(new_n852), .ZN(G1343gat));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n836), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n676), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n675), .A2(new_n838), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n277), .A2(G141gat), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n854), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n864));
  INV_X1    g663(.A(new_n857), .ZN(new_n865));
  XNOR2_X1  g664(.A(KEYINPUT111), .B(KEYINPUT57), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n855), .B2(new_n676), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n386), .B1(new_n371), .B2(KEYINPUT100), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n816), .B1(new_n870), .B2(new_n383), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT112), .B1(new_n871), .B2(new_n814), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n820), .A2(new_n873), .A3(new_n821), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n874), .A3(new_n823), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n266), .A2(new_n875), .A3(new_n819), .A4(new_n276), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n310), .B1(new_n876), .B2(new_n830), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n845), .B1(new_n877), .B2(new_n834), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n869), .B(new_n649), .C1(new_n878), .C2(new_n836), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n865), .B1(new_n868), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n277), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n863), .A2(new_n864), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n864), .B1(new_n863), .B2(new_n881), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n881), .A2(new_n860), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n882), .A2(new_n883), .B1(new_n854), .B2(new_n884), .ZN(G1344gat));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n886));
  INV_X1    g685(.A(G148gat), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n649), .B1(new_n878), .B2(new_n836), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n856), .A2(new_n866), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n390), .B1(new_n857), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n890), .B2(new_n857), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n887), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n888), .A2(KEYINPUT57), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n649), .B(new_n866), .C1(new_n835), .C2(new_n836), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G148gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n390), .B(new_n865), .C1(new_n868), .C2(new_n879), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n887), .A2(KEYINPUT59), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(KEYINPUT115), .A3(new_n902), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n895), .A2(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n858), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(G148gat), .A3(new_n389), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT118), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT117), .B1(new_n899), .B2(KEYINPUT59), .ZN(new_n911));
  AOI211_X1 g710(.A(new_n886), .B(new_n894), .C1(new_n898), .C2(G148gat), .ZN(new_n912));
  INV_X1    g711(.A(new_n906), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT115), .B1(new_n901), .B2(new_n902), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n911), .A2(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  INV_X1    g715(.A(new_n909), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n910), .A2(new_n918), .ZN(G1345gat));
  NOR2_X1   g718(.A1(new_n908), .A2(new_n845), .ZN(new_n920));
  AOI21_X1  g719(.A(G155gat), .B1(new_n920), .B2(KEYINPUT119), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(KEYINPUT119), .B2(new_n920), .ZN(new_n922));
  OR3_X1    g721(.A1(new_n880), .A2(new_n348), .A3(new_n728), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n880), .B2(new_n311), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n311), .A2(G162gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n908), .B2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n741), .A2(new_n564), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n837), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n277), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(new_n422), .ZN(G1348gat));
  OAI22_X1  g730(.A1(new_n929), .A2(new_n389), .B1(KEYINPUT120), .B2(new_n423), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n423), .A2(KEYINPUT120), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n932), .B(new_n933), .Z(G1349gat));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n929), .A2(new_n935), .A3(new_n728), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n929), .B2(new_n728), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G183gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n355), .A2(new_n413), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n936), .A2(new_n938), .B1(new_n929), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT60), .ZN(G1350gat));
  OAI22_X1  g740(.A1(new_n929), .A2(new_n311), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n942), .B(new_n943), .ZN(G1351gat));
  NAND3_X1  g743(.A1(new_n675), .A2(new_n676), .A3(new_n928), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n835), .B2(new_n836), .ZN(new_n946));
  AOI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n278), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n889), .B(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n675), .A2(new_n928), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(G197gat), .A3(new_n278), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(new_n948), .B2(new_n951), .ZN(G1352gat));
  INV_X1    g751(.A(G204gat), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n949), .A2(new_n389), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n948), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n389), .A2(G204gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n946), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n946), .A2(new_n956), .A3(new_n957), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n959), .A2(KEYINPUT62), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT62), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n955), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n955), .B2(new_n963), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1353gat));
  INV_X1    g766(.A(G211gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n946), .A2(new_n968), .A3(new_n355), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n889), .A2(new_n355), .A3(new_n950), .ZN(new_n971));
  AND4_X1   g770(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT63), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(KEYINPUT125), .B2(new_n973), .ZN(new_n974));
  AOI22_X1  g773(.A1(new_n971), .A2(new_n974), .B1(new_n970), .B2(KEYINPUT63), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n969), .B1(new_n972), .B2(new_n975), .ZN(G1354gat));
  AOI21_X1  g775(.A(G218gat), .B1(new_n946), .B2(new_n310), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n310), .A2(G218gat), .ZN(new_n978));
  XOR2_X1   g777(.A(new_n978), .B(KEYINPUT126), .Z(new_n979));
  NOR2_X1   g778(.A1(new_n949), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n977), .B1(new_n948), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g780(.A(new_n981), .B(KEYINPUT127), .Z(G1355gat));
endmodule


