//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G197gat), .ZN(new_n203));
  INV_X1    g002(.A(G204gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  NAND2_X1  g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G211gat), .ZN(new_n211));
  INV_X1    g010(.A(G218gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(new_n208), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n214), .B1(new_n213), .B2(new_n208), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n210), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n217), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(new_n209), .A3(new_n215), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT80), .B1(new_n223), .B2(G141gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(G141gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n224), .A2(new_n227), .A3(KEYINPUT81), .A4(new_n228), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  INV_X1    g033(.A(G162gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT2), .ZN(new_n237));
  NOR2_X1   g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n226), .A2(G148gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT2), .B1(new_n243), .B2(new_n228), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n244), .A2(new_n236), .A3(new_n238), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n222), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n239), .B1(new_n231), .B2(new_n232), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(new_n245), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n218), .A2(new_n248), .A3(new_n220), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n251), .B1(new_n242), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G228gat), .ZN(new_n254));
  INV_X1    g053(.A(G233gat), .ZN(new_n255));
  OAI22_X1  g054(.A1(new_n249), .A2(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n250), .A2(KEYINPUT3), .A3(new_n245), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n221), .B1(new_n257), .B2(KEYINPUT29), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n242), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n250), .B2(new_n245), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n254), .A2(new_n255), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n202), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n264));
  INV_X1    g063(.A(G50gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G78gat), .B(G106gat), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n202), .A3(new_n262), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT89), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n256), .A2(new_n262), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G22gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n276), .A3(G22gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n275), .B1(new_n282), .B2(new_n271), .ZN(new_n283));
  AOI211_X1 g082(.A(KEYINPUT89), .B(new_n270), .C1(new_n280), .C2(new_n281), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n274), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G1gat), .B(G29gat), .Z(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G57gat), .B(G85gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(KEYINPUT1), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294));
  INV_X1    g093(.A(G113gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(G120gat), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G113gat), .ZN(new_n298));
  OAI211_X1 g097(.A(KEYINPUT72), .B(new_n294), .C1(new_n296), .C2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n293), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n292), .A2(KEYINPUT1), .ZN(new_n302));
  INV_X1    g101(.A(new_n300), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(KEYINPUT72), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT3), .B1(new_n250), .B2(new_n245), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n247), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n241), .A2(new_n305), .A3(new_n246), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n305), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT39), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n304), .B(new_n301), .C1(new_n250), .C2(new_n245), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n317), .B1(new_n319), .B2(new_n314), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n290), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n313), .A2(new_n317), .A3(new_n315), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(KEYINPUT40), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G169gat), .ZN(new_n326));
  INV_X1    g125(.A(G176gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT23), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT65), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT24), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(G183gat), .A3(G190gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G183gat), .ZN(new_n339));
  INV_X1    g138(.A(G190gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT66), .B1(new_n331), .B2(KEYINPUT23), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n345), .B(new_n346), .C1(G169gat), .C2(G176gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n333), .A2(new_n342), .A3(new_n343), .A4(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT68), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR3_X1   g152(.A1(KEYINPUT68), .A2(G183gat), .A3(G190gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT67), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n346), .B1(new_n331), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n355), .A2(new_n338), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n343), .A2(KEYINPUT25), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n360), .B1(new_n344), .B2(new_n347), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n351), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n339), .A2(KEYINPUT27), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT27), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G183gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n364), .B1(new_n368), .B2(G190gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT27), .B(G183gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(KEYINPUT69), .A3(new_n340), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(KEYINPUT70), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT28), .A4(new_n340), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n356), .A2(KEYINPUT71), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT26), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(KEYINPUT71), .A2(KEYINPUT26), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT67), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n331), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n385), .A2(new_n343), .B1(G183gat), .B2(G190gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n363), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n389), .B(KEYINPUT79), .Z(new_n390));
  NOR2_X1   g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n363), .B2(new_n387), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n221), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  AOI22_X1  g195(.A1(new_n379), .A2(new_n380), .B1(new_n331), .B2(new_n383), .ZN(new_n397));
  INV_X1    g196(.A(new_n343), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n334), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(new_n373), .B2(new_n377), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n349), .A2(new_n350), .B1(new_n359), .B2(new_n361), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n248), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n389), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n390), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n222), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n393), .A2(new_n396), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n407), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n405), .ZN(new_n410));
  INV_X1    g209(.A(new_n396), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT82), .B1(new_n319), .B2(new_n314), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT5), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n314), .B1(new_n309), .B2(new_n318), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n308), .A2(new_n311), .A3(new_n314), .A4(new_n312), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n311), .A2(new_n312), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n422), .A2(new_n415), .A3(new_n314), .A4(new_n308), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n421), .B1(new_n419), .B2(KEYINPUT5), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(new_n419), .A3(new_n414), .A4(new_n418), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n426), .A3(new_n290), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n321), .A2(new_n322), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n428), .A2(KEYINPUT40), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n325), .A2(new_n413), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  INV_X1    g230(.A(new_n390), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n392), .B1(new_n432), .B2(new_n402), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n405), .B(new_n431), .C1(new_n433), .C2(new_n222), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n393), .A2(KEYINPUT91), .A3(new_n431), .A4(new_n405), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n403), .A2(new_n221), .A3(new_n404), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n439), .A2(KEYINPUT37), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n222), .B1(new_n391), .B2(new_n392), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT38), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n442), .A3(new_n411), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n431), .B1(new_n393), .B2(new_n405), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n396), .B(new_n444), .C1(new_n436), .C2(new_n437), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT38), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n406), .B(new_n443), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n290), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n420), .B1(new_n421), .B2(new_n423), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n416), .A2(new_n417), .ZN(new_n450));
  AOI211_X1 g249(.A(KEYINPUT82), .B(new_n314), .C1(new_n309), .C2(new_n318), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n450), .A2(new_n451), .A3(new_n415), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n425), .B1(new_n452), .B2(new_n419), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n448), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n427), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT6), .A4(new_n290), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n285), .B(new_n430), .C1(new_n447), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n413), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n424), .A2(new_n426), .A3(new_n290), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n290), .B1(new_n424), .B2(new_n426), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT6), .ZN(new_n463));
  INV_X1    g262(.A(new_n457), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n263), .B1(new_n276), .B2(new_n273), .ZN(new_n466));
  INV_X1    g265(.A(new_n281), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n271), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT89), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n282), .A2(new_n275), .A3(new_n271), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n469), .A2(new_n470), .B1(new_n273), .B2(new_n272), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT32), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n305), .B1(new_n400), .B2(new_n401), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n363), .A2(new_n387), .A3(new_n306), .ZN(new_n475));
  NAND2_X1  g274(.A1(G227gat), .A2(G233gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n476), .B(KEYINPUT64), .Z(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT73), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n474), .A2(new_n475), .A3(new_n480), .A4(new_n477), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n473), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT33), .B1(new_n479), .B2(new_n481), .ZN(new_n483));
  XOR2_X1   g282(.A(KEYINPUT74), .B(G71gat), .Z(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(G99gat), .ZN(new_n485));
  XOR2_X1   g284(.A(G15gat), .B(G43gat), .Z(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n482), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  AOI221_X4 g288(.A(new_n473), .B1(KEYINPUT33), .B2(new_n487), .C1(new_n479), .C2(new_n481), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT75), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT75), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n476), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT34), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n477), .A2(KEYINPUT34), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n474), .B2(new_n475), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT76), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n489), .A2(new_n490), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n491), .A2(new_n492), .B1(G227gat), .B2(G233gat), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(new_n494), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n491), .A2(new_n497), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT76), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT76), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n499), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n479), .A2(new_n481), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT32), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n515), .A3(new_n487), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n482), .B1(new_n483), .B2(new_n488), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT77), .B1(new_n502), .B2(new_n518), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n501), .B1(new_n489), .B2(new_n490), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT77), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n459), .A2(new_n472), .A3(new_n521), .A4(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n413), .B1(new_n456), .B2(new_n457), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n285), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n522), .A2(new_n526), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n456), .B2(new_n457), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(new_n285), .A3(new_n460), .A4(new_n519), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n528), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G57gat), .B(G64gat), .Z(new_n537));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n540), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  XNOR2_X1  g340(.A(G71gat), .B(G78gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT21), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G127gat), .ZN(new_n548));
  XOR2_X1   g347(.A(G15gat), .B(G22gat), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(G1gat), .ZN(new_n550));
  INV_X1    g349(.A(G1gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT16), .ZN(new_n552));
  OAI221_X1 g351(.A(new_n550), .B1(KEYINPUT95), .B2(G8gat), .C1(new_n549), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(KEYINPUT95), .A2(G8gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n543), .B2(new_n544), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n548), .A2(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT98), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G155gat), .ZN(new_n562));
  XOR2_X1   g361(.A(G183gat), .B(G211gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n557), .A2(new_n558), .A3(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G29gat), .ZN(new_n570));
  INV_X1    g369(.A(G36gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT14), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT14), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(G29gat), .B2(G36gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT94), .Z(new_n576));
  INV_X1    g375(.A(G43gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G50gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n265), .A2(G43gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT93), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT15), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n580), .B(new_n581), .C1(KEYINPUT93), .C2(new_n578), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT15), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G29gat), .A2(G36gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT92), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n576), .A2(new_n582), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n584), .B1(new_n586), .B2(new_n575), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT17), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n589), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT8), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n596), .B(new_n598), .C1(G85gat), .C2(G92gat), .ZN(new_n599));
  XOR2_X1   g398(.A(G99gat), .B(G106gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT99), .B1(new_n599), .B2(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n591), .A2(new_n594), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT41), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n606), .B(new_n608), .C1(new_n590), .C2(new_n605), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G134gat), .B(G162gat), .Z(new_n612));
  NOR2_X1   g411(.A1(new_n607), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n614), .A2(KEYINPUT100), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(KEYINPUT100), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n611), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n543), .A2(new_n601), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n620), .B1(new_n543), .B2(new_n605), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OR3_X1    g422(.A1(new_n605), .A2(new_n543), .A3(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT101), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  OAI211_X1 g431(.A(new_n629), .B(new_n632), .C1(new_n628), .C2(new_n621), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n627), .B1(new_n623), .B2(new_n624), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n621), .A2(new_n628), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n633), .A2(KEYINPUT102), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT102), .B1(new_n633), .B2(new_n637), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n569), .A2(new_n619), .A3(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(KEYINPUT103), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n555), .A2(new_n590), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n555), .A2(new_n594), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n591), .ZN(new_n645));
  NAND2_X1  g444(.A1(G229gat), .A2(G233gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(KEYINPUT18), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n555), .B(new_n590), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n646), .B(KEYINPUT13), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G113gat), .B(G141gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G197gat), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT11), .B(G169gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT12), .Z(new_n656));
  NOR2_X1   g455(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n645), .A2(new_n646), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT96), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(new_n662), .A3(new_n659), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n657), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n660), .A2(new_n650), .A3(new_n647), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n656), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n641), .A2(KEYINPUT103), .ZN(new_n668));
  AND4_X1   g467(.A1(new_n536), .A2(new_n642), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n458), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n413), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n673), .A2(KEYINPUT104), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(KEYINPUT104), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(G8gat), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT16), .B(G8gat), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n673), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n674), .B2(new_n675), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n676), .B(new_n679), .C1(new_n680), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g480(.A(G15gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n532), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n669), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n521), .A2(new_n527), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n669), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n684), .B1(new_n687), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n471), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NAND3_X1  g490(.A1(new_n568), .A2(new_n640), .A3(new_n667), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n619), .A2(KEYINPUT44), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n528), .B(KEYINPUT105), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n533), .A2(new_n535), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n533), .A2(KEYINPUT106), .A3(new_n535), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n695), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  INV_X1    g502(.A(new_n619), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n536), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n693), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n458), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n536), .A2(new_n704), .A3(new_n693), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n570), .A3(new_n670), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n708), .A2(new_n571), .A3(new_n413), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT46), .Z(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n706), .B2(new_n460), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n528), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n685), .A2(KEYINPUT105), .A3(new_n459), .A4(new_n472), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n533), .A2(KEYINPUT106), .A3(new_n535), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT106), .B1(new_n533), .B2(new_n535), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n705), .B1(new_n721), .B2(new_n694), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n722), .A2(new_n685), .A3(new_n692), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(KEYINPUT109), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(KEYINPUT109), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(G43gat), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n532), .A2(G43gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(KEYINPUT47), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n728), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n686), .B(new_n693), .C1(new_n702), .C2(new_n705), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G43gat), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n730), .B1(new_n732), .B2(KEYINPUT107), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n734), .A3(G43gat), .ZN(new_n735));
  AOI211_X1 g534(.A(KEYINPUT108), .B(KEYINPUT47), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT107), .B1(new_n723), .B2(new_n577), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n735), .A3(new_n728), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n729), .B1(new_n736), .B2(new_n741), .ZN(G1330gat));
  NAND3_X1  g541(.A1(new_n708), .A2(new_n265), .A3(new_n471), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n706), .A2(new_n285), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n265), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g545(.A(new_n640), .ZN(new_n747));
  INV_X1    g546(.A(new_n667), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n569), .A2(new_n747), .A3(new_n748), .A4(new_n619), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n696), .B2(new_n701), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n458), .B(KEYINPUT110), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n413), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT49), .B(G64gat), .Z(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(G1333gat));
  NAND2_X1  g557(.A1(new_n750), .A2(new_n683), .ZN(new_n759));
  INV_X1    g558(.A(G71gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n685), .A2(new_n760), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n750), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n750), .B2(new_n763), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n471), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g568(.A1(new_n640), .A2(G85gat), .A3(new_n458), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n568), .A2(new_n748), .ZN(new_n771));
  AOI211_X1 g570(.A(new_n619), .B(new_n771), .C1(new_n696), .C2(new_n701), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n773), .A2(KEYINPUT112), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT112), .B1(new_n773), .B2(new_n774), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n770), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n722), .A2(new_n640), .A3(new_n771), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779), .B2(new_n458), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(G1336gat));
  NOR2_X1   g580(.A1(new_n640), .A2(new_n460), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n460), .A2(new_n786), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n778), .B2(new_n790), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n787), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n788), .B1(new_n787), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(G1337gat));
  NOR3_X1   g593(.A1(new_n640), .A2(G99gat), .A3(new_n532), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT114), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n775), .B2(new_n776), .ZN(new_n797));
  OAI21_X1  g596(.A(G99gat), .B1(new_n779), .B2(new_n685), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1338gat));
  INV_X1    g598(.A(G106gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n778), .A2(new_n471), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n773), .A2(new_n774), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n640), .A2(G106gat), .A3(new_n285), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n800), .B1(new_n778), .B2(new_n471), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n632), .B1(new_n635), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n629), .A2(KEYINPUT54), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n625), .A2(new_n628), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT55), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n633), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n816), .A2(new_n813), .A3(new_n635), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n634), .B1(new_n629), .B2(KEYINPUT54), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n704), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n645), .A2(new_n646), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n648), .A2(new_n649), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n655), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n664), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n664), .B(new_n826), .C1(new_n638), .C2(new_n639), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n667), .A2(new_n822), .A3(new_n633), .A4(new_n817), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n704), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT116), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n828), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n835), .A2(new_n569), .B1(new_n667), .B2(new_n641), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n752), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n520), .A2(new_n471), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n460), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n667), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n641), .A2(new_n667), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n833), .A2(new_n834), .ZN(new_n846));
  INV_X1    g645(.A(new_n828), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n848), .B2(new_n568), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n683), .A2(new_n285), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n458), .A2(new_n413), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n748), .A2(new_n295), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n844), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  AOI21_X1  g657(.A(G120gat), .B1(new_n843), .B2(new_n747), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n640), .A2(new_n297), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n856), .B2(new_n860), .ZN(G1341gat));
  AND2_X1   g660(.A1(new_n569), .A2(G127gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n838), .A2(new_n841), .A3(new_n569), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(G127gat), .B1(new_n863), .B2(new_n864), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n856), .A2(new_n862), .B1(new_n865), .B2(new_n866), .ZN(G1342gat));
  OR4_X1    g666(.A1(G134gat), .A2(new_n837), .A3(new_n840), .A4(new_n619), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n855), .B2(new_n619), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1343gat));
  NOR3_X1   g671(.A1(new_n686), .A2(new_n285), .A3(new_n413), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n837), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT119), .B1(new_n836), .B2(new_n752), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n748), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n685), .A2(new_n852), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n831), .A2(new_n619), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n569), .B1(new_n847), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n471), .B1(new_n880), .B2(new_n845), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n878), .B1(new_n881), .B2(KEYINPUT57), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n836), .A2(new_n471), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n667), .A2(G141gat), .ZN(new_n885));
  OAI22_X1  g684(.A1(new_n877), .A2(G141gat), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI221_X1 g687(.A(KEYINPUT58), .B1(new_n884), .B2(new_n885), .C1(new_n877), .C2(G141gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n876), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n223), .A3(new_n747), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT57), .B1(new_n849), .B2(new_n285), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n823), .A2(KEYINPUT120), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n818), .A2(new_n704), .A3(new_n896), .A4(new_n822), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n895), .A2(new_n664), .A3(new_n826), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n879), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n568), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n642), .A2(new_n668), .A3(new_n748), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n285), .A2(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n878), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n894), .A2(new_n904), .A3(new_n747), .A4(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n223), .B1(new_n906), .B2(KEYINPUT121), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n883), .A2(KEYINPUT57), .B1(new_n902), .B2(new_n903), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n747), .A4(new_n905), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n893), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n884), .A2(new_n640), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(KEYINPUT59), .A3(new_n223), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n892), .B1(new_n911), .B2(new_n913), .ZN(G1345gat));
  NOR3_X1   g713(.A1(new_n884), .A2(new_n234), .A3(new_n568), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n891), .A2(new_n569), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  AOI21_X1  g716(.A(G155gat), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n891), .A2(KEYINPUT122), .A3(new_n569), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1346gat));
  NOR2_X1   g719(.A1(new_n619), .A2(G162gat), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n891), .A2(KEYINPUT123), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT123), .B1(new_n891), .B2(new_n921), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(new_n884), .B2(new_n619), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(G162gat), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n884), .A2(new_n924), .A3(new_n619), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n922), .A2(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n752), .A2(new_n460), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n851), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(new_n326), .A3(new_n748), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n849), .A2(new_n670), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n520), .A2(new_n471), .A3(new_n460), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n667), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n931), .B1(new_n326), .B2(new_n936), .ZN(G1348gat));
  NOR3_X1   g736(.A1(new_n930), .A2(new_n327), .A3(new_n640), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n747), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n327), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n942), .A3(new_n327), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n938), .B1(new_n941), .B2(new_n943), .ZN(G1349gat));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(KEYINPUT60), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n945), .A2(KEYINPUT60), .ZN(new_n947));
  OAI21_X1  g746(.A(G183gat), .B1(new_n930), .B2(new_n568), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n374), .A2(new_n376), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n932), .A2(new_n949), .A3(new_n569), .A4(new_n933), .ZN(new_n950));
  AOI211_X1 g749(.A(new_n946), .B(new_n947), .C1(new_n948), .C2(new_n950), .ZN(new_n951));
  AND4_X1   g750(.A1(new_n945), .A2(new_n948), .A3(KEYINPUT60), .A4(new_n950), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n935), .A2(new_n340), .A3(new_n704), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n851), .A2(new_n704), .A3(new_n929), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n955), .A2(new_n956), .A3(G190gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n955), .B2(G190gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  NAND2_X1  g758(.A1(new_n929), .A2(new_n685), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n908), .A2(new_n961), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n962), .A2(new_n203), .A3(new_n748), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n686), .A2(new_n285), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n932), .A2(new_n413), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n667), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n963), .A2(new_n966), .ZN(G1352gat));
  NAND4_X1  g766(.A1(new_n932), .A2(new_n204), .A3(new_n782), .A4(new_n964), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT62), .Z(new_n969));
  AND3_X1   g768(.A1(new_n908), .A2(new_n747), .A3(new_n961), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n204), .B2(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n965), .A2(new_n211), .A3(new_n569), .ZN(new_n972));
  NOR2_X1   g771(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n973));
  OAI211_X1 g772(.A(G211gat), .B(new_n973), .C1(new_n962), .C2(new_n568), .ZN(new_n974));
  INV_X1    g773(.A(new_n962), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n211), .B1(new_n975), .B2(new_n569), .ZN(new_n976));
  XNOR2_X1  g775(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n972), .B(new_n974), .C1(new_n976), .C2(new_n977), .ZN(G1354gat));
  OAI21_X1  g777(.A(G218gat), .B1(new_n962), .B2(new_n619), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n965), .A2(new_n212), .A3(new_n704), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1355gat));
endmodule


