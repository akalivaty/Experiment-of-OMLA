

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  INV_X1 U323 ( .A(n522), .ZN(n524) );
  XNOR2_X1 U324 ( .A(n407), .B(n342), .ZN(n343) );
  XNOR2_X1 U325 ( .A(n391), .B(KEYINPUT48), .ZN(n522) );
  XNOR2_X1 U326 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n444) );
  INV_X1 U327 ( .A(n376), .ZN(n342) );
  XNOR2_X1 U328 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U329 ( .A(n344), .B(n343), .ZN(n386) );
  XOR2_X1 U330 ( .A(n466), .B(KEYINPUT28), .Z(n528) );
  XNOR2_X1 U331 ( .A(KEYINPUT89), .B(n464), .ZN(n570) );
  XNOR2_X1 U332 ( .A(n449), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U333 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  INV_X1 U334 ( .A(KEYINPUT121), .ZN(n448) );
  XOR2_X1 U335 ( .A(G71GAT), .B(G120GAT), .Z(n292) );
  XNOR2_X1 U336 ( .A(G127GAT), .B(KEYINPUT20), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U338 ( .A(G183GAT), .B(KEYINPUT81), .Z(n294) );
  XNOR2_X1 U339 ( .A(G15GAT), .B(KEYINPUT80), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U341 ( .A(n296), .B(n295), .Z(n301) );
  XOR2_X1 U342 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n298) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U345 ( .A(G176GAT), .B(n299), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n307) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G190GAT), .Z(n305) );
  XOR2_X1 U348 ( .A(KEYINPUT0), .B(KEYINPUT79), .Z(n303) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n431) );
  XNOR2_X1 U351 ( .A(G134GAT), .B(n431), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(n307), .B(n306), .Z(n312) );
  XOR2_X1 U354 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n309) );
  XNOR2_X1 U355 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U357 ( .A(G169GAT), .B(n310), .Z(n403) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(n403), .ZN(n311) );
  XOR2_X1 U359 ( .A(n312), .B(n311), .Z(n468) );
  INV_X1 U360 ( .A(n468), .ZN(n526) );
  XOR2_X1 U361 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n314) );
  XNOR2_X1 U362 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U364 ( .A(G8GAT), .B(G183GAT), .Z(n394) );
  XOR2_X1 U365 ( .A(n394), .B(G78GAT), .Z(n316) );
  XOR2_X1 U366 ( .A(G22GAT), .B(G15GAT), .Z(n360) );
  XNOR2_X1 U367 ( .A(n360), .B(G211GAT), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U369 ( .A(n318), .B(n317), .Z(n320) );
  NAND2_X1 U370 ( .A1(G231GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U372 ( .A(KEYINPUT73), .B(KEYINPUT76), .Z(n322) );
  XNOR2_X1 U373 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U375 ( .A(n324), .B(n323), .Z(n329) );
  XNOR2_X1 U376 ( .A(G1GAT), .B(G127GAT), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n325), .B(G155GAT), .ZN(n436) );
  XOR2_X1 U378 ( .A(KEYINPUT69), .B(KEYINPUT13), .Z(n327) );
  XNOR2_X1 U379 ( .A(G71GAT), .B(G57GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n436), .B(n332), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n578) );
  XOR2_X1 U383 ( .A(n578), .B(KEYINPUT109), .Z(n564) );
  XOR2_X1 U384 ( .A(G64GAT), .B(G92GAT), .Z(n331) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n399) );
  XNOR2_X1 U387 ( .A(n399), .B(n332), .ZN(n334) );
  INV_X1 U388 ( .A(KEYINPUT71), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n339) );
  XOR2_X1 U390 ( .A(KEYINPUT70), .B(KEYINPUT32), .Z(n336) );
  NAND2_X1 U391 ( .A1(G230GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(n337), .B(KEYINPUT33), .Z(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U395 ( .A(G120GAT), .B(G148GAT), .Z(n434) );
  XNOR2_X1 U396 ( .A(n434), .B(KEYINPUT31), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n344) );
  XOR2_X1 U398 ( .A(G106GAT), .B(G78GAT), .Z(n407) );
  XNOR2_X1 U399 ( .A(G99GAT), .B(G85GAT), .ZN(n376) );
  XOR2_X1 U400 ( .A(KEYINPUT41), .B(n386), .Z(n547) );
  XOR2_X1 U401 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n346) );
  XNOR2_X1 U402 ( .A(G8GAT), .B(KEYINPUT64), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n358) );
  XOR2_X1 U404 ( .A(G197GAT), .B(G50GAT), .Z(n348) );
  XNOR2_X1 U405 ( .A(G36GAT), .B(G29GAT), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n356) );
  XOR2_X1 U407 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n350) );
  XNOR2_X1 U408 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U410 ( .A(G1GAT), .B(G113GAT), .Z(n352) );
  XNOR2_X1 U411 ( .A(G169GAT), .B(G141GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U413 ( .A(n354), .B(n353), .Z(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n364) );
  XNOR2_X1 U416 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n359), .B(KEYINPUT7), .ZN(n377) );
  XOR2_X1 U418 ( .A(n377), .B(n360), .Z(n362) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U421 ( .A(n364), .B(n363), .Z(n529) );
  INV_X1 U422 ( .A(n529), .ZN(n573) );
  AND2_X1 U423 ( .A1(n547), .A2(n573), .ZN(n366) );
  XNOR2_X1 U424 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  NOR2_X1 U426 ( .A1(n564), .A2(n367), .ZN(n382) );
  XOR2_X1 U427 ( .A(KEYINPUT72), .B(KEYINPUT10), .Z(n369) );
  XNOR2_X1 U428 ( .A(G106GAT), .B(G162GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n381) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n371) );
  NAND2_X1 U431 ( .A1(G232GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U433 ( .A(n372), .B(G92GAT), .Z(n374) );
  XOR2_X1 U434 ( .A(G50GAT), .B(G218GAT), .Z(n408) );
  XOR2_X1 U435 ( .A(G29GAT), .B(G134GAT), .Z(n437) );
  XNOR2_X1 U436 ( .A(n408), .B(n437), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U438 ( .A(G36GAT), .B(G190GAT), .Z(n396) );
  XOR2_X1 U439 ( .A(n375), .B(n396), .Z(n379) );
  XOR2_X1 U440 ( .A(n377), .B(n376), .Z(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n551) );
  INV_X1 U443 ( .A(n551), .ZN(n453) );
  NAND2_X1 U444 ( .A1(n382), .A2(n453), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n383), .B(KEYINPUT47), .ZN(n390) );
  XOR2_X1 U446 ( .A(KEYINPUT36), .B(n453), .Z(n580) );
  NAND2_X1 U447 ( .A1(n578), .A2(n580), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n384), .B(KEYINPUT111), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n385), .B(KEYINPUT45), .ZN(n387) );
  INV_X1 U450 ( .A(n386), .ZN(n452) );
  NAND2_X1 U451 ( .A1(n387), .A2(n452), .ZN(n388) );
  NOR2_X1 U452 ( .A1(n573), .A2(n388), .ZN(n389) );
  NOR2_X1 U453 ( .A1(n390), .A2(n389), .ZN(n391) );
  XOR2_X1 U454 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n393) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U457 ( .A(n395), .B(n394), .Z(n398) );
  XNOR2_X1 U458 ( .A(G218GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U460 ( .A(n400), .B(n399), .Z(n405) );
  XOR2_X1 U461 ( .A(G211GAT), .B(KEYINPUT21), .Z(n402) );
  XNOR2_X1 U462 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n403), .B(n412), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n513) );
  NOR2_X1 U466 ( .A1(n522), .A2(n513), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n406), .B(KEYINPUT54), .ZN(n569) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n411) );
  XOR2_X1 U469 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n410) );
  XNOR2_X1 U470 ( .A(G141GAT), .B(G162GAT), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n430) );
  XNOR2_X1 U472 ( .A(n411), .B(n430), .ZN(n416) );
  XOR2_X1 U473 ( .A(G22GAT), .B(n412), .Z(n414) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U476 ( .A(n416), .B(n415), .Z(n424) );
  XOR2_X1 U477 ( .A(KEYINPUT85), .B(KEYINPUT87), .Z(n418) );
  XNOR2_X1 U478 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U480 ( .A(G148GAT), .B(G155GAT), .Z(n420) );
  XNOR2_X1 U481 ( .A(KEYINPUT24), .B(G204GAT), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n466) );
  XOR2_X1 U485 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n426) );
  XNOR2_X1 U486 ( .A(G85GAT), .B(KEYINPUT1), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n441) );
  XOR2_X1 U488 ( .A(KEYINPUT6), .B(KEYINPUT88), .Z(n428) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U491 ( .A(n429), .B(G57GAT), .Z(n433) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U494 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U497 ( .A(n441), .B(n440), .Z(n464) );
  INV_X1 U498 ( .A(n570), .ZN(n442) );
  NOR2_X1 U499 ( .A1(n466), .A2(n442), .ZN(n443) );
  AND2_X1 U500 ( .A1(n569), .A2(n443), .ZN(n445) );
  NOR2_X1 U501 ( .A1(n526), .A2(n446), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n565) );
  NAND2_X1 U503 ( .A1(n565), .A2(n551), .ZN(n451) );
  XOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n449) );
  NAND2_X1 U505 ( .A1(n573), .A2(n452), .ZN(n485) );
  XOR2_X1 U506 ( .A(KEYINPUT16), .B(KEYINPUT77), .Z(n455) );
  NAND2_X1 U507 ( .A1(n578), .A2(n453), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n472) );
  NOR2_X1 U509 ( .A1(n526), .A2(n513), .ZN(n456) );
  XOR2_X1 U510 ( .A(KEYINPUT93), .B(n456), .Z(n457) );
  NOR2_X1 U511 ( .A1(n466), .A2(n457), .ZN(n458) );
  XOR2_X1 U512 ( .A(KEYINPUT94), .B(n458), .Z(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT25), .ZN(n462) );
  XNOR2_X1 U514 ( .A(n513), .B(KEYINPUT27), .ZN(n465) );
  NAND2_X1 U515 ( .A1(n466), .A2(n526), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT26), .ZN(n572) );
  NOR2_X1 U517 ( .A1(n465), .A2(n572), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n471) );
  NOR2_X1 U520 ( .A1(n570), .A2(n465), .ZN(n523) );
  NAND2_X1 U521 ( .A1(n523), .A2(n528), .ZN(n467) );
  XNOR2_X1 U522 ( .A(KEYINPUT92), .B(n467), .ZN(n469) );
  NOR2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U524 ( .A1(n471), .A2(n470), .ZN(n482) );
  NOR2_X1 U525 ( .A1(n472), .A2(n482), .ZN(n473) );
  XNOR2_X1 U526 ( .A(n473), .B(KEYINPUT95), .ZN(n499) );
  OR2_X1 U527 ( .A1(n485), .A2(n499), .ZN(n479) );
  NOR2_X1 U528 ( .A1(n570), .A2(n479), .ZN(n474) );
  XOR2_X1 U529 ( .A(G1GAT), .B(n474), .Z(n475) );
  XNOR2_X1 U530 ( .A(KEYINPUT34), .B(n475), .ZN(G1324GAT) );
  NOR2_X1 U531 ( .A1(n513), .A2(n479), .ZN(n476) );
  XOR2_X1 U532 ( .A(G8GAT), .B(n476), .Z(G1325GAT) );
  NOR2_X1 U533 ( .A1(n526), .A2(n479), .ZN(n478) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NOR2_X1 U536 ( .A1(n528), .A2(n479), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT96), .B(n480), .Z(n481) );
  XNOR2_X1 U538 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  NOR2_X1 U539 ( .A1(n578), .A2(n482), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n580), .A2(n483), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT37), .B(n484), .Z(n509) );
  NOR2_X1 U542 ( .A1(n509), .A2(n485), .ZN(n487) );
  XNOR2_X1 U543 ( .A(KEYINPUT97), .B(KEYINPUT38), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(n494) );
  NOR2_X1 U545 ( .A1(n494), .A2(n570), .ZN(n489) );
  XNOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NOR2_X1 U548 ( .A1(n513), .A2(n494), .ZN(n490) );
  XOR2_X1 U549 ( .A(G36GAT), .B(n490), .Z(G1329GAT) );
  XNOR2_X1 U550 ( .A(KEYINPUT98), .B(KEYINPUT40), .ZN(n492) );
  NOR2_X1 U551 ( .A1(n526), .A2(n494), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U553 ( .A(G43GAT), .B(n493), .Z(G1330GAT) );
  XNOR2_X1 U554 ( .A(G50GAT), .B(KEYINPUT99), .ZN(n496) );
  NOR2_X1 U555 ( .A1(n528), .A2(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1331GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n498) );
  XNOR2_X1 U558 ( .A(G57GAT), .B(KEYINPUT101), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n547), .B(KEYINPUT100), .ZN(n561) );
  NAND2_X1 U561 ( .A1(n529), .A2(n561), .ZN(n508) );
  OR2_X1 U562 ( .A1(n508), .A2(n499), .ZN(n504) );
  NOR2_X1 U563 ( .A1(n570), .A2(n504), .ZN(n500) );
  XOR2_X1 U564 ( .A(n501), .B(n500), .Z(G1332GAT) );
  NOR2_X1 U565 ( .A1(n513), .A2(n504), .ZN(n502) );
  XOR2_X1 U566 ( .A(G64GAT), .B(n502), .Z(G1333GAT) );
  NOR2_X1 U567 ( .A1(n526), .A2(n504), .ZN(n503) );
  XOR2_X1 U568 ( .A(G71GAT), .B(n503), .Z(G1334GAT) );
  NOR2_X1 U569 ( .A1(n528), .A2(n504), .ZN(n506) );
  XNOR2_X1 U570 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U572 ( .A(G78GAT), .B(n507), .Z(G1335GAT) );
  NOR2_X1 U573 ( .A1(n509), .A2(n508), .ZN(n510) );
  XOR2_X1 U574 ( .A(KEYINPUT104), .B(n510), .Z(n518) );
  NOR2_X1 U575 ( .A1(n518), .A2(n570), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT105), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NOR2_X1 U578 ( .A1(n513), .A2(n518), .ZN(n514) );
  XOR2_X1 U579 ( .A(KEYINPUT106), .B(n514), .Z(n515) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(n515), .ZN(G1337GAT) );
  XNOR2_X1 U581 ( .A(G99GAT), .B(KEYINPUT107), .ZN(n517) );
  NOR2_X1 U582 ( .A1(n526), .A2(n518), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1338GAT) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT108), .ZN(n520) );
  NOR2_X1 U585 ( .A1(n528), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U587 ( .A(G106GAT), .B(n521), .Z(G1339GAT) );
  NAND2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT112), .B(n525), .ZN(n541) );
  NOR2_X1 U590 ( .A1(n526), .A2(n541), .ZN(n527) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n532) );
  NOR2_X1 U592 ( .A1(n529), .A2(n532), .ZN(n531) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n534) );
  INV_X1 U596 ( .A(n532), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n538), .A2(n561), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n536) );
  NAND2_X1 U600 ( .A1(n538), .A2(n564), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U602 ( .A(G127GAT), .B(n537), .Z(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U604 ( .A1(n538), .A2(n551), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  XOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT115), .Z(n543) );
  NOR2_X1 U607 ( .A1(n572), .A2(n541), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n552), .A2(n573), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n545) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U613 ( .A(KEYINPUT52), .B(n546), .Z(n549) );
  NAND2_X1 U614 ( .A1(n552), .A2(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n552), .A2(n578), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n554) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n573), .A2(n565), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT122), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n559) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(n560), .Z(n563) );
  NAND2_X1 U629 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT60), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(n568), .Z(n575) );
  NAND2_X1 U636 ( .A1(n569), .A2(n570), .ZN(n571) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n581), .A2(n386), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n583) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

