//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  OR3_X1    g0020(.A1(new_n209), .A2(KEYINPUT64), .A3(G13), .ZN(new_n221));
  OAI21_X1  g0021(.A(KEYINPUT64), .B1(new_n209), .B2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n207), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n220), .B(new_n225), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G226), .B(G232), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n211), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n242), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n226), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n251), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n206), .A2(G20), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n257), .A2(G68), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n206), .A2(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n211), .A2(G20), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT12), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n254), .A2(new_n211), .A3(new_n256), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(KEYINPUT12), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT72), .ZN(new_n265));
  OR3_X1    g0065(.A1(new_n259), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n259), .B2(new_n264), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n207), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n261), .B1(new_n268), .B2(new_n269), .C1(new_n271), .C2(new_n243), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n251), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT11), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n266), .A2(new_n267), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT14), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT71), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n202), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n280), .B2(KEYINPUT71), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT70), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G226), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n287), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n279), .A2(KEYINPUT70), .A3(G226), .A4(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n283), .A2(new_n286), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G274), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  INV_X1    g0102(.A(G45), .ZN(new_n303));
  AOI21_X1  g0103(.A(G1), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n304), .ZN(new_n306));
  OAI211_X1 g0106(.A(G1), .B(G13), .C1(new_n284), .C2(new_n302), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n305), .B1(new_n212), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n278), .B1(new_n299), .B2(new_n310), .ZN(new_n311));
  AOI211_X1 g0111(.A(KEYINPUT13), .B(new_n309), .C1(new_n297), .C2(new_n298), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n277), .B(G169), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n281), .A2(new_n282), .B1(new_n294), .B2(new_n295), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n307), .B1(new_n314), .B2(new_n286), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT13), .B1(new_n315), .B2(new_n309), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n299), .A2(new_n278), .A3(new_n310), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(G179), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n277), .B1(new_n320), .B2(G169), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n276), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G226), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n305), .B1(new_n323), .B2(new_n308), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n279), .A2(G222), .A3(new_n292), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n279), .A2(G1698), .ZN(new_n326));
  INV_X1    g0126(.A(G223), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n325), .B1(new_n269), .B2(new_n279), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT67), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n307), .B1(new_n328), .B2(KEYINPUT67), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n324), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT8), .B(G58), .ZN(new_n332));
  INV_X1    g0132(.A(G150), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n332), .A2(new_n268), .B1(new_n333), .B2(new_n271), .ZN(new_n334));
  NOR2_X1   g0134(.A1(G58), .A2(G68), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n207), .B1(new_n335), .B2(new_n243), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n251), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n253), .A2(new_n251), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n258), .A2(G50), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n340), .A2(new_n341), .B1(G50), .B2(new_n252), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n331), .A2(G169), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n331), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n338), .A2(new_n342), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT9), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(KEYINPUT9), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n348), .C1(new_n331), .C2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n331), .A2(G190), .ZN(new_n351));
  OR3_X1    g0151(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT10), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT10), .B1(new_n350), .B2(new_n351), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n345), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(G200), .B1(new_n311), .B2(new_n312), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n316), .A2(new_n317), .A3(G190), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n275), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n251), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n332), .B(KEYINPUT68), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n270), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n361), .A2(new_n268), .B1(new_n207), .B2(new_n269), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n358), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n257), .A2(G77), .A3(new_n258), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n254), .A2(new_n256), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(G77), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n279), .A2(G232), .A3(new_n292), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n369), .B1(new_n203), .B2(new_n279), .C1(new_n326), .C2(new_n212), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n298), .ZN(new_n371));
  INV_X1    g0171(.A(new_n308), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G244), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n305), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n374), .A2(G179), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n368), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n374), .A2(G200), .ZN(new_n381));
  INV_X1    g0181(.A(G190), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n374), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  AND4_X1   g0184(.A1(new_n322), .A2(new_n354), .A3(new_n357), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT76), .ZN(new_n386));
  INV_X1    g0186(.A(G232), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n305), .B1(new_n387), .B2(new_n308), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n279), .A2(G223), .A3(new_n292), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n389), .B1(new_n284), .B2(new_n213), .C1(new_n326), .C2(new_n323), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n388), .B1(new_n390), .B2(new_n298), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n391), .A2(G179), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n375), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n386), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(G179), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n395), .B(KEYINPUT76), .C1(new_n375), .C2(new_n391), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G58), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(new_n211), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n399), .B2(new_n335), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n270), .A2(G159), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n279), .A2(new_n405), .A3(G20), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n289), .A2(G33), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT73), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT73), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n288), .A2(new_n290), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n207), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n405), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n406), .B1(new_n413), .B2(KEYINPUT74), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n415), .A3(new_n405), .ZN(new_n416));
  AOI211_X1 g0216(.A(KEYINPUT75), .B(new_n211), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT75), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n288), .A2(new_n290), .A3(new_n410), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n410), .B1(new_n288), .B2(new_n290), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n419), .A2(new_n420), .A3(G20), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT74), .B1(new_n421), .B2(KEYINPUT7), .ZN(new_n422));
  INV_X1    g0222(.A(new_n406), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n416), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n418), .B1(new_n424), .B2(G68), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n404), .B1(new_n417), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n402), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT7), .B1(new_n291), .B2(new_n207), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n406), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(new_n211), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n403), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n251), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n332), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n258), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n340), .A2(new_n434), .B1(new_n252), .B2(new_n433), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  AOI211_X1 g0236(.A(KEYINPUT18), .B(new_n397), .C1(new_n432), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(new_n436), .ZN(new_n439));
  INV_X1    g0239(.A(new_n397), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n391), .A2(new_n382), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G200), .B2(new_n391), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n432), .A2(new_n436), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT17), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n432), .A2(KEYINPUT17), .A3(new_n436), .A4(new_n444), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n385), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n279), .A2(new_n207), .A3(G68), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT19), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n268), .B2(new_n202), .ZN(new_n454));
  AOI21_X1  g0254(.A(G20), .B1(new_n285), .B2(KEYINPUT19), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n204), .A2(G87), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n452), .B(new_n454), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n251), .ZN(new_n458));
  INV_X1    g0258(.A(new_n366), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n361), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n339), .B1(G1), .B2(new_n284), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n458), .B(new_n460), .C1(new_n461), .C2(new_n361), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n303), .A2(G1), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n214), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n307), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n307), .A2(G274), .ZN(new_n466));
  INV_X1    g0266(.A(new_n463), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n279), .A2(G244), .A3(G1698), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n279), .A2(G238), .A3(new_n292), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G116), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n468), .B1(new_n298), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n344), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n462), .B(new_n474), .C1(G169), .C2(new_n473), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n339), .B(G87), .C1(G1), .C2(new_n284), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n458), .A2(new_n460), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(new_n298), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n301), .A2(new_n463), .B1(new_n307), .B2(new_n464), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G200), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n473), .A2(G190), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n477), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n288), .A2(new_n290), .A3(new_n207), .A4(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT22), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n279), .A2(new_n487), .A3(new_n207), .A4(G87), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT24), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n471), .A2(G20), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n207), .B2(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n489), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n490), .B1(new_n489), .B2(new_n495), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n251), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n253), .A2(new_n203), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT25), .ZN(new_n500));
  INV_X1    g0300(.A(new_n461), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(G107), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n279), .A2(G257), .A3(G1698), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G294), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n288), .A2(new_n290), .A3(G250), .A4(new_n292), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g0308(.A(KEYINPUT5), .B(G41), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n298), .B1(new_n463), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n508), .A2(new_n298), .B1(G264), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n509), .A2(new_n463), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n301), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(new_n382), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(G200), .B2(new_n514), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n484), .B1(new_n504), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n509), .A2(new_n463), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(G257), .A3(new_n307), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT80), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT80), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n510), .A2(new_n521), .A3(G257), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n520), .A2(new_n522), .B1(new_n301), .B2(new_n512), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n288), .A2(new_n290), .A3(G244), .A4(new_n292), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(KEYINPUT79), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n288), .A2(new_n290), .A3(G250), .A4(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(new_n524), .C2(new_n525), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT79), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n524), .B2(new_n525), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n527), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n523), .B1(new_n533), .B2(new_n307), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n270), .A2(G77), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT77), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n539), .A2(new_n202), .A3(G107), .ZN(new_n540));
  XNOR2_X1  g0340(.A(G97), .B(G107), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n538), .B1(new_n543), .B2(G20), .ZN(new_n544));
  OAI21_X1  g0344(.A(G107), .B1(new_n406), .B2(new_n428), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n358), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n252), .A2(G97), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n461), .B2(new_n202), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT78), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n526), .A2(KEYINPUT79), .ZN(new_n551));
  OR2_X1    g0351(.A1(new_n524), .A2(new_n525), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n528), .A2(new_n529), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n298), .B1(new_n554), .B2(new_n527), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(G190), .A3(new_n523), .ZN(new_n556));
  INV_X1    g0356(.A(new_n545), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n536), .B(KEYINPUT77), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n207), .B2(new_n542), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n251), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT78), .ZN(new_n561));
  INV_X1    g0361(.A(new_n549), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n535), .A2(new_n550), .A3(new_n556), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n534), .A2(G169), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n555), .A2(G179), .A3(new_n523), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n546), .A2(new_n549), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT81), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT81), .ZN(new_n571));
  AOI211_X1 g0371(.A(new_n571), .B(new_n568), .C1(new_n565), .C2(new_n566), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n517), .B(new_n564), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n508), .A2(new_n298), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n510), .A2(G264), .ZN(new_n575));
  AND4_X1   g0375(.A1(new_n344), .A2(new_n574), .A3(new_n513), .A4(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(G169), .B1(new_n511), .B2(new_n513), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n578), .A2(new_n503), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n579), .B1(new_n578), .B2(new_n503), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(G116), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n206), .B2(G33), .ZN(new_n585));
  INV_X1    g0385(.A(new_n256), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n252), .A2(new_n255), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n358), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G116), .B2(new_n366), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n529), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT83), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n284), .A2(G97), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT83), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n207), .A4(new_n529), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n584), .A2(G20), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n251), .A2(KEYINPUT82), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n251), .A2(new_n596), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT82), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n251), .A2(KEYINPUT82), .A3(new_n596), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT82), .B1(new_n251), .B2(new_n596), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(KEYINPUT20), .A3(new_n595), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n589), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n510), .A2(G270), .B1(new_n512), .B2(new_n301), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n288), .A2(new_n290), .A3(G264), .A4(G1698), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n288), .A2(new_n290), .A3(G257), .A4(new_n292), .ZN(new_n611));
  INV_X1    g0411(.A(G303), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n279), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n298), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n608), .B(new_n616), .C1(new_n382), .C2(new_n615), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(G169), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n608), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n459), .A2(new_n584), .B1(new_n257), .B2(new_n585), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n601), .A2(new_n602), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT20), .B1(new_n606), .B2(new_n595), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n613), .A2(new_n298), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n518), .A2(G270), .A3(new_n307), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n513), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n624), .A2(G179), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n375), .B1(new_n609), .B2(new_n614), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n624), .A2(KEYINPUT21), .A3(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n617), .A2(new_n620), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  NOR4_X1   g0432(.A1(new_n451), .A2(new_n573), .A3(new_n583), .A4(new_n632), .ZN(G372));
  NOR2_X1   g0433(.A1(new_n377), .A2(new_n378), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n357), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n322), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n449), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n392), .A2(new_n393), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n432), .B2(new_n436), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT18), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n352), .A2(new_n353), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n345), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n475), .A2(new_n483), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n550), .A2(new_n563), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n644), .A2(new_n645), .A3(new_n567), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n475), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n555), .A2(G179), .A3(new_n523), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n375), .B1(new_n555), .B2(new_n523), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n569), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n571), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n567), .A2(KEYINPUT81), .A3(new_n569), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n644), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n648), .B1(KEYINPUT26), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n564), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n652), .B2(new_n653), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n578), .A2(new_n503), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n620), .A2(new_n631), .A3(new_n629), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT85), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n620), .A2(new_n629), .A3(new_n631), .A4(KEYINPUT85), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT86), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n657), .B(new_n517), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n655), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n643), .B1(new_n451), .B2(new_n669), .ZN(G369));
  OR2_X1    g0470(.A1(new_n632), .A2(KEYINPUT87), .ZN(new_n671));
  OR3_X1    g0471(.A1(new_n260), .A2(KEYINPUT27), .A3(G20), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT27), .B1(new_n260), .B2(G20), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n608), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n632), .B2(KEYINPUT87), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n662), .A2(new_n663), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n671), .A2(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n516), .A2(new_n504), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n582), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n504), .A2(new_n677), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n685), .A2(new_n686), .B1(new_n658), .B2(new_n677), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n660), .A2(new_n677), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n659), .B2(new_n677), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n223), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n456), .A2(new_n584), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n694), .A2(new_n206), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n228), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  NOR3_X1   g0499(.A1(new_n632), .A2(new_n580), .A3(new_n581), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n657), .A2(new_n517), .A3(new_n700), .A4(new_n677), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n628), .A2(G179), .A3(new_n473), .A4(new_n511), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n534), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n478), .A2(new_n574), .A3(new_n479), .A4(new_n575), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n609), .A2(G179), .A3(new_n614), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(KEYINPUT30), .A3(new_n555), .A4(new_n523), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n473), .A2(G179), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n534), .A2(new_n514), .A3(new_n615), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n704), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT88), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n704), .A2(new_n708), .A3(KEYINPUT88), .A4(new_n710), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n676), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n701), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT89), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT89), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n722), .A3(G330), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n668), .A2(new_n677), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT29), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n583), .A2(new_n660), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n573), .ZN(new_n728));
  INV_X1    g0528(.A(new_n475), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n644), .A2(new_n567), .A3(new_n646), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(KEYINPUT26), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n652), .A2(new_n653), .A3(new_n645), .A4(new_n644), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(KEYINPUT29), .B(new_n677), .C1(new_n728), .C2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n724), .B1(new_n726), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n699), .B1(new_n735), .B2(G1), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT90), .Z(G364));
  AOI21_X1  g0537(.A(new_n226), .B1(G20), .B2(new_n375), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n344), .A2(G200), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G20), .A3(G190), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n279), .B1(new_n742), .B2(G322), .ZN(new_n743));
  INV_X1    g0543(.A(G311), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n207), .A2(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n740), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n207), .A2(new_n344), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n382), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(KEYINPUT33), .A2(G317), .ZN(new_n751));
  AND2_X1   g0551(.A1(KEYINPUT33), .A2(G317), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G283), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n207), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(new_n382), .A3(G200), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n753), .B1(new_n754), .B2(new_n756), .C1(new_n612), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n344), .A2(new_n349), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT93), .ZN(new_n760));
  INV_X1    g0560(.A(new_n745), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n747), .B(new_n758), .C1(G329), .C2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n745), .B1(new_n760), .B2(G20), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT94), .ZN(new_n766));
  INV_X1    g0566(.A(G326), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n748), .A2(G190), .A3(G200), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT95), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n763), .B1(new_n764), .B2(new_n766), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n766), .A2(new_n202), .ZN(new_n771));
  INV_X1    g0571(.A(new_n762), .ZN(new_n772));
  INV_X1    g0572(.A(G159), .ZN(new_n773));
  OR3_X1    g0573(.A1(new_n772), .A2(KEYINPUT32), .A3(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n741), .A2(new_n398), .B1(new_n746), .B2(new_n269), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT92), .Z(new_n776));
  OAI22_X1  g0576(.A1(new_n749), .A2(new_n211), .B1(new_n756), .B2(new_n203), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n279), .B1(new_n768), .B2(new_n243), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n757), .A2(new_n213), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT32), .B1(new_n772), .B2(new_n773), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n774), .A2(new_n776), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n770), .B1(new_n771), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT96), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n739), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n207), .A2(G13), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n206), .B1(new_n787), .B2(G45), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n223), .A2(G355), .A3(new_n279), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n419), .A2(new_n420), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n693), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n229), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(G45), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n248), .A2(new_n303), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n790), .B1(G116), .B2(new_n223), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n738), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n694), .B(new_n789), .C1(new_n797), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n800), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n786), .B(new_n802), .C1(new_n681), .C2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT97), .Z(new_n805));
  NOR2_X1   g0605(.A1(new_n681), .A2(G330), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n694), .A2(new_n789), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n683), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT91), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n808), .A2(KEYINPUT91), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n805), .A2(new_n809), .A3(new_n810), .ZN(G396));
  INV_X1    g0611(.A(new_n724), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n379), .A2(KEYINPUT101), .ZN(new_n813));
  OR3_X1    g0613(.A1(new_n377), .A2(KEYINPUT101), .A3(new_n378), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n815), .A2(new_n383), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n668), .A2(new_n677), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n368), .A2(new_n676), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n813), .A2(new_n383), .A3(new_n818), .A4(new_n814), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n379), .B2(new_n677), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n817), .B1(new_n725), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n807), .B1(new_n812), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n812), .B2(new_n821), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n739), .A2(new_n799), .ZN(new_n824));
  INV_X1    g0624(.A(new_n746), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n742), .A2(G143), .B1(new_n825), .B2(G159), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n827), .B2(new_n768), .C1(new_n333), .C2(new_n749), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT98), .Z(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n243), .A2(new_n757), .B1(new_n756), .B2(new_n211), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT99), .Z(new_n832));
  AOI21_X1  g0632(.A(new_n791), .B1(new_n762), .B2(G132), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n766), .C2(new_n398), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n291), .B1(new_n746), .B2(new_n584), .C1(new_n764), .C2(new_n741), .ZN(new_n837));
  INV_X1    g0637(.A(new_n757), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G283), .A2(new_n750), .B1(new_n838), .B2(G107), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n839), .B1(new_n213), .B2(new_n756), .C1(new_n612), .C2(new_n768), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n837), .B(new_n840), .C1(G311), .C2(new_n762), .ZN(new_n841));
  INV_X1    g0641(.A(new_n771), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n835), .A2(new_n836), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n807), .B1(G77), .B2(new_n824), .C1(new_n843), .C2(new_n739), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT100), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n799), .B2(new_n820), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n823), .A2(new_n846), .ZN(G384));
  NOR2_X1   g0647(.A1(new_n275), .A2(new_n677), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n322), .A2(new_n357), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(G169), .B1(new_n311), .B2(new_n312), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT14), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n357), .A2(new_n852), .A3(new_n318), .A4(new_n313), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n848), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n850), .A2(new_n854), .A3(KEYINPUT102), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT102), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n322), .A2(new_n856), .A3(new_n357), .A4(new_n849), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT103), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT103), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n855), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n676), .A4(new_n714), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n701), .A2(new_n717), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n820), .ZN(new_n865));
  NAND2_X1  g0665(.A1(KEYINPUT104), .A2(KEYINPUT40), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n412), .A2(new_n415), .A3(new_n405), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n415), .B1(new_n412), .B2(new_n405), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n868), .A2(new_n869), .A3(new_n406), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT75), .B1(new_n870), .B2(new_n211), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n424), .A2(new_n418), .A3(G68), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n358), .B1(new_n873), .B2(new_n404), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n427), .B1(new_n417), .B2(new_n425), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n403), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n435), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n445), .B1(new_n877), .B2(new_n638), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n674), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT37), .B1(new_n439), .B2(new_n440), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n674), .B1(new_n432), .B2(new_n436), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n445), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n435), .B1(new_n874), .B2(new_n431), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT18), .B1(new_n886), .B2(new_n397), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n439), .A2(new_n438), .A3(new_n440), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(new_n447), .A3(new_n448), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n879), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n885), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n885), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n867), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n861), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n860), .B1(new_n855), .B2(new_n857), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n865), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT104), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n883), .B1(new_n640), .B2(new_n449), .ZN(new_n901));
  INV_X1    g0701(.A(new_n638), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n439), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n883), .A2(new_n445), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n445), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(new_n882), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n904), .A2(KEYINPUT37), .B1(new_n906), .B2(new_n881), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n900), .B1(new_n901), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n885), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n894), .B1(new_n899), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n895), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n450), .A2(new_n864), .ZN(new_n913));
  OAI21_X1  g0713(.A(G330), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n913), .B2(new_n912), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n903), .A2(KEYINPUT18), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n639), .A2(new_n438), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n917), .A2(new_n447), .A3(new_n448), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n882), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n905), .A2(new_n639), .A3(new_n882), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT37), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n884), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n916), .B1(new_n891), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT16), .B1(new_n873), .B2(new_n427), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n426), .A2(new_n251), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n436), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n674), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n445), .C1(new_n638), .C2(new_n877), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(KEYINPUT37), .B1(new_n906), .B2(new_n881), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n930), .B1(new_n442), .B2(new_n449), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n900), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(KEYINPUT39), .A3(new_n909), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n322), .A2(new_n676), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n925), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n640), .A2(new_n929), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n934), .A2(new_n909), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n815), .A2(new_n676), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n817), .A2(new_n941), .B1(new_n859), .B2(new_n861), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n450), .B(new_n734), .C1(new_n725), .C2(KEYINPUT29), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n643), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n944), .B(new_n946), .Z(new_n947));
  OAI22_X1  g0747(.A1(new_n915), .A2(new_n947), .B1(new_n206), .B2(new_n787), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n947), .B2(new_n915), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n543), .A2(KEYINPUT35), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n543), .A2(KEYINPUT35), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n950), .A2(G116), .A3(new_n227), .A4(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT36), .Z(new_n953));
  OAI211_X1 g0753(.A(new_n697), .B(G77), .C1(new_n398), .C2(new_n211), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n206), .B(G13), .C1(new_n954), .C2(new_n244), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n949), .A2(new_n953), .A3(new_n955), .ZN(G367));
  OAI22_X1  g0756(.A1(new_n749), .A2(new_n764), .B1(new_n756), .B2(new_n202), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n791), .B1(new_n754), .B2(new_n746), .C1(new_n612), .C2(new_n741), .ZN(new_n958));
  INV_X1    g0758(.A(new_n769), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n957), .B(new_n958), .C1(G311), .C2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT46), .B1(new_n838), .B2(G116), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n838), .A2(KEYINPUT46), .A3(G116), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n961), .B(new_n962), .C1(G317), .C2(new_n762), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n960), .B(new_n963), .C1(new_n203), .C2(new_n766), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n279), .B1(new_n746), .B2(new_n243), .C1(new_n333), .C2(new_n741), .ZN(new_n965));
  INV_X1    g0765(.A(new_n756), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n838), .A2(G58), .B1(new_n966), .B2(G77), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n773), .B2(new_n749), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n965), .B(new_n968), .C1(G137), .C2(new_n762), .ZN(new_n969));
  INV_X1    g0769(.A(G143), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n970), .B2(new_n769), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n766), .A2(new_n211), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n964), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT47), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n739), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n974), .B2(new_n973), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n793), .A2(new_n238), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n801), .B1(new_n223), .B2(new_n361), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n807), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT108), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n477), .A2(new_n677), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n484), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n729), .A2(new_n984), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n803), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n982), .A2(new_n983), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n646), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n657), .B1(new_n990), .B2(new_n677), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n567), .A2(new_n646), .A3(new_n676), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT105), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n690), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT42), .Z(new_n996));
  INV_X1    g0796(.A(new_n994), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n997), .A2(new_n582), .B1(new_n570), .B2(new_n572), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n677), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n996), .A2(new_n999), .B1(KEYINPUT43), .B2(new_n987), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n688), .A2(new_n997), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n694), .B(KEYINPUT41), .Z(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT106), .B1(new_n691), .B2(new_n994), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n691), .A2(new_n994), .A3(KEYINPUT106), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1010), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n691), .A2(new_n994), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT45), .Z(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n688), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n690), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n689), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1021), .B1(new_n687), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n683), .B(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n735), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1007), .B1(new_n1026), .B2(new_n735), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1006), .B1(new_n1027), .B2(new_n789), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT107), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(KEYINPUT107), .B(new_n1006), .C1(new_n1027), .C2(new_n789), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n989), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT110), .ZN(G387));
  NAND3_X1  g0833(.A1(new_n223), .A2(new_n279), .A3(new_n695), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(G107), .B2(new_n223), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n359), .A2(new_n243), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT50), .Z(new_n1037));
  AOI21_X1  g0837(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1037), .A2(new_n584), .A3(new_n456), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n793), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n235), .B2(G45), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1035), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n801), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n807), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n766), .A2(new_n361), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n773), .A2(new_n768), .B1(new_n749), .B2(new_n332), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n269), .A2(new_n757), .B1(new_n756), .B2(new_n202), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n741), .A2(new_n243), .B1(new_n746), .B2(new_n211), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n791), .B(new_n1049), .C1(new_n762), .C2(G150), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1045), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n742), .A2(G317), .B1(new_n825), .B2(G303), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n744), .B2(new_n749), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G322), .B2(new_n959), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT48), .Z(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n754), .B2(new_n766), .C1(new_n764), .C2(new_n757), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT49), .Z(new_n1057));
  OAI221_X1 g0857(.A(new_n791), .B1(new_n584), .B2(new_n756), .C1(new_n772), .C2(new_n767), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1051), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1044), .B1(new_n1059), .B2(new_n738), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n687), .A2(new_n803), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1060), .A2(new_n1061), .B1(new_n1024), .B2(new_n789), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1025), .A2(new_n694), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n735), .A2(new_n1024), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(G393));
  NAND2_X1  g0865(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1026), .A2(new_n694), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1018), .A2(new_n789), .A3(new_n1019), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1040), .A2(new_n242), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n801), .B1(new_n223), .B2(new_n202), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n807), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n749), .A2(new_n612), .B1(new_n757), .B2(new_n754), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n291), .B1(new_n746), .B2(new_n764), .C1(new_n203), .C2(new_n756), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G322), .C2(new_n762), .ZN(new_n1074));
  INV_X1    g0874(.A(G317), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n768), .A2(new_n1075), .B1(new_n741), .B2(new_n744), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1074), .B(new_n1077), .C1(new_n584), .C2(new_n766), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n766), .A2(new_n269), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n768), .A2(new_n333), .B1(new_n741), .B2(new_n773), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT51), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n791), .B1(G87), .B2(new_n966), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n762), .A2(G143), .B1(new_n359), .B2(new_n825), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G50), .A2(new_n750), .B1(new_n838), .B2(G68), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1078), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1071), .B1(new_n1086), .B2(new_n738), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n994), .B2(new_n803), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n1068), .A2(KEYINPUT111), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT111), .B1(new_n1068), .B2(new_n1088), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1067), .B1(new_n1089), .B2(new_n1090), .ZN(G390));
  NOR3_X1   g0891(.A1(new_n891), .A2(new_n892), .A3(new_n916), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT39), .B1(new_n908), .B2(new_n909), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1092), .A2(new_n1093), .B1(new_n937), .B2(new_n942), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n724), .A2(new_n820), .A3(new_n862), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n816), .B(new_n677), .C1(new_n728), .C2(new_n733), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n941), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n937), .B1(new_n862), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n910), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1094), .A2(new_n1095), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n864), .A2(G330), .A3(new_n820), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n859), .B2(new_n861), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n817), .A2(new_n941), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n937), .B1(new_n1103), .B2(new_n862), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n925), .B2(new_n935), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1098), .A2(new_n910), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1102), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n450), .A2(G330), .A3(new_n864), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n945), .A2(new_n643), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n862), .B1(new_n724), .B2(new_n820), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1103), .B1(new_n1110), .B2(new_n1102), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1097), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n859), .A2(new_n861), .A3(new_n1101), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n719), .A2(new_n722), .A3(G330), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n722), .B1(new_n719), .B2(G330), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n820), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n896), .A2(new_n897), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1112), .B(new_n1113), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1109), .B1(new_n1111), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1100), .A2(new_n1107), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1119), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(KEYINPUT112), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT112), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n694), .B(new_n1120), .C1(new_n1124), .C2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1100), .A2(new_n1107), .A3(new_n789), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n798), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n807), .B1(new_n433), .B2(new_n824), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n749), .A2(new_n203), .B1(new_n768), .B2(new_n754), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n779), .B(new_n1131), .C1(G68), .C2(new_n966), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n291), .B1(new_n741), .B2(new_n584), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G97), .B2(new_n825), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(new_n764), .C2(new_n772), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n766), .A2(new_n773), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n746), .A2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n291), .B(new_n1138), .C1(G132), .C2(new_n742), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n1140));
  NOR3_X1   g0940(.A1(new_n1140), .A2(new_n757), .A3(new_n333), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n762), .B2(G125), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n749), .A2(new_n827), .B1(new_n768), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G50), .B2(new_n966), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1140), .B1(new_n757), .B2(new_n333), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1139), .A2(new_n1142), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1135), .A2(new_n1079), .B1(new_n1136), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1130), .B1(new_n1148), .B2(new_n738), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1129), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1128), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT114), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1127), .A2(new_n1152), .ZN(G378));
  INV_X1    g0953(.A(new_n1109), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1120), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n346), .A2(new_n674), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n354), .B(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(KEYINPUT118), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT119), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n944), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1159), .A2(new_n1165), .A3(new_n1160), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(G330), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n899), .A2(new_n910), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT40), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n867), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(KEYINPUT40), .B2(new_n940), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1167), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n938), .A2(new_n943), .A3(new_n1162), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1164), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(G330), .B(new_n1166), .C1(new_n895), .C2(new_n911), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n938), .A2(new_n943), .A3(new_n1162), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1162), .B1(new_n938), .B2(new_n943), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1155), .A2(KEYINPUT57), .A3(new_n1174), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT120), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1178), .A2(new_n1174), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1182), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n1155), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1120), .A2(new_n1154), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1178), .A2(new_n1174), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1181), .A2(new_n1183), .A3(new_n694), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT121), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1182), .A2(new_n789), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1159), .A2(new_n798), .A3(new_n1160), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n807), .B1(G50), .B2(new_n824), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT117), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n792), .A2(G41), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G50), .B(new_n1194), .C1(new_n284), .C2(new_n302), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT115), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n749), .A2(new_n202), .B1(new_n768), .B2(new_n584), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G58), .B2(new_n966), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n741), .A2(new_n203), .B1(new_n746), .B2(new_n361), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G77), .B2(new_n838), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n762), .A2(G283), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n1194), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n972), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1196), .B1(KEYINPUT58), .B2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n284), .B(new_n302), .C1(new_n756), .C2(new_n773), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n762), .B2(G124), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n766), .A2(new_n333), .ZN(new_n1207));
  INV_X1    g1007(.A(G132), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n749), .A2(new_n1208), .B1(new_n746), .B2(new_n827), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT116), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n742), .A2(G128), .ZN(new_n1211));
  INV_X1    g1011(.A(G125), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n768), .C1(new_n757), .C2(new_n1137), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1207), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT59), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1206), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1214), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1204), .B1(KEYINPUT58), .B2(new_n1203), .C1(new_n1216), .C2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1193), .B1(new_n1219), .B2(new_n738), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1191), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1190), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1188), .A2(new_n1189), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1189), .B1(new_n1188), .B2(new_n1223), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(G375));
  AOI21_X1  g1026(.A(new_n1102), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1103), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1109), .B(new_n1118), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1230), .A2(new_n1119), .A3(new_n1007), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT122), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1208), .A2(new_n768), .B1(new_n749), .B2(new_n1137), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n742), .A2(G137), .B1(new_n825), .B2(G150), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n773), .B2(new_n757), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(G128), .C2(new_n762), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n792), .B1(new_n398), .B2(new_n756), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT124), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1236), .B(new_n1238), .C1(new_n243), .C2(new_n766), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n768), .A2(new_n764), .B1(new_n746), .B2(new_n203), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G116), .B2(new_n750), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT123), .Z(new_n1242));
  AOI21_X1  g1042(.A(new_n279), .B1(new_n742), .B2(G283), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n269), .B2(new_n756), .C1(new_n202), .C2(new_n757), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G303), .B2(new_n762), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1045), .A2(new_n1242), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n739), .B1(new_n1239), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n807), .B1(G68), .B2(new_n824), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n1117), .C2(new_n798), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1118), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n789), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1232), .A2(new_n1251), .ZN(G381));
  OR2_X1    g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(G381), .A2(G390), .A3(G384), .A4(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(G378), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  OR3_X1    g1056(.A1(G387), .A2(G375), .A3(new_n1256), .ZN(G407));
  NAND2_X1  g1057(.A1(new_n1188), .A2(new_n1223), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT121), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1188), .A2(new_n1189), .A3(new_n1223), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G378), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n675), .A2(G213), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(G213), .A3(new_n1264), .ZN(G409));
  NAND3_X1  g1065(.A1(new_n1188), .A2(G378), .A3(new_n1223), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1185), .A2(new_n1186), .A3(new_n1007), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1127), .B(new_n1152), .C1(new_n1222), .C2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1263), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1250), .B2(new_n1154), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT125), .B1(new_n1272), .B2(new_n1230), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1274), .B(new_n1229), .C1(new_n1119), .C2(new_n1271), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n694), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1230), .B2(KEYINPUT60), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1273), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1278), .A2(G384), .A3(new_n1251), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1278), .B2(new_n1251), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT126), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1279), .A2(new_n1280), .A3(KEYINPUT126), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1263), .A2(G2897), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1283), .ZN(new_n1285));
  OAI211_X1 g1085(.A(KEYINPUT126), .B(new_n1285), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT61), .B1(new_n1270), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1290), .B1(new_n1270), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT110), .B1(new_n1253), .B2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(G390), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1253), .A2(new_n1294), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(G390), .B2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(new_n1032), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1269), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1289), .A2(new_n1293), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1269), .A2(new_n1302), .A3(new_n1291), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1269), .B2(new_n1287), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1302), .B1(new_n1269), .B2(new_n1291), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1303), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1301), .B1(new_n1307), .B2(new_n1299), .ZN(G405));
  NAND2_X1  g1108(.A1(new_n1258), .A2(G378), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1291), .B1(new_n1261), .B2(new_n1310), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1292), .B(new_n1309), .C1(G375), .C2(G378), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1311), .A2(new_n1299), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1299), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(G402));
endmodule


