//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT75), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT24), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(G183gat), .A3(G190gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n209));
  XNOR2_X1  g008(.A(G183gat), .B(G190gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n209), .C1(new_n210), .C2(new_n206), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n212), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT25), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n207), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n217), .B1(new_n222), .B2(KEYINPUT24), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n213), .A2(new_n214), .ZN(new_n224));
  INV_X1    g023(.A(new_n208), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n212), .A2(G169gat), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT25), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n223), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  INV_X1    g032(.A(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT26), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n208), .A2(KEYINPUT66), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT27), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G183gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n243), .A3(new_n220), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT28), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT28), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n220), .ZN(new_n248));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n240), .A2(new_n245), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n216), .A2(new_n232), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(G226gat), .A3(G233gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT29), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n251), .A2(new_n254), .B1(G226gat), .B2(G233gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT73), .ZN(new_n256));
  INV_X1    g055(.A(G197gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(G204gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(G197gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n256), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(G197gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(G204gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT73), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(KEYINPUT74), .A2(KEYINPUT22), .ZN(new_n266));
  NOR2_X1   g065(.A1(KEYINPUT74), .A2(KEYINPUT22), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G211gat), .ZN(new_n270));
  INV_X1    g069(.A(G218gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(G211gat), .A2(G218gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n266), .B2(new_n267), .ZN(new_n276));
  INV_X1    g075(.A(new_n272), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n265), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n253), .A2(new_n255), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n251), .A2(new_n254), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n280), .B1(new_n285), .B2(new_n252), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n205), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n281), .B1(new_n253), .B2(new_n255), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n280), .A3(new_n252), .ZN(new_n289));
  INV_X1    g088(.A(new_n205), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(KEYINPUT30), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n288), .A2(new_n289), .A3(new_n293), .A4(new_n290), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G225gat), .A2(G233gat), .ZN(new_n297));
  INV_X1    g096(.A(G134gat), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT67), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G113gat), .B2(G120gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(G113gat), .A2(G120gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(G127gat), .A2(G134gat), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n303), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G127gat), .A2(G134gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n304), .B1(new_n311), .B2(new_n309), .ZN(new_n312));
  OR2_X1    g111(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(G113gat), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G113gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT69), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G113gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n319), .A3(G120gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n312), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT76), .B1(new_n310), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(new_n320), .ZN(new_n323));
  INV_X1    g122(.A(new_n312), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n326));
  INV_X1    g125(.A(G120gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n316), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n304), .A3(new_n306), .ZN(new_n329));
  INV_X1    g128(.A(new_n309), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT67), .B(G127gat), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n329), .B(new_n330), .C1(new_n298), .C2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n325), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G141gat), .B(G148gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n334), .B(new_n337), .C1(new_n338), .C2(KEYINPUT2), .ZN(new_n339));
  INV_X1    g138(.A(G141gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G148gat), .ZN(new_n341));
  INV_X1    g140(.A(G148gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G141gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n337), .A2(new_n334), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n334), .A2(KEYINPUT2), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n339), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n322), .A2(new_n333), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n325), .A2(new_n332), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT78), .B1(new_n353), .B2(new_n348), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n300), .A2(new_n302), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n309), .B1(new_n355), .B2(G134gat), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n329), .A2(new_n356), .B1(new_n323), .B2(new_n324), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n339), .A2(new_n347), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT4), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n353), .A2(new_n348), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n297), .B(new_n352), .C1(new_n361), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT5), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n322), .A2(new_n348), .A3(new_n333), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(new_n354), .A3(new_n360), .ZN(new_n368));
  INV_X1    g167(.A(new_n297), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n360), .A3(KEYINPUT4), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n362), .A2(new_n363), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n322), .A2(new_n333), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n349), .A2(new_n351), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n371), .A2(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n369), .A2(KEYINPUT5), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n365), .A2(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G1gat), .B(G29gat), .Z(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G57gat), .B(G85gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT6), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n372), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n352), .A3(new_n376), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n369), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT5), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n352), .A2(new_n297), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n353), .A2(KEYINPUT78), .A3(new_n348), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n359), .B1(new_n357), .B2(new_n358), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n362), .A2(new_n363), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n383), .B(new_n388), .C1(new_n390), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT80), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n377), .B2(new_n383), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n388), .B1(new_n390), .B2(new_n397), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(KEYINPUT81), .A3(new_n382), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n386), .A2(new_n401), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n296), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n251), .A2(new_n357), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n353), .A2(new_n216), .A3(new_n250), .A4(new_n232), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G227gat), .ZN(new_n412));
  INV_X1    g211(.A(G233gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n411), .B(new_n415), .C1(new_n412), .C2(new_n413), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT71), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n409), .A2(G227gat), .A3(G233gat), .A4(new_n410), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT32), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G71gat), .B(G99gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT70), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(G15gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G43gat), .ZN(new_n428));
  INV_X1    g227(.A(G15gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n426), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G43gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n422), .A2(new_n424), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT32), .B(new_n421), .C1(new_n433), .C2(new_n423), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n420), .B(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G22gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n351), .A2(new_n254), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n281), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n261), .A2(new_n264), .B1(new_n276), .B2(new_n277), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n266), .A2(new_n267), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n261), .B2(new_n264), .ZN(new_n445));
  INV_X1    g244(.A(new_n274), .ZN(new_n446));
  OAI22_X1  g245(.A1(new_n443), .A2(KEYINPUT84), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n265), .A2(KEYINPUT84), .A3(new_n278), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n254), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT85), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT85), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n451), .B(new_n254), .C1(new_n447), .C2(new_n448), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n350), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n442), .B1(new_n453), .B2(new_n348), .ZN(new_n454));
  INV_X1    g253(.A(G228gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n413), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT83), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT86), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n452), .A2(new_n350), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n279), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n443), .A2(KEYINPUT84), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n275), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n451), .B1(new_n464), .B2(new_n254), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n348), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n441), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n457), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n459), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT3), .B1(new_n280), .B2(new_n254), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n441), .B(new_n456), .C1(new_n471), .C2(new_n358), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n439), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  AOI211_X1 g273(.A(G22gat), .B(new_n474), .C1(new_n459), .C2(new_n469), .ZN(new_n475));
  XNOR2_X1  g274(.A(G78gat), .B(G106gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT31), .B(G50gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  NOR3_X1   g277(.A1(new_n473), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(KEYINPUT82), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n468), .B1(new_n467), .B2(new_n457), .ZN(new_n481));
  AOI211_X1 g280(.A(KEYINPUT86), .B(new_n458), .C1(new_n466), .C2(new_n441), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n472), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G22gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n470), .A2(new_n439), .A3(new_n472), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n408), .B(new_n438), .C1(new_n479), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n377), .A2(new_n383), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n407), .B1(new_n400), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT35), .B1(new_n292), .B2(new_n294), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n435), .A2(new_n436), .A3(new_n417), .A4(new_n418), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT88), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n435), .A2(new_n436), .B1(new_n417), .B2(new_n418), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n437), .A2(new_n419), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT88), .B1(new_n497), .B2(new_n492), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n490), .B(new_n491), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n480), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n473), .B2(new_n475), .ZN(new_n501));
  INV_X1    g300(.A(new_n478), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n485), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT36), .B1(new_n497), .B2(new_n492), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n438), .B2(KEYINPUT36), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n501), .A2(new_n503), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n407), .B(new_n291), .C1(new_n400), .C2(new_n489), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT37), .B1(new_n282), .B2(new_n286), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n288), .A2(new_n289), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n205), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT38), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT38), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n511), .A2(new_n516), .A3(new_n205), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n404), .A2(new_n382), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n387), .A2(new_n352), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n369), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT39), .B1(new_n368), .B2(new_n369), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT87), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(KEYINPUT39), .C1(new_n368), .C2(new_n369), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n297), .B1(new_n387), .B2(new_n352), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT39), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n382), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n520), .A2(KEYINPUT40), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n527), .A2(KEYINPUT40), .A3(new_n530), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n531), .A2(new_n532), .A3(new_n295), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n519), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n508), .B1(new_n509), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n403), .B(new_n405), .C1(new_n384), .C2(new_n385), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n400), .A2(KEYINPUT80), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n407), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n295), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(new_n501), .A3(new_n503), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n506), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n538), .ZN(new_n543));
  NAND2_X1  g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  INV_X1    g343(.A(G71gat), .ZN(new_n545));
  INV_X1    g344(.A(G78gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT9), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n544), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G57gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G64gat), .ZN(new_n552));
  INV_X1    g351(.A(G64gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(G57gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n547), .A2(new_n544), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n544), .A2(new_n549), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G127gat), .B(G155gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT20), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G8gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572));
  INV_X1    g371(.A(G1gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT16), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n572), .A2(G1gat), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT92), .B(new_n571), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n571), .A2(KEYINPUT92), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n571), .A2(KEYINPUT92), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n579), .A2(new_n575), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n560), .B2(new_n559), .ZN(new_n584));
  XOR2_X1   g383(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n586), .A3(new_n569), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT91), .B(KEYINPUT17), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G36gat), .ZN(new_n593));
  AND2_X1   g392(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G29gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G43gat), .B(G50gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT15), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G50gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(G43gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n431), .A2(G50gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT89), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT15), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n431), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n610), .A2(new_n599), .A3(KEYINPUT90), .A4(new_n601), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n602), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n596), .A2(new_n598), .B1(new_n600), .B2(KEYINPUT15), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT90), .B1(new_n613), .B2(new_n610), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n592), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n610), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT90), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n618), .A2(KEYINPUT17), .A3(new_n602), .A4(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT7), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT7), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(G85gat), .A3(G92gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  INV_X1    g425(.A(G92gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(KEYINPUT8), .A2(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G99gat), .B(G106gat), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n624), .B2(new_n628), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n615), .B(new_n619), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n602), .A3(new_n611), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n631), .A2(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT97), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n634), .A2(new_n635), .B1(KEYINPUT41), .B2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G190gat), .B(G218gat), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n633), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n633), .B2(new_n639), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n638), .A2(KEYINPUT41), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OR3_X1    g446(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n642), .B2(new_n643), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n590), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G230gat), .A2(G233gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n559), .B1(new_n631), .B2(new_n632), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n624), .A2(new_n628), .ZN(new_n660));
  INV_X1    g459(.A(new_n629), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n662), .A2(new_n550), .A3(new_n558), .A4(new_n630), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n659), .A2(KEYINPUT98), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n559), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n635), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT10), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n663), .A2(new_n669), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n658), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n664), .A2(new_n667), .A3(new_n658), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT99), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n664), .A2(new_n667), .A3(new_n676), .A4(new_n658), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n656), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT10), .B1(new_n664), .B2(new_n667), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n657), .B1(new_n680), .B2(new_n671), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n681), .A2(new_n655), .A3(new_n677), .A4(new_n675), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n652), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n634), .A2(new_n578), .A3(new_n582), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n583), .A2(new_n618), .A3(new_n602), .A4(new_n611), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(G229gat), .A2(G233gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT93), .Z(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n615), .A2(new_n583), .A3(new_n619), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n693), .A2(KEYINPUT18), .A3(new_n685), .A4(new_n689), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n685), .A3(new_n689), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT18), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(G113gat), .B(G141gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G197gat), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT11), .B(G169gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT12), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n695), .B(new_n698), .C1(KEYINPUT94), .C2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n692), .A2(new_n694), .A3(KEYINPUT94), .ZN(new_n707));
  INV_X1    g506(.A(new_n698), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n694), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n707), .B(new_n704), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n684), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n542), .A2(new_n543), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g513(.A(new_n534), .B1(new_n479), .B2(new_n486), .ZN(new_n715));
  INV_X1    g514(.A(new_n508), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n715), .A2(new_n540), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n504), .B1(new_n487), .B2(KEYINPUT35), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n296), .B(new_n712), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT16), .B(G8gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT101), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n719), .A2(KEYINPUT100), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT100), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n542), .A2(new_n725), .A3(new_n296), .A4(new_n712), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n722), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n726), .A3(G8gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  OAI221_X1 g530(.A(new_n723), .B1(KEYINPUT42), .B2(new_n727), .C1(new_n730), .C2(new_n731), .ZN(G1325gat));
  NAND2_X1  g531(.A1(new_n542), .A2(new_n712), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n508), .B(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G15gat), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n496), .ZN(new_n738));
  INV_X1    g537(.A(new_n498), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n429), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n737), .B1(new_n733), .B2(new_n741), .ZN(G1326gat));
  INV_X1    g541(.A(new_n509), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n542), .A2(new_n743), .A3(new_n712), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT104), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT43), .B(G22gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1327gat));
  AOI21_X1  g546(.A(new_n650), .B1(new_n506), .B2(new_n541), .ZN(new_n748));
  INV_X1    g547(.A(new_n590), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n679), .A2(new_n682), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n749), .A2(new_n711), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n748), .A2(new_n597), .A3(new_n543), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT45), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n488), .A2(new_n505), .B1(new_n535), .B2(new_n540), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(new_n650), .ZN(new_n756));
  OAI211_X1 g555(.A(KEYINPUT44), .B(new_n651), .C1(new_n717), .C2(new_n718), .ZN(new_n757));
  AND4_X1   g556(.A1(new_n543), .A2(new_n756), .A3(new_n757), .A4(new_n751), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n597), .B2(new_n758), .ZN(G1328gat));
  AOI211_X1 g558(.A(G36gat), .B(new_n295), .C1(KEYINPUT105), .C2(KEYINPUT46), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n748), .A2(new_n751), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AND4_X1   g562(.A1(new_n296), .A2(new_n756), .A3(new_n757), .A4(new_n751), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n593), .B2(new_n764), .ZN(G1329gat));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n751), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n740), .A2(new_n431), .ZN(new_n767));
  AND4_X1   g566(.A1(new_n508), .A2(new_n756), .A3(new_n757), .A4(new_n751), .ZN(new_n768));
  OAI221_X1 g567(.A(KEYINPUT47), .B1(new_n766), .B2(new_n767), .C1(new_n768), .C2(new_n431), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n766), .A2(new_n767), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n756), .A2(new_n735), .A3(new_n757), .A4(new_n751), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(G43gat), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n772), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g572(.A1(new_n748), .A2(new_n743), .A3(new_n751), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n774), .A2(new_n603), .B1(new_n775), .B2(KEYINPUT48), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n509), .A2(new_n603), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n756), .A2(new_n757), .A3(new_n751), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n775), .A2(KEYINPUT48), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1331gat));
  NAND3_X1  g580(.A1(new_n652), .A2(new_n711), .A3(new_n750), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n755), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n543), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G57gat), .ZN(G1332gat));
  OAI21_X1  g584(.A(KEYINPUT107), .B1(new_n755), .B2(new_n782), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n787));
  INV_X1    g586(.A(new_n782), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n787), .B(new_n788), .C1(new_n717), .C2(new_n718), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n790), .A2(new_n295), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT49), .B(G64gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n786), .A2(new_n296), .A3(new_n789), .A4(new_n793), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n792), .B1(new_n791), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(G1333gat));
  OAI21_X1  g596(.A(G71gat), .B1(new_n790), .B2(new_n736), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n545), .A3(new_n740), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g599(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n801), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1334gat));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n509), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(new_n546), .ZN(G1335gat));
  NAND2_X1  g606(.A1(new_n590), .A2(new_n711), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT110), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n750), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n756), .A2(new_n543), .A3(new_n757), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G85gat), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT51), .B1(new_n748), .B2(new_n809), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n651), .B(new_n809), .C1(new_n717), .C2(new_n718), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n543), .A2(new_n626), .A3(new_n750), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n812), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n812), .B(KEYINPUT111), .C1(new_n817), .C2(new_n818), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1336gat));
  NAND4_X1  g622(.A1(new_n756), .A2(new_n296), .A3(new_n757), .A4(new_n810), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G92gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT112), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n295), .A2(new_n683), .A3(G92gat), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n813), .B2(new_n816), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n825), .B(new_n828), .C1(KEYINPUT112), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1337gat));
  NAND4_X1  g632(.A1(new_n756), .A2(new_n735), .A3(new_n757), .A4(new_n810), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G99gat), .ZN(new_n835));
  AOI211_X1 g634(.A(G99gat), .B(new_n683), .C1(new_n738), .C2(new_n739), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT113), .Z(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n817), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n835), .B(new_n840), .C1(new_n817), .C2(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(G1338gat));
  XNOR2_X1  g641(.A(new_n814), .B(new_n815), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n509), .A2(G106gat), .A3(new_n683), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n756), .A2(new_n743), .A3(new_n757), .A4(new_n810), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G106gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n845), .B(KEYINPUT116), .Z(new_n851));
  AOI22_X1  g650(.A1(new_n851), .A2(new_n843), .B1(G106gat), .B2(new_n848), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n852), .B2(new_n847), .ZN(G1339gat));
  NAND3_X1  g652(.A1(new_n652), .A2(new_n711), .A3(new_n683), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n687), .A2(new_n691), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n689), .B1(new_n693), .B2(new_n685), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n704), .B1(new_n696), .B2(new_n697), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n857), .A2(new_n702), .B1(new_n695), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n648), .A3(new_n649), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n670), .A2(new_n658), .A3(new_n672), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n862), .A2(KEYINPUT54), .A3(new_n681), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n656), .B1(new_n681), .B2(KEYINPUT54), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n655), .B1(new_n673), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n862), .A2(KEYINPUT54), .A3(new_n681), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(KEYINPUT55), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n682), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n860), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n702), .B1(new_n855), .B2(new_n856), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n698), .A2(new_n705), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n709), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT117), .B1(new_n683), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n876), .A3(new_n750), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n875), .B(new_n877), .C1(new_n711), .C2(new_n870), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n871), .B1(new_n878), .B2(new_n650), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n854), .B1(new_n879), .B2(new_n749), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT118), .B(new_n854), .C1(new_n879), .C2(new_n749), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n543), .A2(new_n295), .A3(new_n740), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n882), .A2(new_n509), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT119), .ZN(new_n886));
  INV_X1    g685(.A(new_n711), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n509), .A2(new_n438), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n882), .A2(new_n543), .A3(new_n889), .A4(new_n883), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT120), .B1(new_n890), .B2(new_n296), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n890), .A2(KEYINPUT120), .A3(new_n296), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n887), .A2(new_n317), .A3(new_n319), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n888), .A2(new_n316), .B1(new_n894), .B2(new_n895), .ZN(G1340gat));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n327), .B1(new_n886), .B2(new_n750), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n750), .A2(new_n313), .A3(new_n314), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT121), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n890), .A2(KEYINPUT120), .A3(new_n296), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n891), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n897), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n885), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n885), .A2(new_n905), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n750), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G120gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n900), .B1(new_n892), .B2(new_n893), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n904), .A2(new_n911), .ZN(G1341gat));
  NOR3_X1   g711(.A1(new_n890), .A2(new_n296), .A3(new_n590), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT123), .Z(new_n914));
  NOR2_X1   g713(.A1(new_n590), .A2(new_n331), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n914), .A2(new_n331), .B1(new_n886), .B2(new_n915), .ZN(G1342gat));
  NOR4_X1   g715(.A1(new_n890), .A2(G134gat), .A3(new_n296), .A4(new_n650), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT56), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n886), .A2(new_n651), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n298), .ZN(G1343gat));
  NAND3_X1  g719(.A1(new_n716), .A2(new_n543), .A3(new_n295), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n882), .A2(new_n743), .A3(new_n883), .ZN(new_n922));
  XOR2_X1   g721(.A(KEYINPUT124), .B(KEYINPUT57), .Z(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n711), .A2(new_n870), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n859), .A2(new_n750), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n650), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n871), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n749), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n854), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(new_n509), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT57), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n921), .B1(new_n924), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n340), .B1(new_n935), .B2(new_n887), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n882), .A2(new_n883), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(new_n538), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n735), .A2(new_n509), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n711), .A2(G141gat), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n938), .A2(new_n295), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT58), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT58), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n711), .B(new_n921), .C1(new_n924), .C2(new_n934), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n941), .B(new_n944), .C1(new_n945), .C2(new_n340), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n946), .ZN(G1344gat));
  NAND2_X1  g746(.A1(new_n938), .A2(new_n939), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n296), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n342), .A3(new_n750), .ZN(new_n950));
  AOI211_X1 g749(.A(KEYINPUT59), .B(new_n342), .C1(new_n935), .C2(new_n750), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n952));
  INV_X1    g751(.A(new_n923), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n882), .A2(new_n743), .A3(new_n883), .A4(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT57), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n955), .B1(new_n932), .B2(new_n509), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n921), .A2(new_n683), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n952), .B1(new_n959), .B2(G148gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n950), .B1(new_n951), .B2(new_n960), .ZN(G1345gat));
  INV_X1    g760(.A(new_n935), .ZN(new_n962));
  OAI21_X1  g761(.A(G155gat), .B1(new_n962), .B2(new_n590), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n949), .A2(new_n335), .A3(new_n749), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1346gat));
  OAI21_X1  g764(.A(G162gat), .B1(new_n962), .B2(new_n650), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n651), .A2(new_n336), .A3(new_n295), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n948), .B2(new_n967), .ZN(G1347gat));
  NOR2_X1   g767(.A1(new_n543), .A2(new_n295), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n969), .A2(new_n740), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n882), .A2(new_n509), .A3(new_n883), .A4(new_n970), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n971), .A2(new_n233), .A3(new_n711), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n937), .A2(new_n543), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n889), .A2(new_n296), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(new_n887), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n972), .B1(new_n977), .B2(new_n233), .ZN(G1348gat));
  NOR3_X1   g777(.A1(new_n971), .A2(new_n229), .A3(new_n683), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(new_n750), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(new_n234), .ZN(G1349gat));
  OAI21_X1  g780(.A(G183gat), .B1(new_n971), .B2(new_n590), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n749), .A2(new_n246), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n982), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g784(.A1(new_n976), .A2(new_n220), .A3(new_n651), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n971), .A2(new_n650), .ZN(new_n987));
  XNOR2_X1  g786(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(G190gat), .A3(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n988), .B1(new_n987), .B2(G190gat), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n986), .B1(new_n990), .B2(new_n991), .ZN(G1351gat));
  NAND2_X1  g791(.A1(new_n736), .A2(new_n969), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n993), .B1(new_n954), .B2(new_n956), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n995), .A2(new_n257), .A3(new_n711), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n939), .A2(new_n296), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(new_n973), .ZN(new_n999));
  INV_X1    g798(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(new_n887), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n996), .B1(new_n1001), .B2(new_n257), .ZN(G1352gat));
  NAND2_X1  g801(.A1(new_n750), .A2(new_n259), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1004), .B1(KEYINPUT127), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g805(.A(G204gat), .B1(new_n995), .B2(new_n683), .ZN(new_n1007));
  XOR2_X1   g806(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1008));
  OAI21_X1  g807(.A(new_n1008), .B1(new_n999), .B2(new_n1003), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(G1353gat));
  NAND3_X1  g809(.A1(new_n1000), .A2(new_n270), .A3(new_n749), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n749), .ZN(new_n1012));
  AND3_X1   g811(.A1(new_n1012), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1013));
  AOI21_X1  g812(.A(KEYINPUT63), .B1(new_n1012), .B2(G211gat), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(G1354gat));
  OAI21_X1  g814(.A(G218gat), .B1(new_n995), .B2(new_n650), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n651), .A2(new_n271), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1016), .B1(new_n999), .B2(new_n1017), .ZN(G1355gat));
endmodule


