//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT72), .B(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT74), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT16), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n192), .A3(G125), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n191), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n191), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n190), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n203));
  XNOR2_X1  g017(.A(G125), .B(G140), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(KEYINPUT16), .ZN(new_n205));
  OAI211_X1 g019(.A(G146), .B(new_n200), .C1(new_n205), .C2(new_n191), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n206), .A3(KEYINPUT75), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT75), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n208), .B(new_n190), .C1(new_n199), .C2(new_n201), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT68), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n215), .A3(G128), .ZN(new_n216));
  AOI21_X1  g030(.A(G128), .B1(new_n213), .B2(new_n215), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n211), .B(new_n216), .C1(new_n217), .C2(KEYINPUT23), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT73), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n212), .B2(G128), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n210), .A2(KEYINPUT73), .A3(G119), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n216), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT24), .B(G110), .Z(new_n223));
  AOI22_X1  g037(.A1(G110), .A2(new_n218), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n207), .A2(new_n209), .A3(new_n224), .ZN(new_n225));
  OAI22_X1  g039(.A1(new_n218), .A2(G110), .B1(new_n222), .B2(new_n223), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n193), .A2(new_n195), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n204), .A2(KEYINPUT76), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT65), .A2(G146), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT65), .A2(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n206), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G953), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(G221), .A3(G234), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n237), .B(KEYINPUT77), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT22), .B(G137), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n225), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n225), .B2(new_n235), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT25), .B1(new_n243), .B2(new_n188), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n225), .A2(new_n235), .ZN(new_n245));
  INV_X1    g059(.A(new_n240), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n225), .A2(new_n235), .A3(new_n240), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n189), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT78), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n188), .A3(new_n248), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n249), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT78), .A3(new_n189), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n189), .A2(G902), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n243), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(G472), .A2(G902), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT2), .B(G113), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n212), .B2(G116), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT68), .B(G119), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G116), .ZN(new_n268));
  AND4_X1   g082(.A1(KEYINPUT69), .A2(new_n213), .A3(new_n215), .A4(G116), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n264), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n213), .A2(new_n215), .A3(G116), .ZN(new_n271));
  INV_X1    g085(.A(new_n266), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n267), .A2(KEYINPUT69), .A3(G116), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n263), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n190), .B2(G143), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n233), .B2(G143), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n190), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT65), .A2(G146), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(KEYINPUT66), .A3(G143), .A4(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n278), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT11), .ZN(new_n288));
  INV_X1    g102(.A(G134), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(G137), .ZN(new_n290));
  INV_X1    g104(.A(G137), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT11), .A3(G134), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(G137), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G131), .ZN(new_n295));
  INV_X1    g109(.A(G131), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n290), .A2(new_n292), .A3(new_n296), .A4(new_n293), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(KEYINPUT67), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n294), .A2(new_n299), .A3(G131), .ZN(new_n300));
  INV_X1    g114(.A(G143), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n231), .B2(new_n232), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT64), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n301), .B2(G146), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n190), .A2(KEYINPUT64), .A3(G143), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(KEYINPUT0), .A2(G128), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n278), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n287), .A2(new_n298), .A3(new_n300), .A4(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n293), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n289), .A2(G137), .ZN(new_n313));
  OAI21_X1  g127(.A(G131), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n314), .A2(new_n297), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n283), .A2(G143), .A3(new_n284), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT1), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n304), .A2(new_n305), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n317), .A2(G128), .B1(new_n318), .B2(new_n302), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n280), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n321), .B1(new_n323), .B2(new_n285), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n315), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n311), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n311), .B2(new_n325), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n276), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT26), .B(G101), .ZN(new_n330));
  NOR2_X1   g144(.A1(G237), .A2(G953), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G210), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n268), .A2(new_n269), .A3(new_n264), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n263), .B1(new_n273), .B2(new_n274), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n311), .A2(new_n325), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n329), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT31), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT31), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n329), .A2(new_n343), .A3(new_n336), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n311), .A2(new_n325), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n276), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n348), .B2(new_n340), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n340), .A2(new_n346), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT71), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT71), .B1(new_n340), .B2(new_n346), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n336), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n262), .B1(new_n345), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT32), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT32), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n358), .B(new_n262), .C1(new_n345), .C2(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n352), .A2(KEYINPUT29), .A3(new_n336), .A4(new_n354), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n311), .A2(new_n325), .A3(new_n339), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n339), .B1(new_n311), .B2(new_n325), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT28), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n350), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n335), .B(new_n353), .C1(new_n365), .C2(KEYINPUT71), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT29), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n329), .A2(new_n340), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(new_n336), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n188), .B(new_n361), .C1(new_n366), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G472), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n261), .B1(new_n360), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G214), .B1(G237), .B2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G210), .B1(G237), .B2(G902), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G101), .ZN(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n378), .B2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G104), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(G107), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n377), .B1(new_n384), .B2(KEYINPUT79), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n379), .A2(new_n382), .A3(new_n386), .A4(new_n383), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n379), .A2(new_n382), .A3(new_n377), .A4(new_n383), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT4), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n393), .A3(new_n387), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n276), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n378), .A2(G107), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n381), .A2(G104), .ZN(new_n397));
  OAI21_X1  g211(.A(G101), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n389), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n273), .B2(new_n274), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n213), .A2(new_n215), .A3(new_n401), .A4(G116), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G113), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n270), .B(new_n400), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n395), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G110), .B(G122), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n405), .A3(new_n407), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT83), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n320), .B1(new_n281), .B2(new_n286), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT1), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n233), .B2(G143), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n306), .B1(new_n416), .B2(new_n210), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n417), .A3(new_n194), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n277), .B1(new_n323), .B2(new_n285), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n308), .B1(new_n318), .B2(new_n302), .ZN(new_n420));
  OAI21_X1  g234(.A(G125), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G224), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(G953), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n422), .B(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n406), .B(new_n408), .C1(KEYINPUT83), .C2(new_n411), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n413), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G902), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n418), .A2(new_n421), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT86), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n418), .A2(new_n421), .A3(new_n433), .A4(new_n430), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT7), .B1(new_n423), .B2(G953), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n422), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n410), .A2(new_n432), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n407), .B(KEYINPUT8), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT5), .B1(new_n268), .B2(new_n269), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n403), .A2(new_n441), .A3(G113), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n404), .A2(KEYINPUT84), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n338), .A2(new_n399), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT85), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n270), .B1(new_n402), .B2(new_n404), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n446), .A2(new_n447), .B1(new_n399), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT85), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n439), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n428), .B1(new_n437), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n376), .B1(new_n427), .B2(new_n452), .ZN(new_n453));
  AND4_X1   g267(.A1(new_n410), .A2(new_n432), .A3(new_n434), .A4(new_n436), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n449), .A2(new_n450), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n438), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n413), .A2(new_n425), .A3(new_n426), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n375), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n374), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT9), .B(G234), .ZN(new_n461));
  OAI21_X1  g275(.A(G221), .B1(new_n461), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n188), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n298), .A2(new_n300), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT10), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT1), .B1(new_n301), .B2(G146), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G128), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n323), .A2(new_n285), .A3(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n465), .B(new_n400), .C1(new_n468), .C2(new_n324), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n399), .B1(new_n414), .B2(new_n417), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n465), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n419), .A2(new_n420), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n392), .A2(new_n472), .A3(new_n394), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n464), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n400), .B1(new_n319), .B2(new_n324), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT10), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n384), .A2(KEYINPUT79), .ZN(new_n478));
  AND4_X1   g292(.A1(new_n393), .A2(new_n478), .A3(G101), .A4(new_n387), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n390), .B1(new_n385), .B2(new_n387), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n477), .A2(new_n469), .B1(new_n481), .B2(new_n472), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n298), .A2(new_n483), .A3(new_n300), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n298), .B2(new_n300), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT81), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n471), .A2(new_n486), .A3(KEYINPUT81), .A4(new_n473), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n475), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G110), .B(G140), .ZN(new_n491));
  INV_X1    g305(.A(G227), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(G953), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n491), .B(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n471), .A2(new_n473), .A3(new_n486), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT81), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n488), .ZN(new_n499));
  INV_X1    g313(.A(new_n494), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT82), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n400), .B1(new_n468), .B2(new_n324), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n414), .A2(new_n417), .A3(new_n399), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n464), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT12), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT12), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n507), .B(new_n464), .C1(new_n502), .C2(new_n503), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n501), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n319), .A2(new_n324), .A3(new_n400), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n323), .A2(new_n285), .A3(new_n467), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n399), .B1(new_n414), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n505), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n507), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n504), .A2(KEYINPUT12), .A3(new_n505), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(KEYINPUT82), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n499), .A2(new_n500), .A3(new_n509), .A4(new_n516), .ZN(new_n517));
  AOI211_X1 g331(.A(G469), .B(new_n463), .C1(new_n495), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n499), .A2(new_n475), .A3(new_n500), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n498), .A2(new_n488), .B1(new_n515), .B2(new_n514), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(G469), .C1(new_n500), .C2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G469), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(new_n428), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n460), .B(new_n462), .C1(new_n518), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G113), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n378), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT19), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n229), .A2(new_n230), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n227), .A2(KEYINPUT19), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n233), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G237), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n236), .A3(G214), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n301), .A2(KEYINPUT87), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G143), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n331), .A2(G214), .B1(new_n537), .B2(G143), .ZN(new_n540));
  OAI21_X1  g354(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n538), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT87), .B(G143), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n542), .B(new_n296), .C1(new_n535), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n533), .A2(new_n545), .A3(new_n206), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n227), .A2(G146), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n234), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n542), .B1(new_n543), .B2(new_n535), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(KEYINPUT18), .A3(G131), .ZN(new_n550));
  NAND2_X1  g364(.A1(KEYINPUT18), .A2(G131), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n542), .B(new_n551), .C1(new_n535), .C2(new_n543), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n529), .B1(new_n546), .B2(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n207), .A2(new_n209), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n541), .A2(new_n557), .A3(new_n544), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n549), .A2(KEYINPUT17), .A3(G131), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n555), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n554), .B1(new_n561), .B2(new_n529), .ZN(new_n562));
  NOR2_X1   g376(.A1(G475), .A2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT20), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT20), .ZN(new_n566));
  INV_X1    g380(.A(new_n529), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n567), .B(new_n555), .C1(new_n556), .C2(new_n560), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n566), .B(new_n563), .C1(new_n568), .C2(new_n554), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n561), .A2(new_n529), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n428), .B1(new_n571), .B2(new_n568), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT88), .B(G475), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n570), .A2(KEYINPUT89), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT89), .B1(new_n570), .B2(new_n575), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n461), .A2(new_n187), .A3(G953), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(G128), .B(G143), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(new_n289), .ZN(new_n581));
  INV_X1    g395(.A(G122), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G116), .ZN(new_n583));
  INV_X1    g397(.A(G116), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G122), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n585), .A3(new_n381), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n583), .B1(new_n585), .B2(KEYINPUT14), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT14), .B1(new_n582), .B2(G116), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT91), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n585), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n581), .B(new_n586), .C1(new_n381), .C2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT92), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n580), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n301), .A2(G128), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n596), .B(G134), .C1(new_n597), .C2(new_n595), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n580), .A2(new_n289), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n583), .A2(new_n585), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G107), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n586), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n593), .A2(new_n594), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n594), .B1(new_n593), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n579), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n593), .A2(new_n603), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT92), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n593), .A2(new_n603), .A3(new_n594), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n578), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n606), .A2(new_n610), .A3(new_n188), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(G478), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(KEYINPUT15), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n606), .A2(new_n610), .A3(KEYINPUT93), .A4(new_n188), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n611), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g432(.A1(G234), .A2(G237), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n619), .A2(G952), .A3(new_n236), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT21), .B(G898), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT94), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n463), .A2(G953), .A3(new_n619), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n617), .A2(new_n618), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n576), .A2(new_n577), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n372), .A2(new_n527), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  NOR3_X1   g443(.A1(new_n427), .A2(new_n452), .A3(new_n376), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n375), .B1(new_n457), .B2(new_n458), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n373), .B(new_n625), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n606), .A2(new_n610), .A3(KEYINPUT33), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT33), .B1(new_n606), .B2(new_n610), .ZN(new_n635));
  OAI211_X1 g449(.A(G478), .B(new_n188), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n556), .A2(new_n560), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n529), .A3(new_n553), .ZN(new_n640));
  INV_X1    g454(.A(new_n554), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n566), .B1(new_n642), .B2(new_n563), .ZN(new_n643));
  AOI211_X1 g457(.A(KEYINPUT20), .B(new_n564), .C1(new_n640), .C2(new_n641), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n639), .A2(new_n553), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n567), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n646), .B2(new_n640), .ZN(new_n647));
  OAI22_X1  g461(.A1(new_n643), .A2(new_n644), .B1(new_n647), .B2(new_n573), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT89), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n570), .A2(new_n575), .A3(KEYINPUT89), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n638), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(KEYINPUT95), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n636), .A2(new_n637), .ZN(new_n654));
  OAI211_X1 g468(.A(KEYINPUT95), .B(new_n654), .C1(new_n576), .C2(new_n577), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n633), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n462), .ZN(new_n658));
  OAI22_X1  g472(.A1(new_n487), .A2(new_n489), .B1(new_n508), .B2(new_n506), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n494), .B1(new_n498), .B2(new_n488), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n659), .A2(new_n494), .B1(new_n660), .B2(new_n475), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n523), .B1(new_n661), .B2(G469), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n500), .B1(new_n487), .B2(new_n489), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n509), .A2(new_n516), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n474), .B1(new_n498), .B2(new_n488), .ZN(new_n665));
  OAI22_X1  g479(.A1(new_n663), .A2(new_n664), .B1(new_n665), .B2(new_n500), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n522), .A3(new_n188), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n658), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n261), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n188), .B1(new_n345), .B2(new_n355), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n353), .B1(new_n365), .B2(KEYINPUT71), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n342), .B(new_n344), .C1(new_n671), .C2(new_n336), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n670), .A2(G472), .B1(new_n672), .B2(new_n262), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n657), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT34), .B(G104), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G6));
  OR2_X1    g491(.A1(new_n570), .A2(KEYINPUT96), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n617), .A2(new_n618), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n643), .A2(KEYINPUT96), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n678), .A2(new_n575), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n674), .A2(new_n632), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT35), .B(G107), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  NOR2_X1   g498(.A1(new_n246), .A2(KEYINPUT36), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT97), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n245), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n259), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n253), .A2(new_n258), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n670), .A2(G472), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n689), .A2(new_n356), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n527), .A2(new_n691), .A3(new_n627), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  AOI22_X1  g508(.A1(new_n357), .A2(new_n359), .B1(G472), .B2(new_n370), .ZN(new_n695));
  INV_X1    g509(.A(new_n689), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n695), .A2(new_n526), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n678), .A2(new_n680), .ZN(new_n698));
  INV_X1    g512(.A(new_n679), .ZN(new_n699));
  INV_X1    g513(.A(G900), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n623), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(new_n620), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n575), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n698), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT98), .B(G128), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G30));
  NOR2_X1   g521(.A1(new_n630), .A2(new_n631), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n576), .A2(new_n577), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n699), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n710), .A2(new_n373), .A3(new_n696), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n702), .B(KEYINPUT39), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n668), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n715), .B(KEYINPUT104), .Z(new_n716));
  AOI21_X1  g530(.A(new_n713), .B1(new_n716), .B2(KEYINPUT40), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n335), .B1(new_n362), .B2(new_n363), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n341), .A2(KEYINPUT100), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n428), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT100), .B1(new_n341), .B2(new_n718), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT101), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(KEYINPUT101), .B(G472), .C1(new_n720), .C2(new_n721), .ZN(new_n725));
  INV_X1    g539(.A(new_n359), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n358), .B1(new_n672), .B2(new_n262), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n724), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n360), .A2(KEYINPUT102), .A3(new_n724), .A4(new_n725), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT103), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n717), .B(new_n733), .C1(KEYINPUT40), .C2(new_n716), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT105), .B(G143), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G45));
  OAI211_X1 g550(.A(new_n654), .B(new_n702), .C1(new_n576), .C2(new_n577), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n697), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  AND2_X1   g554(.A1(new_n509), .A2(new_n516), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n660), .A2(new_n741), .B1(new_n490), .B2(new_n494), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n742), .B2(new_n463), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n462), .A3(new_n667), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n371), .B1(new_n726), .B2(new_n727), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n743), .A2(KEYINPUT106), .A3(new_n462), .A4(new_n667), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n669), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n657), .ZN(new_n750));
  XOR2_X1   g564(.A(KEYINPUT41), .B(G113), .Z(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G15));
  AOI21_X1  g566(.A(new_n522), .B1(new_n666), .B2(new_n188), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n518), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT106), .B1(new_n754), .B2(new_n462), .ZN(new_n755));
  INV_X1    g569(.A(new_n748), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n681), .A2(new_n632), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(KEYINPUT107), .A3(new_n372), .A4(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n372), .A2(new_n758), .A3(new_n746), .A4(new_n748), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT108), .B(G116), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G18));
  NAND3_X1  g579(.A1(new_n746), .A2(new_n460), .A3(new_n748), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n747), .A2(new_n627), .A3(new_n689), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT109), .B(G119), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G21));
  AOI21_X1  g584(.A(KEYINPUT78), .B1(new_n257), .B2(new_n189), .ZN(new_n771));
  INV_X1    g585(.A(new_n189), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n252), .B(new_n772), .C1(new_n256), .C2(new_n249), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT111), .A3(new_n260), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n261), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n670), .A2(new_n779), .A3(G472), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n690), .A2(KEYINPUT110), .B1(new_n672), .B2(new_n262), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n746), .A2(new_n633), .A3(new_n712), .A4(new_n748), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n582), .ZN(G24));
  NAND4_X1  g599(.A1(new_n781), .A2(new_n738), .A3(new_n689), .A4(new_n780), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n766), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT112), .B(G125), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G27));
  NAND3_X1  g603(.A1(new_n453), .A2(new_n373), .A3(new_n459), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n658), .B(new_n790), .C1(new_n667), .C2(new_n662), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n778), .A2(new_n791), .A3(new_n747), .A4(new_n738), .ZN(new_n792));
  INV_X1    g606(.A(new_n790), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n793), .B(new_n462), .C1(new_n518), .C2(new_n525), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n695), .A3(new_n261), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n792), .A2(KEYINPUT42), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G131), .ZN(G33));
  NAND3_X1  g612(.A1(new_n372), .A2(new_n791), .A3(new_n704), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G134), .ZN(G36));
  NAND2_X1  g614(.A1(new_n711), .A2(new_n654), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT43), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT43), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n711), .A2(new_n803), .A3(new_n654), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n673), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n689), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n790), .B1(new_n807), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n661), .A2(KEYINPUT45), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n519), .B1(new_n500), .B2(new_n520), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(new_n814), .A3(G469), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n524), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT46), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n667), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n816), .A2(new_n817), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n462), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n809), .A2(new_n810), .A3(new_n714), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(KEYINPUT113), .B(G137), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(G39));
  INV_X1    g639(.A(KEYINPUT47), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(KEYINPUT47), .B(new_n462), .C1(new_n819), .C2(new_n820), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n747), .A2(new_n669), .A3(new_n737), .A4(new_n790), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G140), .ZN(G42));
  INV_X1    g646(.A(new_n778), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n710), .A2(new_n374), .A3(new_n658), .ZN(new_n834));
  INV_X1    g648(.A(new_n754), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n801), .B1(new_n835), .B2(KEYINPUT49), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n834), .B(new_n836), .C1(KEYINPUT49), .C2(new_n835), .ZN(new_n837));
  OR3_X1    g651(.A1(new_n733), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n702), .B(KEYINPUT114), .Z(new_n840));
  NAND3_X1  g654(.A1(new_n668), .A2(new_n696), .A3(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n460), .B(new_n679), .C1(new_n577), .C2(new_n576), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n732), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n739), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n527), .A2(new_n747), .A3(new_n689), .ZN(new_n846));
  INV_X1    g660(.A(new_n704), .ZN(new_n847));
  OAI22_X1  g661(.A1(new_n846), .A2(new_n847), .B1(new_n766), .B2(new_n786), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n845), .A2(new_n848), .A3(KEYINPUT52), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  INV_X1    g664(.A(new_n786), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n746), .A2(new_n460), .A3(new_n748), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n851), .A2(new_n852), .B1(new_n697), .B2(new_n704), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n732), .A2(new_n843), .B1(new_n697), .B2(new_n738), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n372), .A2(new_n746), .A3(new_n748), .ZN(new_n857));
  INV_X1    g671(.A(new_n657), .ZN(new_n858));
  INV_X1    g672(.A(new_n767), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n857), .A2(new_n858), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n784), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n763), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n668), .A2(new_n460), .A3(new_n627), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n747), .A2(new_n669), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n673), .A2(new_n689), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n654), .B1(new_n576), .B2(new_n577), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n650), .A2(new_n651), .A3(new_n679), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n633), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n674), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n698), .A2(new_n679), .A3(new_n703), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n747), .A3(new_n689), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n786), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n791), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n797), .A2(new_n799), .A3(new_n872), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n862), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n856), .A2(new_n878), .A3(KEYINPUT53), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT52), .B1(new_n845), .B2(new_n848), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n853), .A2(new_n854), .A3(new_n850), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n749), .A2(new_n657), .B1(new_n766), .B2(new_n767), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n784), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT111), .B1(new_n774), .B2(new_n260), .ZN(new_n886));
  AND4_X1   g700(.A1(KEYINPUT111), .A2(new_n253), .A3(new_n258), .A4(new_n260), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n747), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n738), .A2(new_n668), .A3(new_n793), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT42), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n372), .A2(new_n791), .A3(new_n796), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n890), .A2(new_n891), .A3(new_n799), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n632), .B1(new_n867), .B2(new_n868), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n669), .A3(new_n668), .A4(new_n673), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n628), .A2(new_n894), .A3(new_n692), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n794), .B1(new_n786), .B2(new_n874), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n885), .A2(new_n892), .A3(new_n897), .A4(new_n763), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n880), .B1(new_n883), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n879), .A2(KEYINPUT54), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT54), .B1(new_n879), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n839), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n733), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n793), .A2(new_n620), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n757), .A2(new_n669), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n903), .A2(new_n905), .A3(new_n711), .A4(new_n638), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n754), .A2(new_n658), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n827), .A2(new_n828), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT116), .ZN(new_n909));
  INV_X1    g723(.A(new_n782), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n802), .A2(new_n620), .A3(new_n804), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n912), .B2(new_n790), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT116), .A4(new_n793), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n908), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n805), .A2(new_n757), .A3(new_n904), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n690), .A2(KEYINPUT110), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n918), .A2(new_n356), .A3(new_n689), .A4(new_n780), .ZN(new_n919));
  OR3_X1    g733(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n917), .B1(new_n916), .B2(new_n919), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n906), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT50), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n710), .A2(new_n373), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n757), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n912), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n926), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n928), .A2(KEYINPUT50), .A3(new_n910), .A4(new_n911), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n927), .B2(new_n929), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT51), .B1(new_n923), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT51), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n927), .B2(new_n929), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n906), .A2(new_n915), .A3(new_n936), .A4(new_n922), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n910), .A2(new_n852), .A3(new_n911), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(KEYINPUT119), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n236), .A2(G952), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n938), .B2(KEYINPUT119), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OR3_X1    g756(.A1(new_n916), .A2(KEYINPUT48), .A3(new_n888), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT48), .B1(new_n916), .B2(new_n888), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n903), .B(new_n905), .C1(new_n653), .C2(new_n656), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n937), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n934), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT54), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT53), .B1(new_n856), .B2(new_n878), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n883), .A2(new_n898), .A3(new_n880), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n879), .A2(new_n899), .A3(KEYINPUT54), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n952), .A2(KEYINPUT115), .A3(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n902), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(G952), .A2(G953), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT120), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n838), .B1(new_n955), .B2(new_n957), .ZN(G75));
  NAND2_X1  g772(.A1(new_n879), .A2(new_n899), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n463), .A3(new_n376), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT56), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n413), .A2(new_n426), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT121), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n425), .B(KEYINPUT55), .Z(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n960), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n960), .B2(new_n961), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n236), .A2(G952), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(G51));
  XNOR2_X1  g783(.A(new_n523), .B(KEYINPUT57), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n952), .A2(new_n953), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(KEYINPUT122), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n952), .A2(new_n973), .A3(new_n953), .A4(new_n970), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n742), .B(KEYINPUT123), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n959), .A2(new_n463), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n977), .A2(new_n815), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n968), .B1(new_n976), .B2(new_n978), .ZN(G54));
  NAND2_X1  g793(.A1(KEYINPUT58), .A2(G475), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n562), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n968), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n977), .A2(new_n562), .A3(new_n980), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(G60));
  NOR2_X1   g799(.A1(new_n634), .A2(new_n635), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(G478), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT59), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n952), .A2(new_n987), .A3(new_n953), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n982), .ZN(new_n991));
  INV_X1    g805(.A(new_n954), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT115), .B1(new_n952), .B2(new_n953), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n991), .B1(new_n994), .B2(new_n986), .ZN(G63));
  NAND2_X1  g809(.A1(G217), .A2(G902), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT60), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n879), .B2(new_n899), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n998), .A2(new_n243), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n687), .B(KEYINPUT124), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n999), .A2(new_n982), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT61), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n999), .A2(new_n1001), .A3(KEYINPUT61), .A4(new_n982), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G66));
  OAI21_X1  g820(.A(G953), .B1(new_n622), .B2(new_n423), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n862), .A2(new_n895), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1008), .A2(G953), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT125), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1008), .A2(new_n1011), .A3(G953), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1007), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(KEYINPUT126), .ZN(new_n1014));
  INV_X1    g828(.A(G898), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n963), .B1(new_n1015), .B2(G953), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT126), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1017), .B(new_n1007), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n1014), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1016), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1019), .A2(new_n1020), .ZN(G69));
  OR2_X1    g835(.A1(new_n327), .A2(new_n328), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n531), .A2(new_n532), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1022), .B(new_n1023), .Z(new_n1024));
  NAND2_X1  g838(.A1(G900), .A2(G953), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n853), .A2(new_n739), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n831), .A2(new_n892), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n888), .A2(new_n842), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n822), .A2(new_n714), .A3(new_n1029), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n823), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1024), .B(new_n1025), .C1(new_n1032), .C2(G953), .ZN(new_n1033));
  OAI21_X1  g847(.A(G953), .B1(new_n492), .B2(new_n700), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT127), .Z(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n734), .A2(new_n1027), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT62), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT62), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n734), .A2(new_n1039), .A3(new_n1027), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n372), .A2(new_n793), .A3(new_n869), .ZN(new_n1041));
  OR2_X1    g855(.A1(new_n716), .A2(new_n1041), .ZN(new_n1042));
  AND3_X1   g856(.A1(new_n823), .A2(new_n831), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1038), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n1044), .A2(new_n236), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1033), .B(new_n1036), .C1(new_n1045), .C2(new_n1024), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1032), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1047), .B1(new_n1048), .B2(new_n236), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1024), .B1(new_n1044), .B2(new_n236), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1035), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n1046), .A2(new_n1051), .ZN(G72));
  NAND4_X1  g866(.A1(new_n1038), .A2(new_n1043), .A3(new_n1008), .A4(new_n1040), .ZN(new_n1053));
  NAND2_X1  g867(.A1(G472), .A2(G902), .ZN(new_n1054));
  XOR2_X1   g868(.A(new_n1054), .B(KEYINPUT63), .Z(new_n1055));
  AOI211_X1 g869(.A(new_n335), .B(new_n368), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n368), .A2(new_n336), .ZN(new_n1057));
  INV_X1    g871(.A(new_n341), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1059), .B1(new_n879), .B2(new_n899), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n368), .A2(new_n335), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1028), .A2(new_n1031), .A3(new_n1008), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1061), .B1(new_n1062), .B2(new_n1055), .ZN(new_n1063));
  NOR4_X1   g877(.A1(new_n1056), .A2(new_n1060), .A3(new_n1063), .A4(new_n968), .ZN(G57));
endmodule


