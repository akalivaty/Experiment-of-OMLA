//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G122), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT91), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G122), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT14), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(KEYINPUT95), .A3(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(KEYINPUT14), .B2(new_n193), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT95), .B1(new_n191), .B2(new_n194), .ZN(new_n197));
  OAI21_X1  g011(.A(G107), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT92), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n191), .A2(new_n207), .A3(new_n193), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n207), .B1(new_n191), .B2(new_n193), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n198), .A2(new_n205), .A3(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT9), .B(G234), .ZN(new_n213));
  INV_X1    g027(.A(G217), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n213), .A2(new_n214), .A3(G953), .ZN(new_n215));
  INV_X1    g029(.A(new_n210), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(G107), .A3(new_n208), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT93), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n203), .A2(new_n204), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT94), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n202), .A2(KEYINPUT13), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n200), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n199), .A2(KEYINPUT13), .A3(G128), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n204), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n218), .B1(new_n211), .B2(new_n217), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n212), .B(new_n215), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(G107), .B1(new_n216), .B2(new_n208), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n209), .A2(new_n206), .A3(new_n210), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT93), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n219), .A3(new_n226), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n215), .B1(new_n234), .B2(new_n212), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n187), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G478), .ZN(new_n238));
  INV_X1    g052(.A(G478), .ZN(new_n239));
  OAI221_X1 g053(.A(new_n187), .B1(KEYINPUT15), .B2(new_n239), .C1(new_n230), .C2(new_n235), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT90), .B(G475), .ZN(new_n242));
  INV_X1    g056(.A(G237), .ZN(new_n243));
  INV_X1    g057(.A(G953), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G214), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(G143), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n246), .B(G131), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT17), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n251), .A2(new_n248), .ZN(new_n252));
  XNOR2_X1  g066(.A(G125), .B(G140), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT16), .ZN(new_n254));
  INV_X1    g068(.A(G140), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G125), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(G146), .C1(KEYINPUT16), .C2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n254), .B1(KEYINPUT16), .B2(new_n256), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n249), .A2(new_n252), .A3(new_n257), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT18), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n251), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G140), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT73), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n253), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n269), .A3(new_n259), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n259), .B2(new_n253), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n246), .B1(new_n262), .B2(new_n250), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n263), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n261), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G113), .B(G122), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT89), .B(G104), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n275), .B(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n242), .B1(new_n279), .B2(G902), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n261), .A2(new_n278), .A3(new_n274), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT88), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT19), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n266), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n267), .A2(new_n269), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n283), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n282), .B(new_n257), .C1(new_n286), .C2(G146), .ZN(new_n287));
  INV_X1    g101(.A(new_n247), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n257), .B1(new_n286), .B2(G146), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT88), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n289), .A2(new_n291), .B1(new_n263), .B2(new_n273), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n281), .B1(new_n292), .B2(new_n278), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT20), .ZN(new_n294));
  NOR2_X1   g108(.A1(G475), .A2(G902), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n294), .B1(new_n293), .B2(new_n295), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n280), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(G234), .A2(G237), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n300), .A2(G952), .A3(new_n244), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n300), .A2(G902), .A3(G953), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT21), .B(G898), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n241), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  XNOR2_X1  g120(.A(G116), .B(G119), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT2), .B(G113), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n206), .A2(G104), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n312));
  INV_X1    g126(.A(G104), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G107), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n206), .A2(G104), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT76), .B1(new_n316), .B2(KEYINPUT3), .ZN(new_n317));
  OAI211_X1 g131(.A(KEYINPUT76), .B(KEYINPUT3), .C1(new_n313), .C2(G107), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n315), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G101), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(G107), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n316), .B2(KEYINPUT3), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n314), .B2(new_n312), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n324), .B1(new_n326), .B2(new_n318), .ZN(new_n327));
  INV_X1    g141(.A(G101), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT4), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n315), .B(new_n328), .C1(new_n317), .C2(new_n319), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n310), .B(new_n322), .C1(new_n329), .C2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(new_n316), .B2(new_n323), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n327), .B2(new_n328), .ZN(new_n334));
  INV_X1    g148(.A(new_n307), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n335), .A2(new_n308), .ZN(new_n336));
  INV_X1    g150(.A(G113), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n192), .A2(KEYINPUT5), .A3(G119), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(KEYINPUT82), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n307), .A2(KEYINPUT5), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G116), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n341), .B1(new_n343), .B2(KEYINPUT5), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n339), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n334), .A2(new_n336), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n332), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G110), .B(G122), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n332), .A2(new_n346), .A3(new_n348), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT6), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n353), .A3(new_n349), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n259), .A2(G143), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n199), .A2(G146), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(KEYINPUT0), .A2(G128), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT64), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n199), .B2(G146), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n259), .A2(KEYINPUT64), .A3(G143), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n356), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(KEYINPUT0), .B(G128), .Z(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n355), .B1(new_n366), .B2(new_n264), .ZN(new_n367));
  INV_X1    g181(.A(new_n356), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n357), .A2(KEYINPUT64), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n361), .A2(new_n199), .A3(G146), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n365), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(KEYINPUT83), .B(G125), .C1(new_n373), .C2(new_n360), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n356), .A3(new_n357), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n201), .B1(new_n356), .B2(KEYINPUT1), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n264), .B(new_n376), .C1(new_n371), .C2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n367), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n244), .A2(G224), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n367), .A2(new_n374), .A3(KEYINPUT84), .A4(new_n378), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n352), .B(new_n354), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n382), .A2(KEYINPUT7), .ZN(new_n387));
  AND4_X1   g201(.A1(new_n374), .A2(new_n367), .A3(new_n378), .A4(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n348), .B(KEYINPUT8), .Z(new_n389));
  AOI21_X1  g203(.A(KEYINPUT85), .B1(new_n307), .B2(KEYINPUT5), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n192), .A2(G119), .ZN(new_n391));
  AND4_X1   g205(.A1(KEYINPUT85), .A2(new_n343), .A3(new_n391), .A4(KEYINPUT5), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n344), .B(new_n339), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n334), .A2(new_n336), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n336), .A2(new_n345), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n331), .B2(new_n333), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n389), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n364), .A2(new_n365), .ZN(new_n398));
  INV_X1    g212(.A(new_n360), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G125), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n387), .B1(new_n401), .B2(new_n378), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n388), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(G902), .B1(new_n403), .B2(new_n351), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n386), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT86), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n386), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G210), .B1(G237), .B2(G902), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT87), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n386), .A2(new_n407), .A3(new_n404), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n407), .B1(new_n386), .B2(new_n404), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT87), .B(new_n411), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n386), .A2(new_n410), .A3(new_n404), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n305), .B(new_n306), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G221), .B1(new_n213), .B2(G902), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT75), .ZN(new_n422));
  XOR2_X1   g236(.A(KEYINPUT80), .B(G469), .Z(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  INV_X1    g238(.A(G227), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G953), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n424), .B(new_n426), .Z(new_n427));
  OAI21_X1  g241(.A(new_n376), .B1(new_n371), .B2(new_n377), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n334), .A2(KEYINPUT10), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n366), .B(new_n322), .C1(new_n329), .C2(new_n331), .ZN(new_n430));
  INV_X1    g244(.A(new_n333), .ZN(new_n431));
  INV_X1    g245(.A(new_n358), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n376), .B1(new_n432), .B2(new_n377), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n330), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT10), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n435), .B1(new_n434), .B2(new_n436), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n429), .B(new_n430), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G137), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT11), .B1(new_n440), .B2(G134), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(G134), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g257(.A1(KEYINPUT65), .A2(G137), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT65), .A2(G137), .ZN(new_n445));
  AND2_X1   g259(.A1(KEYINPUT11), .A2(G134), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n443), .A2(new_n447), .A3(new_n250), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n250), .B1(new_n443), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT66), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n204), .A2(G137), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n204), .A2(G137), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(KEYINPUT11), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(KEYINPUT65), .A2(G137), .ZN(new_n454));
  NOR2_X1   g268(.A1(KEYINPUT65), .A2(G137), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT11), .A2(G134), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G131), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n443), .A2(new_n447), .A3(new_n250), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n450), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n439), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT79), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT79), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n439), .A2(new_n465), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n430), .A2(new_n429), .ZN(new_n468));
  INV_X1    g282(.A(new_n462), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(new_n469), .C1(new_n437), .C2(new_n438), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n427), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n470), .A2(new_n427), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n434), .B1(new_n334), .B2(new_n428), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT12), .B1(new_n473), .B2(new_n462), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT78), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n458), .A2(new_n460), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(KEYINPUT12), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n474), .B2(new_n475), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n187), .B(new_n423), .C1(new_n471), .C2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n470), .B1(new_n476), .B2(new_n479), .ZN(new_n483));
  INV_X1    g297(.A(new_n427), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n467), .A2(new_n472), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G469), .B1(new_n485), .B2(G902), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n422), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT81), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n420), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT25), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n201), .A2(G119), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT23), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(KEYINPUT71), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n493), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n342), .A2(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n497), .B2(KEYINPUT71), .ZN(new_n498));
  INV_X1    g312(.A(G110), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n496), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT24), .B(G110), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n498), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n257), .A2(new_n270), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT74), .ZN(new_n504));
  OR3_X1    g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n504), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n498), .A2(new_n499), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n508), .A2(KEYINPUT72), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(KEYINPUT72), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n500), .A2(new_n501), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n260), .A2(new_n257), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT22), .B(G137), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n244), .A2(G221), .A3(G234), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n507), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n507), .B2(new_n513), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n491), .B(new_n187), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n214), .B1(G234), .B2(new_n187), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n520), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n518), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n491), .B1(new_n526), .B2(new_n187), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n522), .A2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(G101), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n243), .A2(new_n244), .A3(G210), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n400), .B1(new_n450), .B2(new_n461), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n204), .B1(new_n454), .B2(new_n455), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n250), .B1(new_n539), .B2(new_n442), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n428), .A2(new_n460), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n538), .A2(new_n543), .A3(new_n310), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT28), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n448), .A2(new_n540), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n428), .A2(new_n547), .B1(new_n477), .B2(new_n366), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(new_n309), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT28), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n537), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT66), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n459), .B1(new_n458), .B2(new_n460), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n366), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n542), .A3(new_n309), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n537), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(KEYINPUT30), .A3(new_n542), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT67), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n398), .B(new_n399), .C1(new_n448), .C2(new_n449), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n542), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT30), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n309), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n560), .B1(new_n559), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n558), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT69), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT31), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n538), .A2(new_n543), .A3(new_n563), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n310), .B1(new_n548), .B2(KEYINPUT30), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT67), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n559), .A2(new_n564), .A3(new_n560), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n557), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT31), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT69), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n573), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n577), .B2(new_n558), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n552), .B(new_n569), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(G472), .A2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT32), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(KEYINPUT32), .A3(new_n580), .ZN(new_n584));
  INV_X1    g398(.A(G472), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n546), .A2(new_n537), .A3(new_n550), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT29), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n544), .B1(new_n572), .B2(new_n573), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n537), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n310), .B1(new_n538), .B2(new_n543), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n556), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n545), .B1(new_n591), .B2(KEYINPUT28), .ZN(new_n592));
  INV_X1    g406(.A(new_n537), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n587), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n585), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n583), .A2(new_n584), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT70), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n580), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n551), .B1(new_n578), .B2(new_n568), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n575), .B(new_n558), .C1(new_n565), .C2(new_n566), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n568), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n567), .A2(KEYINPUT31), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI211_X1 g420(.A(new_n582), .B(new_n601), .C1(new_n602), .C2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT32), .B1(new_n579), .B2(new_n580), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(KEYINPUT70), .A3(new_n597), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n532), .B1(new_n600), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n490), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  NAND2_X1  g427(.A1(new_n482), .A2(new_n486), .ZN(new_n614));
  INV_X1    g428(.A(new_n422), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n488), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n487), .A2(KEYINPUT81), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n585), .B1(new_n579), .B2(new_n187), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n601), .B1(new_n602), .B2(new_n606), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n620), .A2(new_n532), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n306), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n405), .A2(new_n411), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n626), .B2(new_n418), .ZN(new_n627));
  INV_X1    g441(.A(new_n304), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n234), .A2(new_n212), .ZN(new_n630));
  INV_X1    g444(.A(new_n215), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT33), .B1(new_n215), .B2(KEYINPUT96), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n229), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n230), .B2(new_n235), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n239), .A2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n236), .A2(new_n239), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(KEYINPUT97), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT97), .B1(new_n638), .B2(new_n639), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n644), .A3(new_n299), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n638), .A2(new_n639), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT97), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n299), .A3(new_n640), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n629), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n624), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  INV_X1    g468(.A(new_n299), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n241), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n629), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n624), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT35), .B(G107), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NAND2_X1  g475(.A1(new_n507), .A2(new_n513), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n517), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT100), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n662), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n530), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n523), .B2(new_n527), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(KEYINPUT101), .B(new_n666), .C1(new_n523), .C2(new_n527), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n671), .A2(new_n621), .A3(new_n620), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT87), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n419), .B1(new_n675), .B2(new_n415), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n625), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n619), .A2(new_n672), .A3(new_n305), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  NAND2_X1  g494(.A1(new_n600), .A2(new_n610), .ZN(new_n681));
  INV_X1    g495(.A(new_n671), .ZN(new_n682));
  INV_X1    g496(.A(new_n627), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n617), .B2(new_n618), .ZN(new_n684));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n302), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n301), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n655), .A2(new_n241), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n681), .A2(new_n682), .A3(new_n684), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  XNOR2_X1  g507(.A(new_n688), .B(KEYINPUT39), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n489), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n417), .B2(new_n419), .ZN(new_n701));
  INV_X1    g515(.A(new_n700), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n676), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n537), .B1(new_n556), .B2(new_n590), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n187), .B1(new_n574), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G472), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n609), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n667), .ZN(new_n709));
  INV_X1    g523(.A(new_n241), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n655), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n708), .A2(new_n306), .A3(new_n709), .A4(new_n711), .ZN(new_n712));
  OR4_X1    g526(.A1(new_n698), .A2(new_n699), .A3(new_n704), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  NAND4_X1  g528(.A1(new_n648), .A2(new_n299), .A3(new_n640), .A4(new_n688), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n671), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n681), .A2(new_n684), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NOR2_X1   g532(.A1(new_n471), .A2(new_n481), .ZN(new_n719));
  OAI21_X1  g533(.A(G469), .B1(new_n719), .B2(G902), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n482), .ZN(new_n721));
  INV_X1    g535(.A(new_n421), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n611), .A2(new_n651), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND3_X1  g540(.A1(new_n611), .A2(new_n657), .A3(new_n723), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NOR3_X1   g542(.A1(new_n721), .A2(new_n722), .A3(new_n683), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n681), .A2(new_n305), .A3(new_n682), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  NOR2_X1   g545(.A1(new_n592), .A2(new_n537), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n578), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n601), .B1(new_n733), .B2(new_n603), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n620), .A2(new_n532), .A3(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n683), .A2(new_n710), .A3(new_n655), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n723), .A2(new_n735), .A3(new_n628), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  INV_X1    g552(.A(new_n715), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n620), .A2(new_n709), .A3(new_n734), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n729), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  OAI211_X1 g556(.A(new_n306), .B(new_n418), .C1(new_n412), .C2(new_n416), .ZN(new_n743));
  NAND2_X1  g557(.A1(G469), .A2(G902), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n744), .B(KEYINPUT104), .Z(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n485), .B2(G469), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n482), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n743), .A2(new_n722), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n611), .A2(new_n739), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n743), .A2(new_n715), .A3(new_n722), .A4(new_n749), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n584), .A2(KEYINPUT105), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n621), .A2(new_n756), .A3(KEYINPUT32), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n755), .A2(new_n757), .A3(new_n583), .A4(new_n597), .ZN(new_n758));
  INV_X1    g572(.A(new_n532), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n754), .A2(new_n760), .A3(new_n761), .A4(KEYINPUT42), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n625), .B(new_n419), .C1(new_n675), .C2(new_n415), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n739), .A2(new_n763), .A3(new_n421), .A4(new_n748), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n758), .A2(KEYINPUT42), .A3(new_n759), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT106), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n753), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G131), .ZN(G33));
  NAND4_X1  g583(.A1(new_n681), .A2(new_n759), .A3(new_n750), .A4(new_n691), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n643), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT108), .B1(new_n641), .B2(new_n642), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n772), .B(new_n773), .C1(new_n777), .C2(new_n299), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n299), .B1(new_n775), .B2(new_n776), .ZN(new_n779));
  INV_X1    g593(.A(new_n773), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT109), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n299), .B(KEYINPUT110), .Z(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT43), .A3(new_n643), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n667), .B1(new_n620), .B2(new_n621), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n788), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n485), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n485), .A2(new_n793), .ZN(new_n795));
  OAI21_X1  g609(.A(G469), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n745), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n482), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT46), .B1(new_n796), .B2(new_n745), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n421), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n695), .A3(new_n743), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n791), .A2(new_n792), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  XNOR2_X1  g617(.A(new_n800), .B(KEYINPUT47), .ZN(new_n804));
  OR4_X1    g618(.A1(new_n681), .A2(new_n759), .A3(new_n715), .A4(new_n743), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  AOI21_X1  g624(.A(new_n687), .B1(new_n782), .B2(new_n785), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n743), .A2(new_n722), .A3(new_n721), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n740), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n609), .A2(new_n759), .A3(new_n707), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n687), .ZN(new_n815));
  INV_X1    g629(.A(new_n643), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(new_n655), .A3(new_n816), .A4(new_n812), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n721), .B(KEYINPUT114), .Z(new_n819));
  OAI21_X1  g633(.A(new_n804), .B1(new_n615), .B2(new_n819), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n735), .A2(new_n811), .A3(new_n820), .A4(new_n763), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT50), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n811), .A2(new_n735), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n704), .A2(new_n625), .A3(new_n723), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n825), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n811), .A2(KEYINPUT50), .A3(new_n735), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n822), .A2(new_n829), .A3(KEYINPUT51), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n811), .A2(new_n729), .A3(new_n735), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n645), .A2(new_n650), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n815), .A2(new_n834), .A3(new_n812), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(G952), .A3(new_n244), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n811), .A2(new_n760), .A3(new_n812), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT48), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT48), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n811), .A2(new_n839), .A3(new_n760), .A4(new_n812), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n836), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n833), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n833), .B2(new_n841), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n826), .A2(new_n845), .A3(new_n828), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n822), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n826), .B2(new_n828), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI221_X1 g663(.A(new_n830), .B1(new_n843), .B2(new_n844), .C1(new_n849), .C2(KEYINPUT51), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n754), .A2(new_n740), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n241), .A2(new_n299), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n669), .A3(new_n670), .A4(new_n688), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n617), .B2(new_n618), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n681), .A2(new_n763), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n770), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n753), .B2(new_n767), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n304), .B1(new_n649), .B2(new_n656), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n619), .A2(new_n858), .A3(new_n677), .A4(new_n622), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT70), .B1(new_n609), .B2(new_n597), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n607), .A2(new_n608), .A3(new_n599), .A4(new_n596), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n759), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n619), .A2(new_n305), .A3(new_n677), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n678), .B(new_n859), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT112), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n612), .A2(new_n866), .A3(new_n678), .A4(new_n859), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n724), .A2(new_n727), .A3(new_n730), .A4(new_n737), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n857), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT113), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n867), .B2(new_n865), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT113), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n857), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n421), .A2(new_n736), .A3(new_n709), .A4(new_n688), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n708), .A3(new_n748), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n692), .A2(new_n717), .A3(new_n877), .A4(new_n741), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n872), .A2(new_n875), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT53), .B1(new_n880), .B2(new_n881), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n871), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n850), .A2(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n816), .A2(new_n422), .A3(new_n625), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n784), .C1(KEYINPUT49), .C2(new_n721), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(KEYINPUT49), .B2(new_n721), .ZN(new_n897));
  INV_X1    g711(.A(new_n814), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n704), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(G75));
  NOR2_X1   g714(.A1(new_n244), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n187), .B1(new_n887), .B2(new_n891), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT56), .B1(new_n903), .B2(G210), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n384), .A2(new_n385), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n352), .A2(new_n354), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n386), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT55), .Z(new_n909));
  OAI21_X1  g723(.A(new_n902), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n904), .B2(new_n909), .ZN(G51));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n187), .B(new_n796), .C1(new_n887), .C2(new_n891), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n745), .B(KEYINPUT57), .Z(new_n914));
  AOI21_X1  g728(.A(new_n888), .B1(new_n887), .B2(new_n891), .ZN(new_n915));
  AOI211_X1 g729(.A(KEYINPUT54), .B(new_n890), .C1(new_n883), .C2(new_n884), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n719), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n912), .B1(new_n919), .B2(new_n901), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n880), .A2(new_n881), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n871), .B2(KEYINPUT113), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT53), .B1(new_n922), .B2(new_n875), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT54), .B1(new_n923), .B2(new_n890), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n892), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n719), .B1(new_n925), .B2(new_n914), .ZN(new_n926));
  OAI211_X1 g740(.A(KEYINPUT118), .B(new_n902), .C1(new_n926), .C2(new_n913), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n920), .A2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  INV_X1    g743(.A(new_n293), .ZN(new_n930));
  OR3_X1    g744(.A1(new_n929), .A2(KEYINPUT119), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT119), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n901), .B1(new_n929), .B2(new_n930), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(G60));
  AND2_X1   g748(.A1(new_n635), .A2(new_n636), .ZN(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n893), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n925), .A2(new_n935), .A3(new_n937), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n901), .A3(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(new_n887), .A2(new_n891), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT60), .B1(new_n214), .B2(new_n187), .ZN(new_n942));
  OR3_X1    g756(.A1(new_n214), .A2(new_n187), .A3(KEYINPUT60), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n526), .B(KEYINPUT120), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n941), .A2(new_n665), .A3(new_n942), .A4(new_n943), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n902), .A3(new_n947), .ZN(new_n948));
  XOR2_X1   g762(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n949), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n946), .A2(new_n902), .A3(new_n947), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(G66));
  NOR2_X1   g767(.A1(new_n873), .A2(G953), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT122), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(KEYINPUT122), .ZN(new_n956));
  INV_X1    g770(.A(G224), .ZN(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n303), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n906), .B1(G898), .B2(new_n244), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G69));
  OAI21_X1  g775(.A(new_n559), .B1(KEYINPUT30), .B2(new_n548), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n286), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n743), .B1(new_n649), .B2(new_n656), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n611), .A2(new_n696), .A3(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n802), .A2(new_n809), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n692), .A2(new_n717), .A3(new_n741), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT123), .Z(new_n968));
  AOI21_X1  g782(.A(KEYINPUT62), .B1(new_n968), .B2(new_n713), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n968), .A2(KEYINPUT62), .A3(new_n713), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n963), .B1(new_n971), .B2(new_n244), .ZN(new_n972));
  NAND2_X1  g786(.A1(G900), .A2(G953), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n800), .A2(new_n695), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n736), .A3(new_n760), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n770), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n807), .B2(new_n808), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n802), .A3(new_n768), .A4(new_n968), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n963), .B(new_n973), .C1(new_n978), .C2(G953), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT124), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n972), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n425), .B2(new_n685), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G72));
  OAI211_X1 g797(.A(new_n966), .B(new_n873), .C1(new_n969), .C2(new_n970), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT63), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT125), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n588), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n537), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n588), .A2(new_n537), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT126), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n986), .B1(new_n992), .B2(new_n567), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n885), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n873), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n987), .B1(new_n978), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n989), .A2(new_n537), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n901), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n990), .A2(new_n994), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n990), .A2(KEYINPUT127), .A3(new_n994), .A4(new_n998), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(G57));
endmodule


