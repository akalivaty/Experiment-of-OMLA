//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G15gat), .ZN(new_n203));
  INV_X1    g002(.A(G15gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT95), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n203), .A2(new_n205), .A3(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n213), .B1(new_n210), .B2(new_n212), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT96), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n208), .B2(new_n212), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  XNOR2_X1  g017(.A(G43gat), .B(G50gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT93), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n220), .B2(new_n219), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT94), .B(G43gat), .ZN(new_n223));
  INV_X1    g022(.A(G50gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n224), .A2(G43gat), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT15), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT14), .ZN(new_n228));
  INV_X1    g027(.A(G36gat), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n228), .A2(new_n229), .A3(G29gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT14), .B(G29gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n230), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n222), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(new_n222), .B2(new_n232), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n217), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n234), .A2(KEYINPUT17), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n217), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(KEYINPUT17), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n241), .A2(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(KEYINPUT18), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n217), .B(new_n234), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n240), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G169gat), .B(G197gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT92), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G113gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n251));
  INV_X1    g050(.A(G141gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n250), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n254), .B(KEYINPUT12), .Z(new_n255));
  OR2_X1    g054(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n255), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(G50gat), .ZN(new_n261));
  XOR2_X1   g060(.A(G78gat), .B(G106gat), .Z(new_n262));
  XOR2_X1   g061(.A(new_n261), .B(new_n262), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n265));
  INV_X1    g064(.A(G148gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n252), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT73), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n272), .A3(new_n268), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(new_n275), .B2(new_n276), .ZN(new_n281));
  INV_X1    g080(.A(G155gat), .ZN(new_n282));
  INV_X1    g081(.A(G162gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(KEYINPUT74), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n271), .B1(G155gat), .B2(G162gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n269), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT75), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT75), .B1(new_n287), .B2(new_n289), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n278), .B(new_n279), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(KEYINPUT72), .B(KEYINPUT29), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT83), .ZN(new_n295));
  NAND2_X1  g094(.A1(G211gat), .A2(G218gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT22), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(G197gat), .A2(G204gat), .ZN(new_n299));
  AND2_X1   g098(.A1(G197gat), .A2(G204gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G211gat), .B(G218gat), .Z(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n298), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n294), .A2(new_n295), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n287), .A2(new_n289), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT75), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n314), .A2(new_n278), .B1(new_n279), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT82), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319));
  AOI221_X4 g118(.A(new_n319), .B1(new_n316), .B2(new_n279), .C1(new_n314), .C2(new_n278), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n309), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n307), .B1(new_n292), .B2(new_n293), .ZN(new_n322));
  OAI211_X1 g121(.A(G228gat), .B(G233gat), .C1(new_n322), .C2(new_n295), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n265), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n278), .B1(new_n290), .B2(new_n291), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n303), .B2(new_n306), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n325), .B1(KEYINPUT3), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n319), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n325), .B(KEYINPUT82), .C1(KEYINPUT3), .C2(new_n326), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n328), .A2(new_n329), .B1(new_n295), .B2(new_n322), .ZN(new_n330));
  NAND2_X1  g129(.A1(G228gat), .A2(G233gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n294), .A2(new_n308), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(KEYINPUT83), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(KEYINPUT84), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n324), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n277), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT2), .B1(new_n269), .B2(KEYINPUT73), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n273), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n312), .B2(new_n313), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT3), .B1(new_n307), .B2(new_n293), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n342), .A2(new_n331), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n335), .A2(new_n202), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n264), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n202), .B1(new_n335), .B2(new_n344), .ZN(new_n349));
  AOI211_X1 g148(.A(G22gat), .B(new_n343), .C1(new_n324), .C2(new_n334), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT86), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT86), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n321), .A2(new_n265), .A3(new_n323), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT84), .B1(new_n330), .B2(new_n333), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n344), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G22gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n356), .B2(new_n345), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n348), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT86), .B1(new_n349), .B2(new_n350), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n352), .A3(new_n345), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n347), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G127gat), .B(G134gat), .Z(new_n367));
  XNOR2_X1  g166(.A(G113gat), .B(G120gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(KEYINPUT1), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G113gat), .B(G120gat), .Z(new_n370));
  INV_X1    g169(.A(KEYINPUT1), .ZN(new_n371));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n325), .B2(KEYINPUT3), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n366), .B1(new_n375), .B2(new_n292), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n374), .B(new_n278), .C1(new_n290), .C2(new_n291), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT4), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n339), .A2(new_n374), .ZN(new_n382));
  INV_X1    g181(.A(new_n377), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n366), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT5), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT76), .B1(new_n377), .B2(KEYINPUT4), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n339), .A2(new_n387), .A3(new_n388), .A4(new_n374), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n377), .A2(KEYINPUT4), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n376), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n385), .B1(new_n392), .B2(KEYINPUT77), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n376), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n381), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n396), .A2(KEYINPUT87), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(KEYINPUT87), .ZN(new_n398));
  XOR2_X1   g197(.A(KEYINPUT78), .B(KEYINPUT0), .Z(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT79), .ZN(new_n400));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n397), .A2(new_n398), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n404), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT6), .B1(new_n396), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n392), .A2(KEYINPUT77), .ZN(new_n409));
  INV_X1    g208(.A(new_n385), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n395), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n380), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(KEYINPUT6), .A3(new_n404), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT89), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT32), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT23), .ZN(new_n417));
  INV_X1    g216(.A(G169gat), .ZN(new_n418));
  INV_X1    g217(.A(G176gat), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT65), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT65), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(G169gat), .A3(G176gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT25), .ZN(new_n430));
  NAND2_X1  g229(.A1(G183gat), .A2(G190gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT24), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT24), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(G183gat), .A3(G190gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT64), .ZN(new_n436));
  OR3_X1    g235(.A1(new_n436), .A2(G183gat), .A3(G190gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(G183gat), .B2(G190gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n429), .A2(new_n430), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G183gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT27), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT68), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT27), .B(G183gat), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n443), .B(new_n447), .C1(new_n448), .C2(new_n446), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT28), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT66), .B(G190gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n450), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n449), .A2(new_n450), .B1(new_n452), .B2(new_n448), .ZN(new_n453));
  NOR2_X1   g252(.A1(G169gat), .A2(G176gat), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT26), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n427), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n431), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n440), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n435), .B1(new_n451), .B2(G183gat), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n428), .B1(new_n460), .B2(KEYINPUT67), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n435), .B(new_n462), .C1(new_n451), .C2(G183gat), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n430), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n374), .ZN(new_n466));
  INV_X1    g265(.A(new_n374), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n459), .B2(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G227gat), .A2(G233gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n416), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n471), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(G71gat), .B(G99gat), .Z(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G43gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n466), .A2(new_n470), .A3(new_n468), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n481), .B(KEYINPUT34), .Z(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(KEYINPUT33), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n474), .A2(KEYINPUT32), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT69), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT69), .B1(new_n472), .B2(new_n483), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n480), .B(new_n482), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n485), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n472), .A2(KEYINPUT69), .A3(new_n483), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n482), .B1(new_n492), .B2(new_n480), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n415), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n480), .B1(new_n486), .B2(new_n487), .ZN(new_n495));
  INV_X1    g294(.A(new_n482), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT89), .A3(new_n488), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT71), .B1(new_n459), .B2(new_n464), .ZN(new_n499));
  INV_X1    g298(.A(new_n435), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n441), .A2(new_n442), .A3(G183gat), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT67), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n463), .A3(new_n429), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT25), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT71), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n454), .B(KEYINPUT26), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n427), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT68), .B1(new_n444), .B2(KEYINPUT27), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n451), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT27), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G183gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n445), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT68), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT28), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n512), .A2(new_n451), .A3(new_n450), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n431), .B(new_n507), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n504), .A2(new_n505), .A3(new_n516), .A4(new_n440), .ZN(new_n517));
  NAND2_X1  g316(.A1(G226gat), .A2(G233gat), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n518), .B(KEYINPUT70), .Z(new_n519));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(new_n465), .B2(KEYINPUT29), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n307), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n465), .A2(new_n518), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n499), .A2(new_n517), .A3(new_n293), .ZN(new_n524));
  INV_X1    g323(.A(new_n519), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n526), .B2(new_n307), .ZN(new_n527));
  XNOR2_X1  g326(.A(G8gat), .B(G36gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(G64gat), .B(G92gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n528), .B(new_n529), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n522), .B(new_n530), .C1(new_n526), .C2(new_n307), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT30), .A3(new_n533), .ZN(new_n534));
  OR3_X1    g333(.A1(new_n527), .A2(KEYINPUT30), .A3(new_n531), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT35), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n494), .A2(new_n498), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n364), .A2(new_n414), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n534), .A2(new_n535), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT80), .B1(new_n396), .B2(new_n406), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT80), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n412), .A2(new_n541), .A3(new_n404), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n407), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n543), .B2(new_n413), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n497), .A2(new_n488), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n544), .A2(new_n358), .A3(new_n362), .A4(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT90), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT35), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n547), .B2(KEYINPUT35), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n538), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n527), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(KEYINPUT88), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT88), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n527), .B2(KEYINPUT37), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n530), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n527), .A2(KEYINPUT37), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT38), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n526), .A2(new_n308), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n520), .A2(new_n521), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n553), .B1(new_n562), .B2(new_n308), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT38), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n557), .A2(new_n564), .B1(new_n552), .B2(new_n530), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n560), .A2(new_n413), .A3(new_n408), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n375), .A2(new_n292), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n365), .B1(new_n378), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT39), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n404), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n382), .A2(new_n383), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT39), .B1(new_n571), .B2(new_n366), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT40), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n405), .A2(new_n539), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n566), .A2(new_n362), .A3(new_n358), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n543), .A2(new_n413), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI22_X1  g377(.A1(new_n359), .A2(new_n363), .B1(new_n578), .B2(new_n539), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n545), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n497), .A2(KEYINPUT36), .A3(new_n488), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n576), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n259), .B1(new_n551), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT21), .ZN(new_n586));
  XNOR2_X1  g385(.A(G57gat), .B(G64gat), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G71gat), .B(G78gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n217), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT99), .Z(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n593), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT98), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n598), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G85gat), .A2(G92gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT7), .ZN(new_n607));
  NAND2_X1  g406(.A1(G99gat), .A2(G106gat), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  INV_X1    g408(.A(G92gat), .ZN(new_n610));
  AOI22_X1  g409(.A1(KEYINPUT8), .A2(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G99gat), .B(G106gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT101), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n236), .A2(new_n615), .A3(new_n238), .ZN(new_n616));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT100), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT41), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n616), .B(new_n620), .C1(new_n234), .C2(new_n615), .ZN(new_n621));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n619), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n591), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n615), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n614), .B(new_n591), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n632), .B1(new_n638), .B2(KEYINPUT102), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(KEYINPUT102), .B2(new_n638), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n636), .A2(new_n631), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT103), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n637), .A2(new_n632), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n649), .B2(new_n642), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n605), .A2(new_n630), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n585), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n577), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n207), .ZN(G1324gat));
  NAND3_X1  g454(.A1(new_n585), .A2(new_n539), .A3(new_n652), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT16), .B(G8gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT42), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(G8gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT104), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT105), .Z(G1325gat));
  AND3_X1   g462(.A1(new_n581), .A2(KEYINPUT106), .A3(new_n582), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT106), .B1(new_n581), .B2(new_n582), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G15gat), .B1(new_n653), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n494), .A2(new_n498), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n204), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n667), .B1(new_n653), .B2(new_n670), .ZN(G1326gat));
  NOR2_X1   g470(.A1(new_n653), .A2(new_n364), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT107), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT43), .B(G22gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(new_n651), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n605), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n629), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n585), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(G29gat), .A3(new_n577), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT45), .Z(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n629), .A2(new_n682), .ZN(new_n683));
  AND4_X1   g482(.A1(new_n362), .A2(new_n537), .A3(new_n358), .A4(new_n414), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT90), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT35), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n576), .A2(new_n579), .A3(new_n583), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n259), .A2(new_n677), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n576), .A2(new_n666), .A3(new_n579), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n629), .B1(new_n551), .B2(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n690), .B(new_n691), .C1(new_n693), .C2(KEYINPUT44), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n577), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n681), .A2(new_n695), .ZN(G1328gat));
  INV_X1    g495(.A(new_n539), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n679), .A2(G36gat), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n694), .B2(new_n697), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  NOR2_X1   g500(.A1(new_n668), .A2(new_n223), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT108), .B1(new_n679), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n585), .A2(new_n705), .A3(new_n678), .A4(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n223), .B1(new_n694), .B2(new_n666), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n694), .B2(new_n666), .ZN(new_n713));
  INV_X1    g512(.A(new_n683), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n551), .B2(new_n584), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n576), .A2(new_n666), .A3(new_n579), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n630), .B1(new_n688), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n715), .B1(new_n717), .B2(new_n682), .ZN(new_n718));
  INV_X1    g517(.A(new_n666), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n718), .A2(KEYINPUT109), .A3(new_n719), .A4(new_n691), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n713), .A2(new_n720), .A3(new_n223), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n710), .B1(new_n704), .B2(new_n706), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n721), .A2(KEYINPUT110), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT110), .B1(new_n721), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n711), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT111), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n711), .B(new_n727), .C1(new_n723), .C2(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(G1330gat));
  OAI21_X1  g528(.A(new_n224), .B1(new_n679), .B2(new_n364), .ZN(new_n730));
  INV_X1    g529(.A(new_n364), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G50gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n694), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g533(.A1(new_n605), .A2(new_n630), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n259), .A2(new_n735), .A3(new_n651), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n551), .B2(new_n692), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n578), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT112), .B(G57gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n539), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT49), .B(G64gat), .Z(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(G1333gat));
  NAND3_X1  g543(.A1(new_n737), .A2(G71gat), .A3(new_n719), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT113), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n737), .A2(new_n669), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748));
  AOI21_X1  g547(.A(G71gat), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n748), .B2(new_n747), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n731), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  INV_X1    g553(.A(new_n605), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n258), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n693), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT51), .Z(new_n758));
  NAND4_X1  g557(.A1(new_n758), .A2(new_n609), .A3(new_n578), .A4(new_n651), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n718), .A2(new_n651), .A3(new_n756), .ZN(new_n760));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n577), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1336gat));
  NAND3_X1  g561(.A1(new_n651), .A2(new_n539), .A3(new_n610), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT115), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n758), .A2(new_n764), .B1(KEYINPUT116), .B2(KEYINPUT52), .ZN(new_n765));
  OAI21_X1  g564(.A(G92gat), .B1(new_n760), .B2(new_n697), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT117), .Z(new_n769));
  XNOR2_X1  g568(.A(new_n767), .B(new_n769), .ZN(G1337gat));
  NOR3_X1   g569(.A1(new_n668), .A2(new_n676), .A3(G99gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n758), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G99gat), .B1(new_n760), .B2(new_n666), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(G1338gat));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n364), .A2(G106gat), .A3(new_n676), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT118), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G106gat), .B1(new_n760), .B2(new_n364), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n779), .B(new_n781), .ZN(G1339gat));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n649), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n646), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n637), .B2(new_n632), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n640), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n648), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n787), .A2(KEYINPUT55), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n258), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n239), .A2(new_n240), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n244), .A2(new_n245), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n254), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n256), .A2(new_n651), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n630), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  AND4_X1   g596(.A1(new_n256), .A2(new_n791), .A3(new_n630), .A4(new_n795), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n605), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n652), .A2(new_n259), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n731), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n802), .A2(new_n578), .A3(new_n697), .A4(new_n669), .ZN(new_n803));
  INV_X1    g602(.A(G113gat), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n803), .A2(new_n804), .A3(new_n259), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n801), .A2(new_n577), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n364), .A3(new_n546), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n539), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n258), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n805), .B1(new_n809), .B2(new_n804), .ZN(G1340gat));
  INV_X1    g609(.A(G120gat), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n803), .A2(new_n811), .A3(new_n676), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n651), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(new_n811), .ZN(G1341gat));
  INV_X1    g613(.A(G127gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n808), .A2(new_n815), .A3(new_n755), .ZN(new_n816));
  OAI21_X1  g615(.A(G127gat), .B1(new_n803), .B2(new_n605), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1342gat));
  NAND2_X1  g617(.A1(new_n630), .A2(new_n697), .ZN(new_n819));
  OR3_X1    g618(.A1(new_n807), .A2(G134gat), .A3(new_n819), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n821));
  OAI21_X1  g620(.A(G134gat), .B1(new_n803), .B2(new_n629), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(G1343gat));
  NAND2_X1  g623(.A1(new_n578), .A2(new_n697), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n719), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n787), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n258), .A2(new_n648), .A3(new_n788), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n630), .B1(new_n830), .B2(new_n796), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n605), .B1(new_n831), .B2(new_n798), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n832), .A2(new_n833), .B1(new_n259), .B2(new_n652), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n364), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n801), .B2(new_n364), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n827), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n258), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G141gat), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n806), .A2(new_n731), .A3(new_n666), .ZN(new_n845));
  NOR4_X1   g644(.A1(new_n845), .A2(G141gat), .A3(new_n259), .A4(new_n539), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n252), .B1(new_n841), .B2(new_n258), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT58), .B1(new_n849), .B2(new_n846), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1344gat));
  NOR2_X1   g650(.A1(new_n845), .A2(new_n539), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n266), .A3(new_n651), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n826), .A2(new_n651), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n832), .A2(new_n800), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n837), .B1(new_n856), .B2(new_n364), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n799), .A2(new_n800), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n838), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n855), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT121), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n266), .B1(new_n860), .B2(KEYINPUT121), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n854), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT59), .B(new_n266), .C1(new_n841), .C2(new_n651), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n853), .B1(new_n863), .B2(new_n864), .ZN(G1345gat));
  AOI21_X1  g664(.A(G155gat), .B1(new_n852), .B2(new_n755), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n605), .A2(new_n282), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT122), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n841), .B2(new_n868), .ZN(G1346gat));
  AOI21_X1  g668(.A(new_n283), .B1(new_n841), .B2(new_n630), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n845), .A2(G162gat), .A3(new_n819), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n870), .A2(new_n871), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n578), .A2(new_n697), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n668), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n802), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n418), .A3(new_n259), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n577), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(KEYINPUT123), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(KEYINPUT123), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR4_X1   g680(.A1(new_n881), .A2(new_n697), .A3(new_n731), .A4(new_n545), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n258), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(new_n418), .ZN(G1348gat));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n419), .A3(new_n651), .ZN(new_n885));
  OAI21_X1  g684(.A(G176gat), .B1(new_n876), .B2(new_n676), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1349gat));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n876), .B2(new_n605), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n802), .A2(KEYINPUT124), .A3(new_n755), .A4(new_n875), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(G183gat), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n731), .A2(new_n697), .A3(new_n545), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n605), .A2(new_n512), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n893), .B(new_n894), .C1(new_n879), .C2(new_n880), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT60), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n891), .A2(new_n892), .A3(new_n898), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n443), .A3(new_n630), .ZN(new_n901));
  OAI21_X1  g700(.A(G190gat), .B1(new_n876), .B2(new_n629), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n902), .A2(KEYINPUT61), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(KEYINPUT61), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(G1351gat));
  NAND2_X1  g704(.A1(new_n857), .A2(new_n859), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n719), .A2(new_n874), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G197gat), .B1(new_n908), .B2(new_n259), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n666), .A2(new_n731), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n881), .A2(new_n697), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n259), .A2(G197gat), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n909), .B1(new_n914), .B2(new_n915), .ZN(G1352gat));
  XOR2_X1   g715(.A(KEYINPUT127), .B(G204gat), .Z(new_n917));
  NOR2_X1   g716(.A1(new_n676), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT62), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n908), .B2(new_n676), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n911), .A2(new_n922), .A3(new_n918), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(G1353gat));
  INV_X1    g723(.A(G211gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n911), .A2(new_n925), .A3(new_n755), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n755), .A3(new_n907), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1354gat));
  INV_X1    g729(.A(G218gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n911), .A2(new_n931), .A3(new_n630), .ZN(new_n932));
  OAI21_X1  g731(.A(G218gat), .B1(new_n908), .B2(new_n629), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1355gat));
endmodule


