//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT3), .A2(G107), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT3), .A2(G107), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(G104), .B2(new_n190), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT79), .A2(G104), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT79), .A2(G104), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n191), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n196), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT79), .A2(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n194), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n194), .A2(G104), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n198), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT80), .B1(new_n199), .B2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(G107), .B1(new_n192), .B2(new_n196), .ZN(new_n207));
  OAI21_X1  g021(.A(G101), .B1(new_n207), .B2(new_n203), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n191), .A2(new_n197), .A3(new_n198), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT10), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n213), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(G143), .B2(new_n214), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n221), .B1(new_n223), .B2(new_n213), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n212), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n206), .A2(new_n211), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT11), .ZN(new_n227));
  INV_X1    g041(.A(G134), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(G137), .ZN(new_n229));
  INV_X1    g043(.A(G137), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT11), .A3(G134), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G131), .ZN(new_n234));
  INV_X1    g048(.A(G131), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n229), .A2(new_n231), .A3(new_n235), .A4(new_n232), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n200), .A2(new_n201), .A3(new_n190), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G107), .ZN(new_n242));
  INV_X1    g056(.A(G104), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n195), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(G101), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n217), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT0), .B(G128), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n221), .A2(new_n250), .A3(KEYINPUT65), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(G101), .C1(new_n241), .C2(new_n244), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n246), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n208), .A2(new_n209), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n216), .A2(new_n217), .ZN(new_n257));
  AND4_X1   g071(.A1(new_n222), .A2(new_n215), .A3(new_n220), .A4(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n212), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n226), .A2(new_n240), .A3(new_n255), .A4(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G110), .B(G140), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT78), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G227), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n263), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n259), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n206), .B2(new_n211), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n256), .A2(new_n259), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n239), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(KEYINPUT12), .B(new_n239), .C1(new_n269), .C2(new_n270), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n267), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n226), .A2(new_n255), .A3(new_n260), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n276), .A2(new_n277), .A3(new_n239), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n276), .B2(new_n239), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n261), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n266), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT74), .B(G902), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n282), .A2(G469), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G469), .ZN(new_n286));
  INV_X1    g100(.A(new_n267), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n278), .B2(new_n279), .ZN(new_n288));
  INV_X1    g102(.A(new_n261), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n273), .B2(new_n274), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n290), .B2(new_n266), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n188), .B1(new_n285), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT82), .ZN(new_n295));
  INV_X1    g109(.A(G237), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n264), .A3(G214), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(KEYINPUT87), .A3(new_n219), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n219), .A2(KEYINPUT87), .ZN(new_n299));
  NOR2_X1   g113(.A1(G237), .A2(G953), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(G214), .A3(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n298), .A2(new_n301), .B1(KEYINPUT18), .B2(G131), .ZN(new_n302));
  AND4_X1   g116(.A1(KEYINPUT18), .A2(new_n298), .A3(G131), .A4(new_n301), .ZN(new_n303));
  XNOR2_X1  g117(.A(G125), .B(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n214), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT75), .A2(G125), .ZN(new_n306));
  INV_X1    g120(.A(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(G146), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT88), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n305), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(new_n305), .B2(new_n310), .ZN(new_n313));
  OAI22_X1  g127(.A1(new_n302), .A2(new_n303), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI221_X1 g130(.A(KEYINPUT89), .B1(new_n312), .B2(new_n313), .C1(new_n302), .C2(new_n303), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G113), .B(G122), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT91), .B(G104), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n319), .B(new_n320), .Z(new_n321));
  NAND2_X1  g135(.A1(new_n298), .A2(new_n301), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT17), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n298), .A2(new_n235), .A3(new_n301), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n327), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n328), .A2(KEYINPUT76), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n308), .A2(new_n309), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT16), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(KEYINPUT76), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n214), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n329), .A2(new_n331), .A3(G146), .A4(new_n332), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n322), .A2(KEYINPUT17), .A3(G131), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n326), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n318), .A2(new_n321), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n321), .B1(new_n318), .B2(new_n337), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n292), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G475), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n323), .A2(new_n325), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT19), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n304), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n308), .A2(KEYINPUT19), .A3(new_n309), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n345), .A2(KEYINPUT90), .A3(new_n214), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n335), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT90), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n346), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(G146), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n316), .A2(new_n317), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n338), .B1(new_n353), .B2(new_n321), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n355));
  NOR2_X1   g169(.A1(G475), .A2(G902), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n354), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n342), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI211_X1 g174(.A(new_n264), .B(new_n283), .C1(G234), .C2(G237), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT21), .B(G898), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G952), .ZN(new_n364));
  AOI211_X1 g178(.A(G953), .B(new_n364), .C1(G234), .C2(G237), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G128), .B(G143), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n228), .ZN(new_n369));
  INV_X1    g183(.A(G116), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT14), .A3(G122), .ZN(new_n371));
  XNOR2_X1  g185(.A(G116), .B(G122), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(G107), .B(new_n371), .C1(new_n373), .C2(KEYINPUT14), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n369), .B(new_n374), .C1(G107), .C2(new_n373), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n368), .A2(KEYINPUT13), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n219), .A2(G128), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n376), .B(G134), .C1(KEYINPUT13), .C2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n372), .B(new_n194), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n368), .A2(new_n228), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G217), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n187), .A2(new_n382), .A3(G953), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n375), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n383), .B1(new_n375), .B2(new_n381), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT92), .B1(new_n386), .B2(new_n284), .ZN(new_n387));
  INV_X1    g201(.A(G478), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(KEYINPUT15), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT92), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n390), .B(new_n283), .C1(new_n384), .C2(new_n385), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  OAI221_X1 g206(.A(new_n283), .B1(KEYINPUT15), .B2(new_n388), .C1(new_n384), .C2(new_n385), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n360), .A2(new_n367), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G214), .B1(G237), .B2(G902), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT2), .B(G113), .Z(new_n398));
  XNOR2_X1  g212(.A(G116), .B(G119), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n370), .A2(G119), .ZN(new_n401));
  INV_X1    g215(.A(G119), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G116), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT5), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n404), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G113), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n400), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n206), .A2(new_n409), .A3(new_n211), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT85), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n256), .A2(new_n412), .A3(new_n408), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n256), .B2(new_n408), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n206), .A2(new_n409), .A3(new_n416), .A4(new_n211), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT8), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n398), .B(new_n399), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n246), .A2(new_n422), .A3(new_n254), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n410), .A2(new_n423), .A3(new_n419), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n252), .A2(G125), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(G125), .B2(new_n259), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n264), .A2(G224), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(KEYINPUT7), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(KEYINPUT7), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n425), .B(new_n429), .C1(G125), .C2(new_n259), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n424), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G210), .B1(G237), .B2(G902), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n427), .B(KEYINPUT84), .Z(new_n434));
  XNOR2_X1  g248(.A(new_n426), .B(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n410), .A2(new_n423), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n419), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n424), .A2(KEYINPUT6), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n436), .A2(KEYINPUT6), .A3(new_n438), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n432), .A2(new_n433), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n433), .B1(new_n432), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n397), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n446), .B(new_n188), .C1(new_n285), .C2(new_n293), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n295), .A2(new_n396), .A3(new_n445), .A4(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n239), .A2(new_n252), .ZN(new_n451));
  INV_X1    g265(.A(new_n422), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n236), .B(KEYINPUT66), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n230), .A2(G134), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n235), .B1(new_n454), .B2(new_n232), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n218), .B2(new_n224), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT28), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT66), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n236), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n455), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n257), .B2(new_n258), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT67), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT67), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n453), .A2(new_n456), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n451), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n422), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n300), .A2(G210), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT27), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT26), .B(G101), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n451), .A2(KEYINPUT30), .A3(new_n457), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n451), .A2(KEYINPUT69), .A3(KEYINPUT30), .A4(new_n457), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n467), .A2(KEYINPUT68), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT68), .B1(new_n467), .B2(new_n480), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n422), .B(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n458), .A2(new_n473), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT70), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT31), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT31), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n474), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(G472), .A2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n450), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT31), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT31), .B1(new_n483), .B2(new_n485), .ZN(new_n496));
  OAI22_X1  g310(.A1(new_n495), .A2(new_n496), .B1(new_n473), .B2(new_n469), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT71), .A3(new_n491), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(KEYINPUT32), .A3(new_n491), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n483), .A2(new_n458), .ZN(new_n501));
  INV_X1    g315(.A(new_n473), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT72), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n469), .A2(new_n473), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT29), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT72), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n507), .B(new_n473), .C1(new_n483), .C2(new_n458), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n503), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n451), .A2(new_n457), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT28), .B1(new_n510), .B2(new_n452), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n458), .A2(KEYINPUT73), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n451), .A2(new_n513), .A3(new_n452), .A4(new_n457), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n512), .B(new_n514), .C1(new_n452), .C2(new_n510), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n511), .B1(new_n515), .B2(KEYINPUT28), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n502), .A2(new_n505), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n284), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G472), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n499), .A2(new_n500), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n382), .B1(new_n283), .B2(G234), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n334), .A2(new_n335), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n213), .A2(KEYINPUT23), .A3(G119), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n402), .A2(G128), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n402), .A2(G128), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(KEYINPUT23), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G110), .ZN(new_n530));
  INV_X1    g344(.A(new_n528), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n531), .A2(new_n527), .ZN(new_n532));
  XOR2_X1   g346(.A(KEYINPUT24), .B(G110), .Z(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n525), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  OAI22_X1  g349(.A1(new_n532), .A2(new_n533), .B1(G110), .B2(new_n529), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n335), .A3(new_n305), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT77), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT22), .B(G137), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n535), .A2(new_n537), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n524), .B1(new_n546), .B2(new_n284), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n544), .A2(KEYINPUT25), .A3(new_n283), .A4(new_n545), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n523), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n522), .A2(G902), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n551), .A3(new_n545), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n449), .A2(new_n521), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(G101), .ZN(G3));
  NAND3_X1  g369(.A1(new_n295), .A2(new_n553), .A3(new_n447), .ZN(new_n556));
  OAI21_X1  g370(.A(G472), .B1(new_n490), .B2(new_n284), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n493), .A2(new_n557), .A3(new_n498), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n559), .B(KEYINPUT93), .Z(new_n560));
  INV_X1    g374(.A(KEYINPUT33), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n386), .A2(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT33), .ZN(new_n563));
  OAI211_X1 g377(.A(G478), .B(new_n283), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n359), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n397), .B(new_n367), .C1(new_n442), .C2(new_n443), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT34), .B(G104), .Z(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(G6));
  NOR3_X1   g386(.A1(new_n568), .A2(new_n359), .A3(new_n395), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n560), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G107), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT94), .B(KEYINPUT35), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G9));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n542), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT95), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n580), .A2(new_n538), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n538), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n551), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n549), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n493), .A2(new_n557), .A3(new_n498), .A4(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n448), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT37), .B(G110), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G12));
  INV_X1    g404(.A(G900), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n365), .B1(new_n361), .B2(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n359), .A2(new_n395), .A3(new_n592), .ZN(new_n593));
  AND4_X1   g407(.A1(new_n445), .A2(new_n295), .A3(new_n447), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n521), .A3(new_n586), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT96), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n594), .A2(new_n521), .A3(new_n597), .A4(new_n586), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G128), .ZN(G30));
  AND2_X1   g414(.A1(new_n295), .A2(new_n447), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n592), .B(KEYINPUT39), .Z(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n603), .B(KEYINPUT40), .Z(new_n604));
  AOI22_X1  g418(.A1(new_n483), .A2(new_n485), .B1(new_n502), .B2(new_n515), .ZN(new_n605));
  OAI21_X1  g419(.A(G472), .B1(new_n605), .B2(G902), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n499), .A2(new_n500), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n442), .A2(new_n443), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT97), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT99), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n608), .B(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n397), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n359), .A2(new_n394), .ZN(new_n614));
  NOR4_X1   g428(.A1(new_n612), .A2(new_n613), .A3(new_n586), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n604), .A2(new_n607), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT100), .B(G143), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G45));
  NOR2_X1   g432(.A1(new_n567), .A2(new_n592), .ZN(new_n619));
  AND4_X1   g433(.A1(new_n445), .A2(new_n295), .A3(new_n447), .A4(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(new_n521), .A3(new_n586), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G146), .ZN(G48));
  NOR2_X1   g436(.A1(new_n286), .A2(KEYINPUT101), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n282), .B2(new_n284), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n273), .A2(new_n274), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n287), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n276), .A2(new_n239), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT81), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n276), .A2(new_n277), .A3(new_n239), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n289), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n626), .B1(new_n630), .B2(new_n266), .ZN(new_n631));
  INV_X1    g445(.A(new_n623), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(new_n283), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n624), .A2(new_n633), .A3(new_n188), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n521), .A2(new_n553), .A3(new_n569), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT41), .B(G113), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G15));
  NAND4_X1  g452(.A1(new_n521), .A2(new_n553), .A3(new_n573), .A4(new_n635), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT102), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n370), .ZN(G18));
  OR3_X1    g455(.A1(new_n634), .A2(KEYINPUT103), .A3(new_n444), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT103), .B1(new_n634), .B2(new_n444), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n521), .A2(new_n644), .A3(new_n396), .A4(new_n586), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT104), .B(G119), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G21));
  NOR3_X1   g461(.A1(new_n634), .A2(new_n614), .A3(new_n568), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n502), .B1(new_n516), .B2(KEYINPUT105), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(KEYINPUT105), .B2(new_n516), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n495), .A2(new_n496), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n491), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n648), .A2(new_n553), .A3(new_n557), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G122), .ZN(G24));
  AND3_X1   g468(.A1(new_n652), .A2(new_n557), .A3(new_n586), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n644), .A2(new_n655), .A3(new_n619), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G125), .ZN(G27));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n658));
  INV_X1    g472(.A(new_n553), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n494), .B1(new_n490), .B2(new_n492), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n500), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n503), .A2(new_n508), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT29), .B1(new_n469), .B2(new_n473), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n518), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n661), .A2(KEYINPUT106), .B1(new_n665), .B2(G472), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n661), .A2(KEYINPUT106), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n659), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n608), .A2(new_n397), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n294), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n619), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n658), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n521), .A2(new_n553), .A3(new_n670), .ZN(new_n673));
  INV_X1    g487(.A(new_n619), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n673), .A2(KEYINPUT42), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT107), .B(G131), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G33));
  NAND4_X1  g492(.A1(new_n521), .A2(new_n553), .A3(new_n593), .A4(new_n670), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G134), .ZN(G36));
  NAND2_X1  g494(.A1(new_n360), .A2(new_n566), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n359), .B2(KEYINPUT109), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n585), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n558), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n669), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n286), .B1(new_n291), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n689), .B2(new_n291), .ZN(new_n691));
  NAND2_X1  g505(.A1(G469), .A2(G902), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n694));
  OR3_X1    g508(.A1(new_n693), .A2(KEYINPUT108), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT108), .B1(new_n693), .B2(new_n694), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n285), .B1(new_n693), .B2(new_n694), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n698), .A2(new_n188), .A3(new_n602), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n688), .B(new_n699), .C1(new_n687), .C2(new_n686), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G137), .ZN(G39));
  NAND2_X1  g515(.A1(new_n698), .A2(new_n188), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT47), .ZN(new_n703));
  OR4_X1    g517(.A1(new_n553), .A2(new_n521), .A3(new_n674), .A4(new_n669), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G140), .ZN(G42));
  AND2_X1   g520(.A1(new_n624), .A2(new_n633), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n703), .B1(new_n188), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n684), .A2(new_n366), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n553), .A3(new_n557), .A4(new_n652), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n669), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT115), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT117), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n612), .A2(new_n613), .A3(new_n635), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n717), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n634), .A2(new_n669), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n711), .A2(new_n655), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n607), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n553), .A3(new_n365), .A4(new_n723), .ZN(new_n726));
  OR3_X1    g540(.A1(new_n726), .A2(new_n359), .A3(new_n566), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n721), .A2(new_n722), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n715), .A2(new_n716), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n668), .A2(new_n711), .A3(new_n723), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n730), .B(KEYINPUT48), .Z(new_n731));
  NOR2_X1   g545(.A1(new_n364), .A2(G953), .ZN(new_n732));
  INV_X1    g546(.A(new_n644), .ZN(new_n733));
  OAI221_X1 g547(.A(new_n732), .B1(new_n726), .B2(new_n567), .C1(new_n733), .C2(new_n712), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n729), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n715), .B(KEYINPUT116), .Z(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n728), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n738));
  OAI21_X1  g552(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n653), .B1(new_n448), .B2(new_n587), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n395), .A2(KEYINPUT111), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n394), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n359), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n359), .A2(new_n566), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n445), .B(new_n367), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n556), .A2(new_n558), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n554), .A3(new_n636), .A4(new_n645), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n640), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n656), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n596), .B2(new_n598), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n549), .A2(new_n584), .A3(new_n592), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n754), .B(new_n188), .C1(new_n285), .C2(new_n293), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT113), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n755), .A2(KEYINPUT113), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n614), .A2(new_n444), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n607), .A2(new_n756), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n759), .A2(new_n621), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n752), .A2(new_n753), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n741), .A2(new_n743), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n669), .A2(new_n359), .A3(new_n762), .A4(new_n592), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n521), .A2(new_n601), .A3(new_n586), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n671), .A2(new_n655), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n679), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n672), .A2(new_n675), .A3(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n750), .A2(new_n761), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n621), .B1(new_n752), .B2(KEYINPUT112), .ZN(new_n769));
  INV_X1    g583(.A(new_n759), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n771), .B(new_n751), .C1(new_n596), .C2(new_n598), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT53), .B(new_n768), .C1(new_n773), .C2(new_n753), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n750), .A2(new_n761), .A3(new_n767), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n753), .B1(new_n752), .B2(new_n760), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n774), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n777), .A2(new_n776), .A3(new_n778), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n768), .B1(new_n773), .B2(new_n753), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(new_n776), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n780), .B1(new_n783), .B2(new_n775), .ZN(new_n784));
  OAI22_X1  g598(.A1(new_n739), .A2(new_n784), .B1(G952), .B2(G953), .ZN(new_n785));
  INV_X1    g599(.A(new_n681), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n553), .A3(new_n397), .A4(new_n188), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n612), .B1(new_n788), .B2(KEYINPUT110), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n707), .B(KEYINPUT49), .Z(new_n792));
  OR3_X1    g606(.A1(new_n789), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n785), .B1(new_n607), .B2(new_n793), .ZN(G75));
  NOR2_X1   g608(.A1(new_n264), .A2(G952), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n283), .B1(new_n774), .B2(new_n779), .ZN(new_n797));
  INV_X1    g611(.A(new_n433), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n439), .A2(new_n440), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(new_n435), .Z(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT55), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n796), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n799), .B2(new_n802), .ZN(G51));
  NAND2_X1  g618(.A1(new_n774), .A2(new_n779), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT54), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n780), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n692), .B(KEYINPUT57), .Z(new_n808));
  AOI21_X1  g622(.A(new_n282), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n691), .B(KEYINPUT118), .Z(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(new_n284), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n797), .A2(KEYINPUT119), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n796), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT120), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n818), .B(new_n796), .C1(new_n809), .C2(new_n815), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(G54));
  NAND3_X1  g634(.A1(new_n797), .A2(KEYINPUT58), .A3(G475), .ZN(new_n821));
  INV_X1    g635(.A(new_n354), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n824), .A3(new_n795), .ZN(G60));
  NOR2_X1   g639(.A1(new_n562), .A2(new_n563), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(G478), .A2(G902), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT59), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n827), .B1(new_n784), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n827), .A2(new_n829), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n795), .B(new_n830), .C1(new_n807), .C2(new_n831), .ZN(G63));
  XNOR2_X1  g646(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n382), .A2(new_n292), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n805), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n795), .B1(new_n836), .B2(new_n546), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n581), .A2(new_n582), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n837), .B1(new_n838), .B2(new_n836), .ZN(new_n839));
  XNOR2_X1  g653(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(G66));
  INV_X1    g655(.A(G224), .ZN(new_n842));
  OAI21_X1  g656(.A(G953), .B1(new_n362), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n750), .B2(G953), .ZN(new_n844));
  INV_X1    g658(.A(G898), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n800), .B1(new_n845), .B2(G953), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT123), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n844), .B(new_n847), .ZN(G69));
  OAI21_X1  g662(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n351), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n591), .A2(G953), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT125), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n699), .A2(new_n668), .A3(new_n758), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n705), .A2(new_n679), .A3(new_n700), .A4(new_n853), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n854), .A2(new_n676), .A3(new_n772), .A4(new_n769), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n850), .B(new_n852), .C1(new_n855), .C2(G953), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n744), .A2(new_n745), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n603), .A2(new_n669), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n553), .A3(new_n521), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n705), .A2(new_n700), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n769), .A2(new_n772), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n616), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(KEYINPUT62), .A3(new_n616), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n850), .A2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n856), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT124), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n264), .B1(G227), .B2(G900), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n869), .B(new_n870), .ZN(G72));
  NAND2_X1  g685(.A1(new_n855), .A2(new_n750), .ZN(new_n872));
  NAND2_X1  g686(.A1(G472), .A2(G902), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT63), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n501), .B(KEYINPUT126), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n473), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n795), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n662), .A2(KEYINPUT127), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n662), .A2(KEYINPUT127), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n486), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n874), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n878), .B1(new_n783), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n876), .A2(new_n473), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n866), .A2(new_n750), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n884), .B1(new_n885), .B2(new_n874), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n883), .A2(new_n886), .ZN(G57));
endmodule


