//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  AND2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT80), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT80), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G155gat), .B2(G162gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n203), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(G141gat), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(G148gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(G148gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(G141gat), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n218), .A2(new_n219), .B1(KEYINPUT2), .B2(new_n210), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(KEYINPUT81), .A3(new_n210), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT81), .ZN(new_n223));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n203), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n220), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G120gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G113gat), .ZN(new_n229));
  INV_X1    g028(.A(G113gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G120gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n232), .B(new_n233), .C1(new_n234), .C2(KEYINPUT70), .ZN(new_n235));
  INV_X1    g034(.A(G127gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G134gat), .ZN(new_n237));
  INV_X1    g036(.A(G134gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G127gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(KEYINPUT70), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n240), .B(new_n241), .C1(new_n242), .C2(KEYINPUT1), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n227), .A2(KEYINPUT83), .A3(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n217), .A2(new_n226), .A3(new_n235), .A4(new_n243), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT87), .ZN(new_n250));
  INV_X1    g049(.A(new_n246), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n250), .B1(new_n249), .B2(new_n253), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n217), .A2(new_n226), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n235), .A2(new_n243), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n217), .A2(new_n226), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n257), .A2(KEYINPUT5), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n246), .B(KEYINPUT83), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT84), .B1(new_n227), .B2(new_n244), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n258), .A2(new_n271), .A3(new_n260), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n264), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n268), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n258), .A2(new_n271), .A3(new_n260), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n271), .B1(new_n258), .B2(new_n260), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n248), .B(new_n245), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n264), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(KEYINPUT85), .A3(KEYINPUT5), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n245), .A2(new_n248), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n251), .A2(new_n252), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n265), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT86), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT86), .ZN(new_n291));
  AOI211_X1 g090(.A(new_n291), .B(new_n288), .C1(new_n276), .C2(new_n282), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n267), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G1gat), .B(G29gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT0), .ZN(new_n295));
  XNOR2_X1  g094(.A(G57gat), .B(G85gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n279), .A2(new_n280), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT39), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n263), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n249), .A2(new_n253), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT87), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n304), .B2(new_n254), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n301), .B1(new_n305), .B2(new_n264), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n263), .B1(new_n255), .B2(new_n256), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(new_n300), .A3(new_n280), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n306), .A2(new_n297), .A3(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n293), .A2(new_n298), .B1(new_n309), .B2(KEYINPUT40), .ZN(new_n310));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(G183gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT27), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G183gat), .ZN(new_n315));
  INV_X1    g114(.A(G190gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT27), .B(G183gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(KEYINPUT28), .A3(new_n316), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n325));
  INV_X1    g124(.A(G169gat), .ZN(new_n326));
  INV_X1    g125(.A(G176gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT26), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n327), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(KEYINPUT26), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n324), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n322), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT65), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT23), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n333), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n344));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n332), .B1(KEYINPUT23), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n339), .B2(new_n341), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT23), .ZN(new_n349));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT66), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n353));
  MUX2_X1   g152(.A(G183gat), .B(new_n353), .S(G190gat), .Z(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(KEYINPUT24), .B2(new_n324), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n328), .A2(KEYINPUT23), .A3(new_n330), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n350), .A2(KEYINPUT25), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n359), .A2(new_n348), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT24), .B1(new_n323), .B2(KEYINPUT68), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(KEYINPUT68), .B2(new_n323), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n354), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n337), .B1(new_n358), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n311), .B1(new_n366), .B2(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT77), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT22), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n369), .A2(KEYINPUT75), .B1(G211gat), .B2(G218gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(KEYINPUT75), .B2(new_n369), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n373));
  XNOR2_X1  g172(.A(G197gat), .B(G204gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G211gat), .B(G218gat), .Z(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n376), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n372), .A2(new_n378), .A3(new_n373), .A4(new_n374), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n358), .A2(new_n365), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT69), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n322), .A2(new_n335), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n322), .B2(new_n335), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n311), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n356), .A2(new_n357), .B1(new_n364), .B2(new_n361), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n337), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n311), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n368), .A2(new_n380), .A3(new_n388), .A4(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n386), .A2(new_n389), .A3(new_n311), .ZN(new_n395));
  INV_X1    g194(.A(new_n380), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n366), .A2(new_n387), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(G8gat), .B(G36gat), .Z(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT78), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n394), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n393), .A2(new_n388), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n392), .B1(new_n391), .B2(new_n311), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n407), .A2(new_n396), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n398), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n402), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n394), .A2(KEYINPUT30), .A3(new_n398), .A4(new_n403), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n406), .A2(new_n411), .A3(KEYINPUT79), .A4(new_n412), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n412), .A2(KEYINPUT79), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n306), .A2(new_n308), .A3(new_n297), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT40), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n310), .A2(new_n413), .A3(new_n414), .A4(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n377), .B2(new_n379), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n258), .B1(new_n419), .B2(KEYINPUT3), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n262), .A2(new_n389), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n396), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n424), .B1(new_n420), .B2(new_n422), .ZN(new_n427));
  NAND2_X1  g226(.A1(G228gat), .A2(G233gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(G22gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OR3_X1    g231(.A1(new_n426), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n432), .B1(new_n426), .B2(new_n427), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n293), .A2(KEYINPUT6), .A3(new_n298), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n293), .B2(new_n298), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT85), .B1(new_n281), .B2(KEYINPUT5), .ZN(new_n439));
  AOI211_X1 g238(.A(new_n268), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n289), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n291), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n283), .A2(KEYINPUT86), .A3(new_n289), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n266), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n297), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n436), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n394), .A2(new_n447), .A3(new_n398), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n402), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n394), .B2(new_n398), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT38), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n395), .A2(new_n397), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n447), .B1(new_n452), .B2(new_n380), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n368), .A2(new_n388), .A3(new_n393), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n380), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT38), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n451), .B(new_n404), .C1(new_n449), .C2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n418), .B(new_n435), .C1(new_n446), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT74), .ZN(new_n460));
  XNOR2_X1  g259(.A(G15gat), .B(G43gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT64), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n336), .A2(KEYINPUT69), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n322), .A2(new_n335), .A3(new_n382), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n468), .A2(new_n390), .A3(new_n260), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n244), .B1(new_n381), .B2(new_n385), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n463), .B1(new_n471), .B2(KEYINPUT32), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n465), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n260), .B1(new_n468), .B2(new_n390), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n381), .A2(new_n385), .A3(new_n244), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT32), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n463), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n481), .A2(KEYINPUT71), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(KEYINPUT71), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(KEYINPUT33), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n472), .A2(new_n474), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n476), .A2(new_n477), .A3(new_n475), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT73), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n471), .A2(KEYINPUT32), .A3(new_n484), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n481), .B1(new_n478), .B2(new_n479), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n478), .A2(KEYINPUT33), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT73), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n486), .B(KEYINPUT34), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n460), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n493), .A2(new_n495), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n472), .A2(new_n474), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n501), .A2(KEYINPUT73), .A3(new_n488), .A4(new_n490), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT74), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n502), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n493), .A2(KEYINPUT72), .A3(new_n495), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT36), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n444), .B2(new_n297), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT6), .B1(new_n444), .B2(new_n297), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n293), .A2(KEYINPUT88), .A3(new_n298), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n436), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n413), .A2(new_n414), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n435), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n511), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n505), .A2(new_n435), .A3(new_n507), .A4(new_n508), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n518), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n497), .A2(new_n499), .A3(new_n503), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT89), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n497), .A2(new_n528), .A3(new_n499), .A4(new_n503), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n518), .A2(new_n530), .A3(new_n435), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n527), .A2(new_n529), .A3(new_n446), .A4(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n459), .A2(new_n521), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT16), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(G1gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n536), .B(new_n537), .C1(G1gat), .C2(new_n534), .ZN(new_n538));
  OR2_X1    g337(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G29gat), .ZN(new_n541));
  INV_X1    g340(.A(G36gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT14), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT14), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n546), .A2(new_n547), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n547), .B2(new_n546), .ZN(new_n549));
  XOR2_X1   g348(.A(G43gat), .B(G50gat), .Z(new_n550));
  INV_X1    g349(.A(KEYINPUT15), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n546), .B1(new_n551), .B2(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(G29gat), .A2(G36gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT92), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n554), .B(new_n556), .C1(new_n551), .C2(new_n550), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT94), .ZN(new_n560));
  NAND2_X1  g359(.A1(G229gat), .A2(G233gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n540), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n553), .A2(KEYINPUT17), .A3(new_n557), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n560), .A2(KEYINPUT18), .A3(new_n561), .A4(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n559), .A2(KEYINPUT94), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n540), .B2(new_n558), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n561), .B(new_n566), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n540), .A2(new_n558), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n568), .B2(new_n570), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n561), .B(KEYINPUT13), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n567), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G169gat), .B(G197gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT12), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n567), .A2(new_n573), .A3(new_n577), .A4(new_n584), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n202), .B1(new_n533), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n413), .A2(new_n414), .ZN(new_n591));
  AOI211_X1 g390(.A(new_n591), .B(new_n522), .C1(new_n516), .C2(new_n436), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n532), .B1(new_n592), .B2(new_n530), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n504), .A2(new_n510), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n516), .B2(new_n436), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n459), .B(new_n594), .C1(new_n595), .C2(new_n435), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(KEYINPUT95), .A3(new_n588), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n517), .ZN(new_n600));
  XNOR2_X1  g399(.A(G57gat), .B(G64gat), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G71gat), .B(G78gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G127gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n564), .B1(new_n607), .B2(new_n606), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n204), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n613), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT7), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G99gat), .B(G106gat), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n621), .B(new_n625), .C1(KEYINPUT96), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(KEYINPUT96), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n563), .A2(new_n565), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n627), .B(new_n628), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n558), .ZN(new_n632));
  NAND3_X1  g431(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT97), .B1(new_n632), .B2(new_n633), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n630), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT98), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n639), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n630), .B(new_n645), .C1(new_n636), .C2(new_n637), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n640), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n640), .B2(new_n646), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n619), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n606), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n626), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n627), .B1(KEYINPUT96), .B2(new_n626), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n605), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n631), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G230gat), .ZN(new_n660));
  INV_X1    g459(.A(G233gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n652), .A2(new_n655), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n665), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n664), .B(new_n669), .C1(new_n665), .C2(new_n663), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT99), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n666), .A2(new_n674), .A3(new_n670), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n651), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n599), .A2(new_n600), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n591), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n590), .B2(new_n598), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT16), .B(G8gat), .Z(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n683), .A2(KEYINPUT100), .A3(KEYINPUT42), .A4(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(G8gat), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT42), .B1(new_n683), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n685), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(G1325gat));
  AND2_X1   g492(.A1(new_n599), .A2(new_n678), .ZN(new_n694));
  INV_X1    g493(.A(G15gat), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n527), .A2(new_n529), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n511), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n699), .B2(new_n695), .ZN(G1326gat));
  NAND3_X1  g499(.A1(new_n599), .A2(new_n520), .A3(new_n678), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT43), .B(G22gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  INV_X1    g502(.A(new_n619), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n676), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n650), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n599), .A2(new_n541), .A3(new_n600), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n533), .B2(new_n650), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n597), .A2(KEYINPUT44), .A3(new_n649), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n705), .A2(new_n589), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(new_n600), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n709), .B(new_n710), .C1(new_n541), .C2(new_n716), .ZN(G1328gat));
  NAND4_X1  g516(.A1(new_n599), .A2(new_n542), .A3(new_n591), .A4(new_n706), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n715), .A2(new_n591), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n719), .B(new_n720), .C1(new_n542), .C2(new_n721), .ZN(G1329gat));
  NAND4_X1  g521(.A1(new_n712), .A2(new_n511), .A3(new_n713), .A4(new_n714), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT44), .B1(new_n597), .B2(new_n649), .ZN(new_n725));
  AOI211_X1 g524(.A(new_n711), .B(new_n650), .C1(new_n593), .C2(new_n596), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n727), .A2(new_n728), .A3(new_n511), .A4(new_n714), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n724), .A2(new_n729), .A3(G43gat), .ZN(new_n730));
  INV_X1    g529(.A(new_n696), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(G43gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n599), .A2(new_n706), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(KEYINPUT47), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n735));
  AND2_X1   g534(.A1(new_n723), .A2(G43gat), .ZN(new_n736));
  INV_X1    g535(.A(new_n733), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(G1330gat));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740));
  INV_X1    g539(.A(G50gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n715), .B2(new_n520), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n435), .A2(G50gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n599), .A2(new_n706), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n740), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n727), .A2(new_n520), .A3(new_n714), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G50gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(KEYINPUT48), .A3(new_n744), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(G1331gat));
  NOR3_X1   g549(.A1(new_n651), .A2(new_n588), .A3(new_n676), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n597), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n600), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n597), .A2(new_n751), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT104), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n518), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n760), .B2(new_n761), .ZN(G1333gat));
  XNOR2_X1  g563(.A(new_n696), .B(KEYINPUT105), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n757), .A2(G71gat), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n756), .A2(new_n511), .A3(new_n758), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(G71gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g568(.A1(new_n759), .A2(new_n435), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g570(.A1(new_n619), .A2(new_n588), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n597), .A2(new_n649), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n597), .A2(KEYINPUT51), .A3(new_n649), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n676), .A2(G85gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n600), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n772), .A2(new_n677), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n725), .A2(new_n726), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n623), .B1(new_n782), .B2(new_n600), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT106), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT106), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n782), .A2(new_n600), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n785), .B(new_n779), .C1(new_n786), .C2(new_n623), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1336gat));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n518), .A2(G92gat), .A3(new_n676), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n777), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n782), .A2(new_n591), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n789), .B(new_n791), .C1(new_n792), .C2(new_n624), .ZN(new_n793));
  INV_X1    g592(.A(new_n791), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n624), .B1(new_n782), .B2(new_n591), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT52), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(G1337gat));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n511), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G99gat), .ZN(new_n799));
  INV_X1    g598(.A(new_n777), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n731), .A2(G99gat), .A3(new_n676), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(G1338gat));
  INV_X1    g601(.A(G106gat), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n782), .B2(new_n520), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n676), .A2(new_n435), .A3(G106gat), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT107), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n775), .B2(new_n776), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT53), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(KEYINPUT108), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n811));
  AOI211_X1 g610(.A(new_n811), .B(new_n806), .C1(new_n775), .C2(new_n776), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n781), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n712), .A2(new_n520), .A3(new_n713), .A4(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n727), .A2(KEYINPUT109), .A3(new_n520), .A4(new_n814), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n817), .A2(new_n818), .A3(G106gat), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n808), .B1(new_n813), .B2(new_n819), .ZN(G1339gat));
  NOR2_X1   g619(.A1(new_n517), .A2(new_n591), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n664), .A2(new_n823), .A3(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n662), .B1(new_n657), .B2(new_n658), .ZN(new_n825));
  XOR2_X1   g624(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n826));
  AOI21_X1  g625(.A(new_n669), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n672), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(KEYINPUT111), .A3(new_n672), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n664), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n834));
  INV_X1    g633(.A(new_n826), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n670), .B1(new_n664), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n831), .A2(new_n588), .A3(new_n832), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT112), .B1(new_n575), .B2(new_n576), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n560), .A2(new_n566), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n561), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n575), .A2(KEYINPUT112), .A3(new_n576), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n583), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(new_n587), .A3(new_n675), .A4(new_n673), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n649), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n843), .B(new_n587), .C1(new_n647), .C2(new_n648), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n832), .A3(new_n837), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n704), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n619), .A2(new_n589), .A3(new_n650), .A4(new_n676), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n822), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n523), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(KEYINPUT114), .Z(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n230), .A3(new_n588), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n850), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n435), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT113), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n731), .A2(new_n822), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n588), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n854), .B1(new_n860), .B2(new_n230), .ZN(G1340gat));
  NAND3_X1  g660(.A1(new_n853), .A2(new_n228), .A3(new_n677), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(new_n858), .ZN(new_n863));
  OAI21_X1  g662(.A(G120gat), .B1(new_n863), .B2(new_n676), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n863), .B2(new_n704), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n619), .A2(new_n236), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n852), .B2(new_n867), .ZN(G1342gat));
  OAI21_X1  g667(.A(G134gat), .B1(new_n863), .B2(new_n650), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n851), .A2(new_n238), .A3(new_n523), .A4(new_n649), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT56), .Z(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n869), .A2(new_n871), .A3(KEYINPUT115), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n822), .A2(new_n511), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n520), .A2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(new_n850), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n834), .B2(new_n836), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n824), .A2(KEYINPUT117), .A3(new_n827), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n833), .A3(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n829), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n588), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n649), .B1(new_n885), .B2(new_n844), .ZN(new_n886));
  OAI22_X1  g685(.A1(new_n886), .A2(KEYINPUT118), .B1(new_n847), .B2(new_n846), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(KEYINPUT118), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n704), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n879), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT119), .B(new_n704), .C1(new_n887), .C2(new_n888), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n878), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n435), .B1(new_n849), .B2(new_n850), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  XOR2_X1   g694(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n896));
  AND2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n588), .B(new_n877), .C1(new_n893), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G141gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n594), .A2(new_n520), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n851), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OR3_X1    g702(.A1(new_n903), .A2(G141gat), .A3(new_n589), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT58), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n899), .A2(new_n907), .A3(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1344gat));
  NOR3_X1   g708(.A1(new_n903), .A2(G148gat), .A3(new_n676), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n704), .B1(new_n886), .B2(new_n848), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n850), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n435), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(KEYINPUT122), .A3(new_n850), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT57), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n895), .A2(new_n896), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n677), .B(new_n877), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n212), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n911), .A2(new_n912), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n877), .B1(new_n893), .B2(new_n897), .ZN(new_n924));
  OAI21_X1  g723(.A(G148gat), .B1(new_n924), .B2(new_n676), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n921), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n926), .ZN(G1345gat));
  OAI21_X1  g726(.A(G155gat), .B1(new_n924), .B2(new_n704), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n619), .A2(new_n204), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n903), .B2(new_n929), .ZN(G1346gat));
  OAI211_X1 g729(.A(new_n649), .B(new_n877), .C1(new_n893), .C2(new_n897), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n205), .B1(new_n931), .B2(KEYINPUT123), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(KEYINPUT123), .B2(new_n931), .ZN(new_n933));
  OR3_X1    g732(.A1(new_n903), .A2(G162gat), .A3(new_n650), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n600), .A2(new_n518), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n855), .A2(new_n523), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n588), .ZN(new_n939));
  INV_X1    g738(.A(new_n936), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n765), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n857), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n589), .A2(new_n326), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(G1348gat));
  OAI21_X1  g744(.A(G176gat), .B1(new_n942), .B2(new_n676), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n938), .A2(new_n327), .A3(new_n677), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1349gat));
  OAI21_X1  g747(.A(G183gat), .B1(new_n942), .B2(new_n704), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n938), .A2(new_n320), .A3(new_n619), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT60), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1350gat));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n316), .A3(new_n649), .ZN(new_n956));
  OAI21_X1  g755(.A(G190gat), .B1(new_n942), .B2(new_n650), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  NOR2_X1   g759(.A1(new_n940), .A2(new_n511), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n894), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n588), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n918), .A2(new_n919), .ZN(new_n965));
  INV_X1    g764(.A(new_n961), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n588), .A2(G197gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1352gat));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n970));
  INV_X1    g769(.A(G204gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n971), .B1(new_n967), .B2(new_n677), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n961), .A2(new_n971), .A3(new_n677), .A4(new_n894), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n974), .A2(new_n975), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n977), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n970), .B1(new_n972), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n977), .B(new_n978), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n965), .A2(new_n676), .A3(new_n966), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n982), .B(KEYINPUT125), .C1(new_n971), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n981), .A2(new_n984), .ZN(G1353gat));
  OAI211_X1 g784(.A(new_n619), .B(new_n961), .C1(new_n918), .C2(new_n919), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT63), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n986), .A2(new_n987), .A3(G211gat), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n704), .A2(G211gat), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n961), .A2(new_n894), .A3(new_n989), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n987), .B1(new_n986), .B2(G211gat), .ZN(new_n994));
  OAI21_X1  g793(.A(KEYINPUT127), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n986), .A2(G211gat), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(KEYINPUT63), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  NAND4_X1  g797(.A1(new_n997), .A2(new_n998), .A3(new_n988), .A4(new_n992), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n995), .A2(new_n999), .ZN(G1354gat));
  INV_X1    g799(.A(G218gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n963), .A2(new_n1001), .A3(new_n649), .ZN(new_n1002));
  NOR3_X1   g801(.A1(new_n965), .A2(new_n650), .A3(new_n966), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1002), .B1(new_n1003), .B2(new_n1001), .ZN(G1355gat));
endmodule


