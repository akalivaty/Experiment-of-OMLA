

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U558 ( .A1(G301), .A2(n743), .ZN(n526) );
  XOR2_X1 U559 ( .A(n750), .B(KEYINPUT31), .Z(n527) );
  NOR2_X1 U560 ( .A1(n758), .A2(n924), .ZN(n716) );
  NAND2_X1 U561 ( .A1(n751), .A2(n527), .ZN(n757) );
  NOR2_X1 U562 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U563 ( .A1(n711), .A2(n710), .ZN(n758) );
  NOR2_X1 U564 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n532), .ZN(n892) );
  NOR2_X1 U566 ( .A1(G651), .A2(n633), .ZN(n664) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n528), .Z(n887) );
  NAND2_X1 U569 ( .A1(G138), .A2(n887), .ZN(n536) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U571 ( .A1(G114), .A2(n891), .ZN(n529) );
  XOR2_X1 U572 ( .A(KEYINPUT83), .B(n529), .Z(n531) );
  INV_X1 U573 ( .A(G2105), .ZN(n532) );
  NAND2_X1 U574 ( .A1(n892), .A2(G126), .ZN(n530) );
  NAND2_X1 U575 ( .A1(n531), .A2(n530), .ZN(n534) );
  AND2_X1 U576 ( .A1(n532), .A2(G2104), .ZN(n888) );
  AND2_X1 U577 ( .A1(G102), .A2(n888), .ZN(n533) );
  NOR2_X1 U578 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U579 ( .A1(n536), .A2(n535), .ZN(n538) );
  INV_X1 U580 ( .A(KEYINPUT84), .ZN(n537) );
  XNOR2_X1 U581 ( .A(n538), .B(n537), .ZN(n691) );
  BUF_X1 U582 ( .A(n691), .Z(G164) );
  XNOR2_X1 U583 ( .A(G2451), .B(G2446), .ZN(n548) );
  XOR2_X1 U584 ( .A(G2430), .B(KEYINPUT105), .Z(n540) );
  XNOR2_X1 U585 ( .A(G2454), .B(G2435), .ZN(n539) );
  XNOR2_X1 U586 ( .A(n540), .B(n539), .ZN(n544) );
  XOR2_X1 U587 ( .A(G2438), .B(KEYINPUT104), .Z(n542) );
  XNOR2_X1 U588 ( .A(G1341), .B(G1348), .ZN(n541) );
  XNOR2_X1 U589 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U590 ( .A(n544), .B(n543), .Z(n546) );
  XNOR2_X1 U591 ( .A(G2443), .B(G2427), .ZN(n545) );
  XNOR2_X1 U592 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U593 ( .A(n548), .B(n547), .ZN(n549) );
  AND2_X1 U594 ( .A1(n549), .A2(G14), .ZN(G401) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U596 ( .A1(G135), .A2(n887), .ZN(n550) );
  XNOR2_X1 U597 ( .A(n550), .B(KEYINPUT72), .ZN(n557) );
  NAND2_X1 U598 ( .A1(G111), .A2(n891), .ZN(n552) );
  NAND2_X1 U599 ( .A1(G99), .A2(n888), .ZN(n551) );
  NAND2_X1 U600 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U601 ( .A1(n892), .A2(G123), .ZN(n553) );
  XOR2_X1 U602 ( .A(KEYINPUT18), .B(n553), .Z(n554) );
  NOR2_X1 U603 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U604 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U605 ( .A(KEYINPUT73), .B(n558), .Z(n1011) );
  XNOR2_X1 U606 ( .A(G2096), .B(n1011), .ZN(n559) );
  OR2_X1 U607 ( .A1(G2100), .A2(n559), .ZN(G156) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G651), .ZN(n564) );
  NOR2_X1 U610 ( .A1(G543), .A2(n564), .ZN(n560) );
  XOR2_X1 U611 ( .A(KEYINPUT1), .B(n560), .Z(n663) );
  NAND2_X1 U612 ( .A1(G65), .A2(n663), .ZN(n563) );
  XOR2_X1 U613 ( .A(G543), .B(KEYINPUT0), .Z(n561) );
  XNOR2_X1 U614 ( .A(KEYINPUT64), .B(n561), .ZN(n633) );
  NAND2_X1 U615 ( .A1(G53), .A2(n664), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n563), .A2(n562), .ZN(n568) );
  NOR2_X1 U617 ( .A1(G543), .A2(G651), .ZN(n659) );
  NAND2_X1 U618 ( .A1(G91), .A2(n659), .ZN(n566) );
  NOR2_X1 U619 ( .A1(n633), .A2(n564), .ZN(n660) );
  NAND2_X1 U620 ( .A1(G78), .A2(n660), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U622 ( .A1(n568), .A2(n567), .ZN(n731) );
  INV_X1 U623 ( .A(n731), .ZN(G299) );
  NAND2_X1 U624 ( .A1(G88), .A2(n659), .ZN(n569) );
  XNOR2_X1 U625 ( .A(n569), .B(KEYINPUT78), .ZN(n571) );
  NAND2_X1 U626 ( .A1(n663), .A2(G62), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U628 ( .A1(G75), .A2(n660), .ZN(n573) );
  NAND2_X1 U629 ( .A1(G50), .A2(n664), .ZN(n572) );
  NAND2_X1 U630 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U631 ( .A1(n575), .A2(n574), .ZN(G166) );
  NAND2_X1 U632 ( .A1(G64), .A2(n663), .ZN(n577) );
  NAND2_X1 U633 ( .A1(G52), .A2(n664), .ZN(n576) );
  NAND2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n582) );
  NAND2_X1 U635 ( .A1(G90), .A2(n659), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G77), .A2(n660), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U638 ( .A(KEYINPUT9), .B(n580), .Z(n581) );
  NOR2_X1 U639 ( .A1(n582), .A2(n581), .ZN(G171) );
  NAND2_X1 U640 ( .A1(n887), .A2(G137), .ZN(n585) );
  NAND2_X1 U641 ( .A1(G101), .A2(n888), .ZN(n583) );
  XOR2_X1 U642 ( .A(KEYINPUT23), .B(n583), .Z(n584) );
  NAND2_X1 U643 ( .A1(n585), .A2(n584), .ZN(n694) );
  NAND2_X1 U644 ( .A1(G113), .A2(n891), .ZN(n587) );
  NAND2_X1 U645 ( .A1(G125), .A2(n892), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(n692) );
  NOR2_X1 U647 ( .A1(n694), .A2(n692), .ZN(G160) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n588) );
  XNOR2_X1 U649 ( .A(n588), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U650 ( .A(G223), .ZN(n833) );
  NAND2_X1 U651 ( .A1(n833), .A2(G567), .ZN(n589) );
  XOR2_X1 U652 ( .A(KEYINPUT11), .B(n589), .Z(G234) );
  NAND2_X1 U653 ( .A1(G56), .A2(n663), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n590), .Z(n596) );
  NAND2_X1 U655 ( .A1(n659), .A2(G81), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n591), .B(KEYINPUT12), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G68), .A2(n660), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(n594), .Z(n595) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U661 ( .A1(n664), .A2(G43), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n942) );
  INV_X1 U663 ( .A(G860), .ZN(n841) );
  OR2_X1 U664 ( .A1(n942), .A2(n841), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n608) );
  NAND2_X1 U667 ( .A1(G54), .A2(n664), .ZN(n605) );
  NAND2_X1 U668 ( .A1(G66), .A2(n663), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G79), .A2(n660), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U671 ( .A1(G92), .A2(n659), .ZN(n601) );
  XNOR2_X1 U672 ( .A(KEYINPUT65), .B(n601), .ZN(n602) );
  NOR2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n606), .B(KEYINPUT15), .ZN(n908) );
  INV_X1 U676 ( .A(n908), .ZN(n960) );
  INV_X1 U677 ( .A(G868), .ZN(n674) );
  NAND2_X1 U678 ( .A1(n960), .A2(n674), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(G284) );
  NAND2_X1 U680 ( .A1(G63), .A2(n663), .ZN(n610) );
  NAND2_X1 U681 ( .A1(G51), .A2(n664), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U683 ( .A(KEYINPUT6), .B(n611), .ZN(n619) );
  NAND2_X1 U684 ( .A1(G89), .A2(n659), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n612), .B(KEYINPUT66), .ZN(n613) );
  XNOR2_X1 U686 ( .A(KEYINPUT4), .B(n613), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n660), .A2(G76), .ZN(n614) );
  XOR2_X1 U688 ( .A(KEYINPUT67), .B(n614), .Z(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U690 ( .A(n617), .B(KEYINPUT5), .Z(n618) );
  NOR2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U692 ( .A(KEYINPUT7), .B(n620), .Z(n621) );
  XNOR2_X1 U693 ( .A(KEYINPUT68), .B(n621), .ZN(G168) );
  XOR2_X1 U694 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U695 ( .A1(G286), .A2(n674), .ZN(n622) );
  XOR2_X1 U696 ( .A(KEYINPUT69), .B(n622), .Z(n624) );
  NOR2_X1 U697 ( .A1(G868), .A2(G299), .ZN(n623) );
  NOR2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U699 ( .A(KEYINPUT70), .B(n625), .ZN(G297) );
  NAND2_X1 U700 ( .A1(n841), .A2(G559), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n626), .A2(n908), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT16), .ZN(n628) );
  XOR2_X1 U703 ( .A(KEYINPUT71), .B(n628), .Z(G148) );
  NOR2_X1 U704 ( .A1(G868), .A2(n942), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G868), .A2(n908), .ZN(n629) );
  NOR2_X1 U706 ( .A1(G559), .A2(n629), .ZN(n630) );
  NOR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT76), .ZN(n638) );
  NAND2_X1 U710 ( .A1(G49), .A2(n664), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G87), .A2(n633), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U713 ( .A1(n663), .A2(n636), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(G288) );
  AND2_X1 U715 ( .A1(n663), .A2(G60), .ZN(n642) );
  NAND2_X1 U716 ( .A1(G85), .A2(n659), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G72), .A2(n660), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n664), .A2(G47), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(G290) );
  NAND2_X1 U722 ( .A1(G73), .A2(n660), .ZN(n645) );
  XNOR2_X1 U723 ( .A(n645), .B(KEYINPUT2), .ZN(n652) );
  NAND2_X1 U724 ( .A1(G61), .A2(n663), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G86), .A2(n659), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U727 ( .A1(G48), .A2(n664), .ZN(n648) );
  XNOR2_X1 U728 ( .A(KEYINPUT77), .B(n648), .ZN(n649) );
  NOR2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(G305) );
  NAND2_X1 U731 ( .A1(G559), .A2(n908), .ZN(n653) );
  XOR2_X1 U732 ( .A(n942), .B(n653), .Z(n840) );
  XNOR2_X1 U733 ( .A(n840), .B(KEYINPUT80), .ZN(n672) );
  XOR2_X1 U734 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n654) );
  XNOR2_X1 U735 ( .A(G288), .B(n654), .ZN(n655) );
  XNOR2_X1 U736 ( .A(n731), .B(n655), .ZN(n657) );
  XNOR2_X1 U737 ( .A(G290), .B(G166), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n658), .B(G305), .ZN(n671) );
  NAND2_X1 U740 ( .A1(G93), .A2(n659), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G80), .A2(n660), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n669) );
  NAND2_X1 U743 ( .A1(G67), .A2(n663), .ZN(n666) );
  NAND2_X1 U744 ( .A1(G55), .A2(n664), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U746 ( .A(KEYINPUT74), .B(n667), .ZN(n668) );
  NOR2_X1 U747 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n670), .B(KEYINPUT75), .ZN(n842) );
  XNOR2_X1 U749 ( .A(n671), .B(n842), .ZN(n911) );
  XNOR2_X1 U750 ( .A(n672), .B(n911), .ZN(n673) );
  NAND2_X1 U751 ( .A1(n673), .A2(G868), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n674), .A2(n842), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2084), .A2(G2078), .ZN(n677) );
  XNOR2_X1 U755 ( .A(n677), .B(KEYINPUT81), .ZN(n678) );
  XNOR2_X1 U756 ( .A(KEYINPUT20), .B(n678), .ZN(n679) );
  NAND2_X1 U757 ( .A1(n679), .A2(G2090), .ZN(n680) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U759 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U761 ( .A1(G132), .A2(G82), .ZN(n682) );
  XNOR2_X1 U762 ( .A(n682), .B(KEYINPUT82), .ZN(n683) );
  XNOR2_X1 U763 ( .A(n683), .B(KEYINPUT22), .ZN(n684) );
  NOR2_X1 U764 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U765 ( .A1(G96), .A2(n685), .ZN(n838) );
  NAND2_X1 U766 ( .A1(n838), .A2(G2106), .ZN(n689) );
  NAND2_X1 U767 ( .A1(G69), .A2(G120), .ZN(n686) );
  NOR2_X1 U768 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U769 ( .A1(G108), .A2(n687), .ZN(n839) );
  NAND2_X1 U770 ( .A1(n839), .A2(G567), .ZN(n688) );
  NAND2_X1 U771 ( .A1(n689), .A2(n688), .ZN(n844) );
  NAND2_X1 U772 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U773 ( .A1(n844), .A2(n690), .ZN(n835) );
  NAND2_X1 U774 ( .A1(n835), .A2(G36), .ZN(G176) );
  INV_X1 U775 ( .A(G166), .ZN(G303) );
  NOR2_X1 U776 ( .A1(G1384), .A2(n691), .ZN(n711) );
  INV_X1 U777 ( .A(G40), .ZN(n693) );
  OR2_X1 U778 ( .A1(n693), .A2(n692), .ZN(n695) );
  OR2_X1 U779 ( .A1(n695), .A2(n694), .ZN(n709) );
  NOR2_X1 U780 ( .A1(n711), .A2(n709), .ZN(n827) );
  NAND2_X1 U781 ( .A1(n887), .A2(G140), .ZN(n696) );
  XNOR2_X1 U782 ( .A(n696), .B(KEYINPUT86), .ZN(n698) );
  NAND2_X1 U783 ( .A1(G104), .A2(n888), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n700) );
  XOR2_X1 U785 ( .A(KEYINPUT87), .B(KEYINPUT34), .Z(n699) );
  XNOR2_X1 U786 ( .A(n700), .B(n699), .ZN(n705) );
  NAND2_X1 U787 ( .A1(G116), .A2(n891), .ZN(n702) );
  NAND2_X1 U788 ( .A1(G128), .A2(n892), .ZN(n701) );
  NAND2_X1 U789 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U790 ( .A(KEYINPUT35), .B(n703), .Z(n704) );
  NOR2_X1 U791 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U792 ( .A(n706), .B(KEYINPUT36), .ZN(n707) );
  XNOR2_X1 U793 ( .A(n707), .B(KEYINPUT88), .ZN(n903) );
  XNOR2_X1 U794 ( .A(KEYINPUT37), .B(G2067), .ZN(n825) );
  NOR2_X1 U795 ( .A1(n903), .A2(n825), .ZN(n1023) );
  NAND2_X1 U796 ( .A1(n827), .A2(n1023), .ZN(n708) );
  XOR2_X1 U797 ( .A(KEYINPUT89), .B(n708), .Z(n823) );
  INV_X1 U798 ( .A(n823), .ZN(n814) );
  XNOR2_X1 U799 ( .A(n709), .B(KEYINPUT93), .ZN(n710) );
  NAND2_X1 U800 ( .A1(G8), .A2(n758), .ZN(n785) );
  NOR2_X1 U801 ( .A1(G2084), .A2(n758), .ZN(n744) );
  NAND2_X1 U802 ( .A1(n744), .A2(G8), .ZN(n756) );
  NOR2_X1 U803 ( .A1(G1966), .A2(n785), .ZN(n753) );
  INV_X1 U804 ( .A(n758), .ZN(n738) );
  NAND2_X1 U805 ( .A1(n738), .A2(G2072), .ZN(n712) );
  XNOR2_X1 U806 ( .A(n712), .B(KEYINPUT27), .ZN(n714) );
  INV_X1 U807 ( .A(G1956), .ZN(n970) );
  NOR2_X1 U808 ( .A1(n970), .A2(n738), .ZN(n713) );
  NOR2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n732) );
  NAND2_X1 U810 ( .A1(n732), .A2(n731), .ZN(n730) );
  INV_X1 U811 ( .A(G1996), .ZN(n924) );
  XNOR2_X1 U812 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n715) );
  XNOR2_X1 U813 ( .A(n716), .B(n715), .ZN(n718) );
  NAND2_X1 U814 ( .A1(n758), .A2(G1341), .ZN(n717) );
  NAND2_X1 U815 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X2 U816 ( .A1(n719), .A2(n942), .ZN(n720) );
  OR2_X1 U817 ( .A1(n908), .A2(n720), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n720), .A2(n908), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n758), .A2(G1348), .ZN(n721) );
  XNOR2_X1 U820 ( .A(n721), .B(KEYINPUT96), .ZN(n723) );
  NAND2_X1 U821 ( .A1(n738), .A2(G2067), .ZN(n722) );
  NAND2_X1 U822 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U823 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U824 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U825 ( .A(KEYINPUT97), .B(n728), .Z(n729) );
  NAND2_X1 U826 ( .A1(n730), .A2(n729), .ZN(n735) );
  NOR2_X1 U827 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U828 ( .A(n733), .B(KEYINPUT28), .Z(n734) );
  NAND2_X1 U829 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U830 ( .A(n736), .B(KEYINPUT29), .ZN(n737) );
  INV_X1 U831 ( .A(n737), .ZN(n742) );
  NOR2_X1 U832 ( .A1(n738), .A2(G1961), .ZN(n739) );
  XNOR2_X1 U833 ( .A(n739), .B(KEYINPUT94), .ZN(n741) );
  XOR2_X1 U834 ( .A(G2078), .B(KEYINPUT25), .Z(n930) );
  NOR2_X1 U835 ( .A1(n758), .A2(n930), .ZN(n740) );
  NOR2_X1 U836 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U837 ( .A1(n742), .A2(n526), .ZN(n751) );
  AND2_X1 U838 ( .A1(G301), .A2(n743), .ZN(n749) );
  NOR2_X1 U839 ( .A1(n753), .A2(n744), .ZN(n745) );
  NAND2_X1 U840 ( .A1(G8), .A2(n745), .ZN(n746) );
  XNOR2_X1 U841 ( .A(KEYINPUT30), .B(n746), .ZN(n747) );
  NOR2_X1 U842 ( .A1(n747), .A2(G168), .ZN(n748) );
  NOR2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n750) );
  INV_X1 U844 ( .A(n757), .ZN(n752) );
  XNOR2_X1 U845 ( .A(KEYINPUT98), .B(n754), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n769) );
  NAND2_X1 U847 ( .A1(n757), .A2(G286), .ZN(n764) );
  NOR2_X1 U848 ( .A1(G2090), .A2(n758), .ZN(n759) );
  XNOR2_X1 U849 ( .A(KEYINPUT99), .B(n759), .ZN(n762) );
  NOR2_X1 U850 ( .A1(G1971), .A2(n785), .ZN(n760) );
  NOR2_X1 U851 ( .A1(G166), .A2(n760), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n765), .A2(G8), .ZN(n767) );
  XNOR2_X1 U855 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n766) );
  XNOR2_X1 U856 ( .A(n767), .B(n766), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n784) );
  NOR2_X1 U858 ( .A1(G1971), .A2(G303), .ZN(n770) );
  NOR2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n949) );
  NOR2_X1 U860 ( .A1(n770), .A2(n949), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n784), .A2(n771), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G1976), .A2(G288), .ZN(n951) );
  NAND2_X1 U863 ( .A1(n772), .A2(n951), .ZN(n773) );
  NOR2_X1 U864 ( .A1(n785), .A2(n773), .ZN(n774) );
  NOR2_X1 U865 ( .A1(KEYINPUT33), .A2(n774), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n949), .A2(KEYINPUT33), .ZN(n775) );
  NOR2_X1 U867 ( .A1(n775), .A2(n785), .ZN(n776) );
  XOR2_X1 U868 ( .A(G1981), .B(G305), .Z(n943) );
  NAND2_X1 U869 ( .A1(n778), .A2(n943), .ZN(n792) );
  NOR2_X1 U870 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XOR2_X1 U871 ( .A(n779), .B(KEYINPUT24), .Z(n780) );
  NOR2_X1 U872 ( .A1(n785), .A2(n780), .ZN(n790) );
  NOR2_X1 U873 ( .A1(G2090), .A2(G303), .ZN(n781) );
  XOR2_X1 U874 ( .A(KEYINPUT101), .B(n781), .Z(n782) );
  NAND2_X1 U875 ( .A1(G8), .A2(n782), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U878 ( .A(KEYINPUT102), .B(n787), .ZN(n788) );
  INV_X1 U879 ( .A(n788), .ZN(n789) );
  NOR2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n812) );
  NAND2_X1 U882 ( .A1(G95), .A2(n888), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G119), .A2(n892), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n887), .A2(G131), .ZN(n795) );
  XOR2_X1 U886 ( .A(KEYINPUT90), .B(n795), .Z(n796) );
  NOR2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n891), .A2(G107), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n880) );
  NAND2_X1 U890 ( .A1(G1991), .A2(n880), .ZN(n809) );
  NAND2_X1 U891 ( .A1(G105), .A2(n888), .ZN(n800) );
  XOR2_X1 U892 ( .A(KEYINPUT38), .B(n800), .Z(n805) );
  NAND2_X1 U893 ( .A1(G117), .A2(n891), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G129), .A2(n892), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U896 ( .A(KEYINPUT91), .B(n803), .Z(n804) );
  NOR2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U898 ( .A1(n887), .A2(G141), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n881) );
  NAND2_X1 U900 ( .A1(G1996), .A2(n881), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n1010) );
  NAND2_X1 U902 ( .A1(n1010), .A2(n827), .ZN(n810) );
  XOR2_X1 U903 ( .A(KEYINPUT92), .B(n810), .Z(n820) );
  INV_X1 U904 ( .A(n820), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n817) );
  XOR2_X1 U907 ( .A(G1986), .B(KEYINPUT85), .Z(n815) );
  XNOR2_X1 U908 ( .A(G290), .B(n815), .ZN(n954) );
  NAND2_X1 U909 ( .A1(n954), .A2(n827), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n830) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n881), .ZN(n1004) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n880), .ZN(n1002) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U914 ( .A1(n1002), .A2(n818), .ZN(n819) );
  NOR2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n1004), .A2(n821), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n903), .A2(n825), .ZN(n1020) );
  NAND2_X1 U920 ( .A1(n826), .A2(n1020), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n832) );
  XOR2_X1 U923 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n831) );
  XNOR2_X1 U924 ( .A(n832), .B(n831), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U927 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G1), .A2(G3), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U930 ( .A(n837), .B(KEYINPUT106), .ZN(G188) );
  INV_X1 U932 ( .A(G132), .ZN(G219) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G82), .ZN(G220) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  NAND2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(G145) );
  INV_X1 U940 ( .A(n844), .ZN(G319) );
  XOR2_X1 U941 ( .A(KEYINPUT109), .B(G1966), .Z(n846) );
  XNOR2_X1 U942 ( .A(G1981), .B(G1961), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U944 ( .A(n847), .B(KEYINPUT41), .Z(n849) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U947 ( .A(G1956), .B(G1971), .Z(n851) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1976), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U950 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U951 ( .A(KEYINPUT108), .B(G2474), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U953 ( .A(G2678), .B(G2084), .Z(n857) );
  XNOR2_X1 U954 ( .A(G2090), .B(G2078), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U956 ( .A(n858), .B(G2100), .Z(n860) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U959 ( .A(G2096), .B(KEYINPUT107), .Z(n862) );
  XNOR2_X1 U960 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n864), .B(n863), .Z(G227) );
  NAND2_X1 U963 ( .A1(G124), .A2(n892), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n891), .A2(G112), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G136), .A2(n887), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G100), .A2(n888), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U970 ( .A1(n871), .A2(n870), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G118), .A2(n891), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G130), .A2(n892), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G142), .A2(n887), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G106), .A2(n888), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(KEYINPUT110), .B(n876), .Z(n877) );
  XNOR2_X1 U978 ( .A(KEYINPUT45), .B(n877), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n902) );
  XOR2_X1 U980 ( .A(n881), .B(n880), .Z(n882) );
  XNOR2_X1 U981 ( .A(n1011), .B(n882), .ZN(n886) );
  XOR2_X1 U982 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n884) );
  XNOR2_X1 U983 ( .A(G162), .B(KEYINPUT46), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U985 ( .A(n886), .B(n885), .Z(n900) );
  NAND2_X1 U986 ( .A1(G139), .A2(n887), .ZN(n890) );
  NAND2_X1 U987 ( .A1(G103), .A2(n888), .ZN(n889) );
  NAND2_X1 U988 ( .A1(n890), .A2(n889), .ZN(n898) );
  NAND2_X1 U989 ( .A1(G115), .A2(n891), .ZN(n894) );
  NAND2_X1 U990 ( .A1(G127), .A2(n892), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U992 ( .A(KEYINPUT47), .B(n895), .ZN(n896) );
  XNOR2_X1 U993 ( .A(KEYINPUT111), .B(n896), .ZN(n897) );
  NOR2_X1 U994 ( .A1(n898), .A2(n897), .ZN(n1013) );
  XNOR2_X1 U995 ( .A(G160), .B(n1013), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n905) );
  XNOR2_X1 U998 ( .A(G164), .B(n903), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(n907) );
  XOR2_X1 U1001 ( .A(KEYINPUT113), .B(n907), .Z(G395) );
  XNOR2_X1 U1002 ( .A(n942), .B(KEYINPUT114), .ZN(n910) );
  XNOR2_X1 U1003 ( .A(G171), .B(n908), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n913) );
  XNOR2_X1 U1005 ( .A(G286), .B(n911), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(KEYINPUT49), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n916), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n917), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(KEYINPUT115), .B(n918), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G96), .ZN(G221) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1018 ( .A(G1991), .B(G25), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(G33), .B(G2072), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n929) );
  XOR2_X1 U1021 ( .A(G2067), .B(G26), .Z(n923) );
  NAND2_X1 U1022 ( .A1(n923), .A2(G28), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT120), .B(n924), .Z(n925) );
  XNOR2_X1 U1024 ( .A(G32), .B(n925), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n932) );
  XNOR2_X1 U1027 ( .A(G27), .B(n930), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1029 ( .A(KEYINPUT53), .B(n933), .Z(n936) );
  XOR2_X1 U1030 ( .A(KEYINPUT54), .B(G34), .Z(n934) );
  XNOR2_X1 U1031 ( .A(G2084), .B(n934), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1033 ( .A(KEYINPUT119), .B(G2090), .Z(n937) );
  XNOR2_X1 U1034 ( .A(G35), .B(n937), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1036 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n1025) );
  XNOR2_X1 U1037 ( .A(n940), .B(n1025), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(G29), .A2(n941), .ZN(n998) );
  XNOR2_X1 U1039 ( .A(G16), .B(KEYINPUT56), .ZN(n969) );
  XNOR2_X1 U1040 ( .A(n942), .B(G1341), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G168), .B(G1966), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n945), .B(KEYINPUT57), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(KEYINPUT121), .B(n946), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n967) );
  INV_X1 U1046 ( .A(n949), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1048 ( .A(KEYINPUT123), .B(n952), .Z(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n958) );
  XOR2_X1 U1050 ( .A(G1971), .B(G166), .Z(n956) );
  XNOR2_X1 U1051 ( .A(G299), .B(G1956), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(KEYINPUT124), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(G301), .B(G1961), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n960), .B(G1348), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1058 ( .A(KEYINPUT122), .B(n963), .Z(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n996) );
  INV_X1 U1062 ( .A(G16), .ZN(n994) );
  XOR2_X1 U1063 ( .A(G1966), .B(G21), .Z(n980) );
  XNOR2_X1 U1064 ( .A(G20), .B(n970), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(G1981), .B(G6), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G1341), .B(G19), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT59), .B(G1348), .Z(n975) );
  XNOR2_X1 U1070 ( .A(G4), .B(n975), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n978), .B(KEYINPUT60), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n981), .B(KEYINPUT125), .ZN(n989) );
  XOR2_X1 U1075 ( .A(G1986), .B(KEYINPUT126), .Z(n982) );
  XNOR2_X1 U1076 ( .A(G24), .B(n982), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G1976), .B(G23), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G22), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1081 ( .A(KEYINPUT58), .B(n987), .Z(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(G5), .B(G1961), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(KEYINPUT61), .B(n992), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(G11), .A2(n999), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(n1000), .B(KEYINPUT127), .ZN(n1029) );
  XOR2_X1 U1091 ( .A(G160), .B(G2084), .Z(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1008) );
  XOR2_X1 U1093 ( .A(G2090), .B(G162), .Z(n1003) );
  XNOR2_X1 U1094 ( .A(KEYINPUT116), .B(n1003), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(KEYINPUT51), .B(n1006), .Z(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1100 ( .A(G2072), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G164), .B(G2078), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT50), .B(n1016), .Z(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT117), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1024), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(G29), .ZN(n1028) );
  NAND2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

