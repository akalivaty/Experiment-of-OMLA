//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1216, new_n1217, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285, new_n1286;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(KEYINPUT64), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT64), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n214), .A2(G1), .A3(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AND2_X1   g0016(.A1(KEYINPUT65), .A2(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(KEYINPUT65), .A2(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(G50), .B1(G58), .B2(G68), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n211), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT66), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n229), .A2(KEYINPUT66), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n208), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  OR2_X1    g0036(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n223), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G226), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n226), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n228), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT69), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G107), .ZN(new_n252));
  INV_X1    g0052(.A(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G68), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G50), .B(G58), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n254), .B(new_n257), .Z(G351));
  INV_X1    g0058(.A(KEYINPUT10), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G150), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n219), .A2(G33), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n261), .B1(new_n206), .B2(new_n201), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n207), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n216), .ZN(new_n266));
  INV_X1    g0066(.A(G50), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n264), .A2(new_n266), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n265), .A2(new_n216), .A3(new_n270), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n205), .A2(G20), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G50), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT9), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G274), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n280), .A2(new_n282), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(G226), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(KEYINPUT70), .A2(G223), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT70), .A2(G223), .ZN(new_n287));
  OAI21_X1  g0087(.A(G1698), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G222), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n213), .A2(new_n215), .A3(new_n279), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n292), .B(new_n294), .C1(G77), .C2(new_n289), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n285), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G190), .B2(new_n296), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n259), .B1(new_n278), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n277), .B(KEYINPUT9), .Z(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n278), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n299), .A2(new_n259), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT73), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n302), .A2(new_n308), .A3(new_n304), .A4(new_n305), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n300), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n260), .A2(G50), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT76), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n311), .A2(new_n312), .B1(G20), .B2(new_n313), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n314), .B1(new_n312), .B2(new_n311), .C1(new_n262), .C2(new_n202), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n266), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT11), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT71), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n273), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(G33), .A2(new_n207), .B1(new_n213), .B2(new_n215), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(G68), .A3(new_n275), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n271), .A2(new_n313), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT12), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(KEYINPUT77), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT77), .B1(new_n323), .B2(new_n325), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT14), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n283), .B1(G238), .B2(new_n284), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT75), .ZN(new_n333));
  NOR2_X1   g0133(.A1(G226), .A2(G1698), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n243), .B2(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n289), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G97), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n293), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT74), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n333), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(new_n333), .B2(new_n339), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n331), .B(G169), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n343), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(G179), .A3(new_n341), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n341), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n331), .B1(new_n348), .B2(G169), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n330), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(G200), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n351), .B(new_n329), .C1(new_n352), .C2(new_n348), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n283), .B1(G244), .B2(new_n284), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G238), .A2(G1698), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n289), .B(new_n355), .C1(new_n243), .C2(G1698), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n356), .B(new_n294), .C1(G107), .C2(new_n289), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(G169), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(new_n358), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n322), .A2(G77), .A3(new_n275), .ZN(new_n362));
  INV_X1    g0162(.A(new_n263), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT65), .B(G20), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n363), .A2(new_n260), .B1(new_n364), .B2(G77), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n262), .B2(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n266), .B1(new_n202), .B2(new_n271), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n358), .A2(new_n297), .ZN(new_n372));
  AOI211_X1 g0172(.A(new_n372), .B(new_n369), .C1(G190), .C2(new_n358), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n350), .A2(new_n353), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n296), .A2(new_n360), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n277), .C1(G169), .C2(new_n296), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n310), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n363), .A2(new_n275), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n273), .A2(new_n380), .B1(new_n270), .B2(new_n363), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  INV_X1    g0183(.A(G33), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT78), .B1(new_n384), .B2(KEYINPUT3), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT78), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT3), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(G33), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(KEYINPUT3), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n217), .A2(new_n218), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n289), .B2(G20), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n313), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n383), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT79), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT79), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n383), .C1(new_n395), .C2(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n387), .A2(G33), .ZN(new_n404));
  AOI21_X1  g0204(.A(G20), .B1(new_n389), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n405), .B2(new_n391), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n364), .A2(new_n289), .A3(KEYINPUT7), .ZN(new_n407));
  OAI211_X1 g0207(.A(KEYINPUT16), .B(new_n397), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n266), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT80), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT80), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n412), .B(new_n409), .C1(new_n400), .C2(new_n402), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n382), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n283), .B1(G232), .B2(new_n284), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n289), .A2(G226), .A3(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT81), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n417), .B(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n290), .A2(G223), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n289), .A2(new_n420), .B1(G33), .B2(G87), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n416), .B1(new_n422), .B2(new_n294), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G179), .ZN(new_n424));
  INV_X1    g0224(.A(G169), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n423), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n414), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT18), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n414), .A2(new_n429), .A3(new_n426), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n422), .A2(new_n294), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(new_n352), .A3(new_n415), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G200), .B2(new_n423), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n382), .B(new_n434), .C1(new_n411), .C2(new_n413), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT17), .ZN(new_n436));
  INV_X1    g0236(.A(new_n405), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n391), .B1(new_n390), .B2(new_n392), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n397), .B1(new_n438), .B2(new_n313), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n401), .B1(new_n439), .B2(new_n383), .ZN(new_n440));
  INV_X1    g0240(.A(new_n402), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n410), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n412), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n403), .A2(KEYINPUT80), .A3(new_n410), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT17), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n382), .A4(new_n434), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT82), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n436), .A2(new_n447), .A3(KEYINPUT82), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n431), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n379), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G107), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT6), .A3(G97), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n456), .A2(KEYINPUT83), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(KEYINPUT83), .ZN(new_n458));
  XOR2_X1   g0258(.A(G97), .B(G107), .Z(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(KEYINPUT6), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n460), .A2(new_n364), .B1(G77), .B2(new_n260), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n393), .A2(new_n394), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G107), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n320), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n270), .A2(G97), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n273), .B1(new_n205), .B2(G33), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(G97), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n389), .A2(new_n404), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT4), .B1(new_n469), .B2(new_n226), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G283), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  INV_X1    g0273(.A(G244), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n289), .A2(KEYINPUT4), .A3(G244), .A4(new_n290), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n471), .A2(new_n472), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n294), .ZN(new_n478));
  INV_X1    g0278(.A(G41), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n205), .B(G45), .C1(new_n479), .C2(KEYINPUT5), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n479), .A2(KEYINPUT5), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(G257), .A3(new_n280), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(G274), .A3(new_n280), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  AOI211_X1 g0287(.A(new_n464), .B(new_n468), .C1(G200), .C2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT84), .B1(new_n487), .B2(new_n352), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT84), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n478), .A2(new_n490), .A3(G190), .A4(new_n486), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(G169), .B1(new_n478), .B2(new_n486), .ZN(new_n493));
  INV_X1    g0293(.A(new_n487), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(new_n360), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n468), .A2(new_n464), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n488), .A2(new_n492), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n269), .A2(G20), .A3(new_n455), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT25), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n466), .B2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n219), .A2(new_n289), .A3(G87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT22), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT22), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n219), .A2(new_n289), .A3(new_n505), .A4(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n364), .A2(new_n508), .A3(new_n455), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT90), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n507), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n507), .B2(new_n513), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT24), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n266), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n502), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G257), .A2(G1698), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT91), .B1(new_n469), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT91), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n289), .A2(new_n526), .A3(G257), .A4(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G294), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n289), .A2(G250), .A3(new_n290), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT92), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n289), .A2(KEYINPUT92), .A3(G250), .A4(new_n290), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n293), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n485), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n483), .A2(G264), .A3(new_n280), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n352), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n539), .B2(G200), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n523), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n225), .A2(new_n227), .A3(new_n455), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT19), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n337), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n543), .B1(new_n364), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n219), .A2(new_n289), .A3(G68), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n219), .A2(G33), .A3(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n544), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT85), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(KEYINPUT85), .A3(new_n544), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n548), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n366), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n554), .A2(new_n320), .B1(new_n270), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n466), .A2(G87), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n558), .B(KEYINPUT86), .ZN(new_n559));
  INV_X1    g0359(.A(G45), .ZN(new_n560));
  OR3_X1    g0360(.A1(new_n560), .A2(G1), .A3(G274), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n226), .B1(new_n560), .B2(G1), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n280), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n474), .A2(G1698), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n289), .B(new_n564), .C1(G238), .C2(G1698), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G116), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G190), .B(new_n563), .C1(new_n567), .C2(new_n293), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n293), .B1(new_n565), .B2(new_n566), .ZN(new_n569));
  INV_X1    g0369(.A(new_n563), .ZN(new_n570));
  OAI21_X1  g0370(.A(G200), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n557), .A2(new_n559), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n563), .B1(new_n567), .B2(new_n293), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n425), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n360), .B(new_n563), .C1(new_n567), .C2(new_n293), .ZN(new_n576));
  INV_X1    g0376(.A(new_n466), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n366), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n575), .B(new_n576), .C1(new_n556), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n498), .A2(new_n542), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n501), .B1(new_n518), .B2(new_n521), .ZN(new_n583));
  INV_X1    g0383(.A(new_n539), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n425), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n539), .A2(new_n360), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n280), .B(G270), .C1(new_n480), .C2(new_n481), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n485), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G257), .A2(G1698), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n290), .A2(G264), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n289), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT87), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n469), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n294), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n593), .B1(new_n592), .B2(new_n595), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n589), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G169), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n472), .B1(new_n227), .B2(G33), .ZN(new_n601));
  OAI22_X1  g0401(.A1(new_n364), .A2(new_n601), .B1(new_n206), .B2(G116), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT20), .ZN(new_n603));
  OR3_X1    g0403(.A1(new_n602), .A2(new_n320), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n603), .B1(new_n602), .B2(new_n320), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n271), .A2(new_n253), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n253), .B1(new_n205), .B2(G33), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n319), .A2(new_n321), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT88), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT88), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n319), .A2(new_n321), .A3(new_n613), .A4(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n600), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT21), .B1(new_n616), .B2(KEYINPUT89), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n609), .A2(new_n615), .ZN(new_n618));
  INV_X1    g0418(.A(new_n599), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(G179), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT89), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT21), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n608), .B1(new_n612), .B2(new_n614), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n600), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n587), .A2(new_n617), .A3(new_n620), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n599), .A2(G200), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n352), .B2(new_n599), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n618), .A2(new_n627), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n582), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n454), .A2(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n579), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n581), .A2(KEYINPUT26), .A3(new_n497), .A4(new_n495), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n495), .A2(new_n497), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n580), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n625), .A2(KEYINPUT93), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n498), .A2(new_n542), .A3(new_n581), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n625), .A2(KEYINPUT93), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n454), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT94), .ZN(new_n643));
  INV_X1    g0443(.A(new_n350), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n353), .A2(new_n371), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT82), .B1(new_n436), .B2(new_n447), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n436), .A2(new_n447), .A3(KEYINPUT82), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n644), .A2(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n414), .A2(new_n429), .A3(new_n426), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n429), .B1(new_n414), .B2(new_n426), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n307), .A2(new_n309), .ZN(new_n653));
  INV_X1    g0453(.A(new_n300), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n378), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n643), .A2(new_n656), .ZN(G369));
  AND3_X1   g0457(.A1(new_n617), .A2(new_n624), .A3(new_n620), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n219), .A2(new_n269), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT95), .Z(new_n660));
  INV_X1    g0460(.A(KEYINPUT27), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(G213), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n658), .A2(new_n623), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n623), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n658), .A2(new_n670), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n668), .A2(new_n671), .B1(new_n618), .B2(new_n627), .ZN(new_n672));
  INV_X1    g0472(.A(G330), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n587), .A2(new_n666), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n583), .A2(new_n666), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n542), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n675), .B1(new_n587), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n658), .A2(new_n666), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n675), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n209), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n205), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n543), .A2(G116), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n685), .A2(new_n686), .B1(new_n222), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n629), .A2(new_n667), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n589), .B(G179), .C1(new_n597), .C2(new_n598), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n574), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n535), .A2(new_n538), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n494), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT97), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n599), .A2(new_n360), .A3(new_n574), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n584), .A2(new_n487), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n696), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n494), .A2(new_n692), .A3(new_n693), .A4(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n697), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT31), .B1(new_n702), .B2(new_n666), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n690), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n641), .A2(new_n667), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n498), .A2(KEYINPUT98), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n580), .B1(new_n523), .B2(new_n541), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n498), .A2(KEYINPUT98), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n713), .A2(new_n714), .A3(new_n625), .A4(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n666), .B1(new_n716), .B2(new_n636), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n709), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n689), .B1(new_n719), .B2(G1), .ZN(G364));
  OR2_X1    g0520(.A1(new_n672), .A2(new_n673), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n364), .A2(new_n268), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G45), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n685), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n672), .A2(new_n673), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n672), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n724), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n209), .A2(new_n289), .ZN(new_n732));
  INV_X1    g0532(.A(G355), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n732), .A2(new_n733), .B1(G116), .B2(new_n209), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n683), .A2(new_n289), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n560), .B2(new_n222), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n257), .A2(G45), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n216), .B1(G20), .B2(new_n425), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n729), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n731), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n364), .A2(new_n352), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n745), .A2(G179), .A3(new_n297), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n745), .A2(new_n360), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G311), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n744), .A2(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n364), .A2(new_n352), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n751), .B1(G329), .B2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n206), .A2(new_n352), .A3(new_n297), .A4(G179), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n289), .B1(new_n756), .B2(G303), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT99), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n219), .A2(new_n360), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n352), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n752), .A2(G190), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n364), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n762), .A2(G322), .B1(G294), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n759), .A2(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n352), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(G190), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G326), .A2(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n755), .A2(new_n758), .A3(new_n765), .A4(new_n770), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT100), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G50), .A2(new_n767), .B1(new_n768), .B2(G68), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n764), .A2(G97), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n756), .A2(G87), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n775), .A3(new_n289), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(G77), .B2(new_n748), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n762), .A2(G58), .B1(new_n746), .B2(G107), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n753), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n773), .A2(new_n777), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n771), .A2(KEYINPUT100), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n772), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n743), .B1(new_n784), .B2(new_n740), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n730), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n726), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  AND2_X1   g0588(.A1(new_n666), .A2(new_n369), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n370), .B1(new_n789), .B2(new_n373), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n371), .A2(new_n667), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n710), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n792), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n641), .A2(new_n667), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n708), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT101), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n731), .B1(new_n796), .B2(new_n708), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n740), .A2(new_n727), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n724), .B1(new_n801), .B2(new_n202), .ZN(new_n802));
  INV_X1    g0602(.A(new_n740), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n746), .A2(G87), .B1(G311), .B2(new_n754), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n805), .B2(new_n761), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n289), .B1(new_n756), .B2(G107), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n807), .A2(new_n774), .ZN(new_n808));
  INV_X1    g0608(.A(new_n768), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n253), .B2(new_n749), .C1(new_n809), .C2(new_n744), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n806), .B(new_n810), .C1(G303), .C2(new_n767), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n762), .A2(G143), .B1(new_n748), .B2(G159), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n767), .A2(G137), .ZN(new_n813));
  INV_X1    g0613(.A(G150), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n809), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT34), .ZN(new_n816));
  INV_X1    g0616(.A(new_n756), .ZN(new_n817));
  INV_X1    g0617(.A(G58), .ZN(new_n818));
  INV_X1    g0618(.A(new_n764), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n289), .B1(new_n817), .B2(new_n267), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n747), .A2(new_n313), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(G132), .C2(new_n754), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n811), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n802), .B1(new_n803), .B2(new_n823), .C1(new_n794), .C2(new_n728), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n800), .A2(new_n824), .ZN(G384));
  OR2_X1    g0625(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n826), .A2(G116), .A3(new_n220), .A4(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT36), .Z(new_n829));
  OAI211_X1 g0629(.A(new_n222), .B(G77), .C1(new_n818), .C2(new_n313), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n267), .A2(G68), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n205), .B(G13), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n644), .A2(new_n667), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT39), .ZN(new_n836));
  INV_X1    g0636(.A(new_n664), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n414), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n427), .A2(new_n838), .A3(new_n839), .A4(new_n435), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n397), .B1(new_n406), .B2(new_n407), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n841), .A2(new_n383), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n382), .B1(new_n842), .B2(new_n409), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n426), .B2(new_n837), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n435), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n837), .A2(new_n843), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n452), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(KEYINPUT38), .B(new_n847), .C1(new_n452), .C2(new_n848), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n836), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n427), .A2(new_n838), .A3(new_n435), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(new_n839), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n838), .B1(new_n651), .B2(new_n448), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n850), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n852), .A2(new_n857), .A3(new_n836), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n835), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n851), .A2(new_n852), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n330), .A2(new_n666), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n350), .A2(new_n353), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n330), .B(new_n666), .C1(new_n347), .C2(new_n349), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n791), .B(KEYINPUT102), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n795), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n860), .A2(new_n867), .B1(new_n431), .B2(new_n664), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT103), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n712), .A2(new_n452), .A3(new_n379), .A4(new_n718), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n656), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n870), .B(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n792), .B1(new_n862), .B2(new_n863), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n707), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n852), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n651), .B1(new_n647), .B2(new_n646), .ZN(new_n878));
  INV_X1    g0678(.A(new_n848), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n880), .B2(new_n847), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n876), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n852), .A2(new_n857), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n707), .A2(new_n874), .A3(KEYINPUT40), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n454), .A2(new_n707), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(G330), .A3(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n873), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT105), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n894), .B1(new_n205), .B2(new_n722), .C1(new_n873), .C2(new_n892), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n893), .A2(KEYINPUT105), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n833), .B1(new_n895), .B2(new_n896), .ZN(G367));
  OAI211_X1 g0697(.A(new_n713), .B(new_n715), .C1(new_n496), .C2(new_n667), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n666), .A2(new_n495), .A3(new_n497), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT42), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n678), .A4(new_n680), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT106), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n678), .A3(new_n680), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n634), .B1(new_n898), .B2(new_n587), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n904), .A2(KEYINPUT42), .B1(new_n667), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n559), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n666), .B1(new_n556), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n909), .A2(new_n579), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n581), .A2(new_n909), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT43), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n907), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n679), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n903), .A2(new_n914), .A3(new_n913), .A4(new_n906), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n900), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n919), .ZN(new_n921));
  INV_X1    g0721(.A(new_n900), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n679), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n684), .B(KEYINPUT41), .Z(new_n924));
  INV_X1    g0724(.A(new_n681), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT45), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n925), .A2(new_n926), .A3(new_n922), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT45), .B1(new_n900), .B2(new_n681), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n918), .A2(KEYINPUT108), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT107), .B(KEYINPUT44), .C1(new_n900), .C2(new_n681), .ZN(new_n932));
  NAND2_X1  g0732(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n933));
  OR2_X1    g0733(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n922), .A2(new_n925), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n930), .A2(new_n931), .A3(new_n932), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n932), .ZN(new_n937));
  OAI211_X1 g0737(.A(KEYINPUT108), .B(new_n918), .C1(new_n929), .C2(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n678), .A2(new_n680), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n678), .A2(new_n680), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n674), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n719), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT109), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT109), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n719), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n936), .A2(new_n938), .A3(new_n944), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n924), .B1(new_n947), .B2(new_n719), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n723), .A2(G1), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n920), .B(new_n923), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n248), .A2(new_n735), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n741), .B1(new_n209), .B2(new_n366), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n817), .A2(new_n253), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT46), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT110), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n744), .B2(new_n749), .C1(new_n594), .C2(new_n761), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n469), .B1(new_n819), .B2(new_n455), .C1(new_n953), .C2(KEYINPUT46), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n746), .A2(G97), .ZN(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n753), .ZN(new_n960));
  INV_X1    g0760(.A(new_n767), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n805), .A2(new_n809), .B1(new_n961), .B2(new_n750), .ZN(new_n962));
  NOR4_X1   g0762(.A1(new_n956), .A2(new_n957), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n746), .A2(G77), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n814), .B2(new_n761), .C1(new_n749), .C2(new_n267), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n819), .A2(new_n313), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n289), .B1(new_n817), .B2(new_n818), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(G137), .C2(new_n754), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n779), .B2(new_n809), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n965), .B(new_n969), .C1(G143), .C2(new_n767), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n963), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT111), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT47), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n731), .B1(new_n951), .B2(new_n952), .C1(new_n973), .C2(new_n803), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n974), .A2(KEYINPUT112), .B1(new_n729), .B2(new_n913), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(KEYINPUT112), .B2(new_n974), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n950), .A2(new_n976), .ZN(G387));
  NAND2_X1  g0777(.A1(new_n944), .A2(new_n946), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n978), .B(new_n684), .C1(new_n719), .C2(new_n942), .ZN(new_n979));
  INV_X1    g0779(.A(G322), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n750), .A2(new_n809), .B1(new_n961), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT114), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT114), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n762), .A2(G317), .B1(new_n748), .B2(G303), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT48), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G283), .A2(new_n764), .B1(new_n756), .B2(G294), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT49), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n289), .B1(new_n754), .B2(G326), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n253), .C2(new_n747), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n768), .A2(new_n363), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n764), .A2(new_n555), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n469), .B1(new_n756), .B2(G77), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n994), .A2(new_n958), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G159), .B2(new_n767), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n748), .A2(G68), .B1(G150), .B2(new_n754), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n267), .C2(new_n761), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n803), .B1(new_n993), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n729), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n678), .A2(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n732), .A2(new_n686), .B1(G107), .B2(new_n209), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n244), .A2(G45), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n686), .ZN(new_n1006));
  AOI211_X1 g0806(.A(G45), .B(new_n1006), .C1(G68), .C2(G77), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n263), .A2(G50), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n736), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1004), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n731), .B1(new_n1011), .B2(new_n742), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n1001), .A2(new_n1003), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n942), .A2(new_n949), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT113), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(KEYINPUT113), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n979), .A2(new_n1017), .ZN(G393));
  OR3_X1    g0818(.A1(new_n929), .A2(new_n918), .A3(new_n937), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n918), .B1(new_n929), .B2(new_n937), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n949), .A3(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n254), .A2(new_n736), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n741), .B1(new_n227), .B2(new_n209), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n731), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n767), .A2(G317), .B1(new_n762), .B2(G311), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT52), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n809), .A2(new_n594), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n289), .B1(new_n756), .B2(G283), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n253), .B2(new_n819), .C1(new_n747), .C2(new_n455), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n749), .A2(new_n805), .B1(new_n980), .B2(new_n753), .ZN(new_n1030));
  NOR4_X1   g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT115), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(KEYINPUT115), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n767), .A2(G150), .B1(new_n762), .B2(G159), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT51), .Z(new_n1035));
  NAND2_X1  g0835(.A1(new_n754), .A2(G143), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n749), .B2(new_n263), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n764), .A2(G77), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n469), .B1(new_n756), .B2(G68), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n747), .C2(new_n225), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(G50), .C2(new_n768), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1035), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1032), .A2(new_n1033), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1024), .B1(new_n1043), .B2(new_n740), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n900), .B2(new_n1002), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1021), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n947), .A2(new_n684), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n978), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(G390));
  NAND4_X1  g0851(.A1(new_n707), .A2(G330), .A3(new_n794), .A4(new_n864), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n867), .A2(new_n835), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n1054), .A2(new_n853), .A3(new_n858), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n717), .A2(new_n790), .B1(new_n371), .B2(new_n667), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n834), .B1(new_n1056), .B2(new_n865), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1057), .A2(new_n886), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1053), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT39), .B1(new_n877), .B2(new_n881), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n852), .A2(new_n857), .A3(new_n836), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1060), .B(new_n1052), .C1(new_n1063), .C2(new_n1054), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n871), .B(new_n656), .C1(new_n453), .C2(new_n708), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n706), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n582), .A2(new_n625), .A3(new_n628), .A4(new_n666), .ZN(new_n1068));
  OAI211_X1 g0868(.A(G330), .B(new_n794), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n865), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n1052), .A3(new_n1056), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1052), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n795), .A2(new_n866), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1071), .A2(KEYINPUT116), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1071), .A2(KEYINPUT116), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1066), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1065), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1059), .A2(new_n1064), .A3(new_n1076), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n684), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1061), .A2(new_n727), .A3(new_n1062), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1038), .A2(new_n775), .A3(new_n469), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1082), .B(new_n821), .C1(G283), .C2(new_n767), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n455), .B2(new_n809), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n748), .A2(G97), .B1(G294), .B2(new_n754), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n253), .B2(new_n761), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n756), .A2(G150), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT53), .Z(new_n1088));
  XOR2_X1   g0888(.A(KEYINPUT54), .B(G143), .Z(new_n1089));
  NAND2_X1  g0889(.A1(new_n748), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n746), .A2(G50), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n754), .A2(G125), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n768), .A2(G137), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n767), .A2(G128), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n762), .A2(G132), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n469), .B1(new_n764), .B2(G159), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1084), .A2(new_n1086), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT117), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n803), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1100), .B2(new_n1099), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n724), .B1(new_n801), .B2(new_n263), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1081), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n949), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1080), .A2(new_n1106), .ZN(G378));
  AOI21_X1  g0907(.A(new_n834), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n860), .A2(new_n867), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n431), .A2(new_n664), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n852), .A2(new_n857), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n707), .A2(new_n874), .A3(KEYINPUT40), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n673), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n655), .A2(new_n377), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n837), .A2(new_n277), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1116), .B1(new_n310), .B2(new_n378), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n875), .B1(new_n851), .B2(new_n852), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1115), .B(new_n1124), .C1(new_n1125), .C2(new_n883), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1124), .B1(new_n885), .B2(new_n1115), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1112), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT120), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1124), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1125), .A2(new_n883), .ZN(new_n1132));
  OAI21_X1  g0932(.A(G330), .B1(new_n886), .B2(new_n887), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n869), .A3(new_n1126), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1112), .B(KEYINPUT120), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n949), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n724), .B1(new_n801), .B2(new_n267), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT119), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n961), .A2(new_n253), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n747), .A2(new_n818), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n479), .B(new_n469), .C1(new_n817), .C2(new_n202), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n1141), .A2(new_n966), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n749), .A2(new_n366), .B1(new_n744), .B2(new_n753), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G107), .B2(new_n762), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(new_n227), .C2(new_n809), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT58), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n479), .B1(new_n387), .B2(new_n384), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1147), .A2(new_n1148), .B1(new_n267), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n768), .A2(G132), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n748), .A2(G137), .B1(G150), .B2(new_n764), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n762), .A2(G128), .B1(new_n756), .B2(new_n1089), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT118), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1153), .B(new_n1155), .C1(G125), .C2(new_n767), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n384), .B(new_n479), .C1(new_n747), .C2(new_n779), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G124), .B2(new_n754), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT59), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1160), .B1(new_n1156), .B2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1150), .B1(new_n1148), .B2(new_n1147), .C1(new_n1158), .C2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1140), .B1(new_n1163), .B2(new_n740), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1131), .B2(new_n728), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1138), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n684), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1129), .A2(KEYINPUT122), .A3(new_n1135), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT122), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1112), .B(new_n1169), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1066), .B(KEYINPUT121), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n1079), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1167), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1079), .A2(new_n1173), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1172), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1166), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(G375));
  NAND2_X1  g0980(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n949), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n724), .B1(new_n801), .B2(new_n313), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1142), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n768), .A2(new_n1089), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n764), .A2(G50), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n469), .B1(new_n756), .B2(G159), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G132), .B2(new_n767), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n754), .A2(G128), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n749), .B2(new_n814), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G137), .B2(new_n762), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n253), .A2(new_n809), .B1(new_n961), .B2(new_n805), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n964), .A2(new_n469), .A3(new_n995), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n749), .A2(new_n455), .B1(new_n744), .B2(new_n761), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n754), .A2(G303), .B1(G97), .B2(new_n756), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT123), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1189), .A2(new_n1192), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1183), .B1(new_n803), .B2(new_n1199), .C1(new_n864), .C2(new_n728), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1182), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT124), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1201), .B(new_n1202), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1066), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n924), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1077), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1203), .A2(new_n1207), .ZN(G381));
  NAND3_X1  g1008(.A1(new_n979), .A2(new_n787), .A3(new_n1017), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(G381), .A2(G384), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(G378), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n950), .A2(new_n1050), .A3(new_n976), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1179), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(G407));
  NAND2_X1  g1014(.A1(new_n665), .A2(G213), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1179), .A2(new_n1211), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(G407), .A2(G213), .A3(new_n1217), .ZN(G409));
  NAND2_X1  g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1209), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1050), .B1(new_n950), .B2(new_n976), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1213), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G387), .A2(G390), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n1212), .A3(new_n1220), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT61), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT60), .B1(new_n1204), .B2(new_n1066), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1204), .A2(KEYINPUT60), .A3(new_n1066), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n684), .A3(new_n1077), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1203), .B(G384), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT124), .B1(new_n1182), .B2(new_n1200), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1232), .A2(new_n1233), .B1(new_n1230), .B2(new_n1228), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n800), .A3(new_n824), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1216), .A2(G2897), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1236), .B(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1166), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1177), .A2(new_n1172), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1176), .A2(new_n1168), .A3(KEYINPUT57), .A4(new_n1170), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n684), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G378), .B(new_n1239), .C1(new_n1240), .C2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1176), .A2(new_n1136), .A3(new_n1206), .A4(new_n1137), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1168), .A2(new_n949), .A3(new_n1170), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1165), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1211), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1215), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1227), .B1(new_n1238), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT63), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1249), .B2(new_n1236), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1216), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(KEYINPUT125), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT125), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1256), .B(new_n1216), .C1(new_n1243), .C2(new_n1247), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1236), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT63), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1255), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT126), .B1(new_n1253), .B2(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1245), .A2(new_n1165), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G378), .B1(new_n1262), .B2(new_n1244), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1179), .B2(G378), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1256), .B1(new_n1264), .B2(new_n1216), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1254), .A2(KEYINPUT125), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(KEYINPUT63), .A4(new_n1258), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1252), .A4(new_n1250), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1261), .A2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1238), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1226), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT62), .B1(new_n1254), .B2(new_n1258), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1258), .A2(KEYINPUT62), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1265), .A2(new_n1266), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1275), .B2(KEYINPUT127), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1265), .A2(new_n1266), .A3(new_n1277), .A4(new_n1274), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1272), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1270), .B1(new_n1279), .B2(new_n1281), .ZN(G405));
  NOR2_X1   g1082(.A1(new_n1179), .A2(G378), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1243), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1258), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(new_n1281), .ZN(G402));
endmodule


