

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761;

  OR2_X1 U374 ( .A1(n474), .A2(KEYINPUT118), .ZN(n419) );
  INV_X1 U375 ( .A(G953), .ZN(n472) );
  NAND2_X1 U376 ( .A1(n668), .A2(n573), .ZN(n583) );
  INV_X1 U377 ( .A(G146), .ZN(n464) );
  XNOR2_X1 U378 ( .A(n644), .B(KEYINPUT32), .ZN(n755) );
  XNOR2_X1 U379 ( .A(n623), .B(KEYINPUT93), .ZN(n757) );
  AND2_X1 U380 ( .A1(n755), .A2(n645), .ZN(n351) );
  XNOR2_X2 U381 ( .A(n616), .B(KEYINPUT0), .ZN(n625) );
  NOR2_X2 U382 ( .A1(n615), .A2(n614), .ZN(n616) );
  INV_X1 U383 ( .A(n621), .ZN(n633) );
  XNOR2_X2 U384 ( .A(G116), .B(G113), .ZN(n491) );
  XNOR2_X2 U385 ( .A(n481), .B(G469), .ZN(n581) );
  OR2_X1 U386 ( .A1(n700), .A2(n662), .ZN(n411) );
  NOR2_X1 U387 ( .A1(n633), .A2(n583), .ZN(n584) );
  XNOR2_X1 U388 ( .A(n414), .B(n413), .ZN(n646) );
  NAND2_X1 U389 ( .A1(n475), .A2(n415), .ZN(n414) );
  NOR2_X1 U390 ( .A1(n663), .A2(n661), .ZN(n432) );
  OR2_X1 U391 ( .A1(n576), .A2(n409), .ZN(n700) );
  NOR2_X1 U392 ( .A1(n597), .A2(n545), .ZN(n547) );
  XNOR2_X1 U393 ( .A(n406), .B(n577), .ZN(n663) );
  XNOR2_X1 U394 ( .A(n408), .B(n355), .ZN(n668) );
  XNOR2_X1 U395 ( .A(n461), .B(n459), .ZN(n594) );
  XNOR2_X1 U396 ( .A(n740), .B(n463), .ZN(n462) );
  XNOR2_X1 U397 ( .A(n537), .B(n538), .ZN(n463) );
  XNOR2_X1 U398 ( .A(n494), .B(G122), .ZN(n486) );
  XOR2_X1 U399 ( .A(KEYINPUT73), .B(KEYINPUT16), .Z(n494) );
  XOR2_X1 U400 ( .A(KEYINPUT67), .B(G101), .Z(n510) );
  XNOR2_X2 U401 ( .A(n468), .B(G472), .ZN(n670) );
  XNOR2_X1 U402 ( .A(n386), .B(n487), .ZN(n503) );
  XNOR2_X1 U403 ( .A(n731), .B(n485), .ZN(n386) );
  XNOR2_X1 U404 ( .A(n498), .B(n433), .ZN(n500) );
  INV_X1 U405 ( .A(KEYINPUT1), .ZN(n480) );
  XNOR2_X1 U406 ( .A(n411), .B(KEYINPUT47), .ZN(n592) );
  NAND2_X1 U407 ( .A1(n582), .A2(n658), .ZN(n588) );
  OR2_X1 U408 ( .A1(n713), .A2(G902), .ZN(n481) );
  XNOR2_X1 U409 ( .A(n360), .B(n497), .ZN(n732) );
  XNOR2_X1 U410 ( .A(KEYINPUT82), .B(G110), .ZN(n497) );
  XNOR2_X1 U411 ( .A(n570), .B(n358), .ZN(n716) );
  XNOR2_X1 U412 ( .A(G143), .B(G131), .ZN(n557) );
  XNOR2_X1 U413 ( .A(n741), .B(n464), .ZN(n524) );
  AND2_X1 U414 ( .A1(n590), .A2(n594), .ZN(n591) );
  NAND2_X1 U415 ( .A1(n373), .A2(n370), .ZN(n369) );
  NOR2_X1 U416 ( .A1(n591), .A2(n707), .ZN(n662) );
  INV_X1 U417 ( .A(n662), .ZN(n429) );
  XNOR2_X1 U418 ( .A(n629), .B(n400), .ZN(n430) );
  INV_X1 U419 ( .A(KEYINPUT88), .ZN(n400) );
  NOR2_X1 U420 ( .A1(n708), .A2(n689), .ZN(n629) );
  XNOR2_X1 U421 ( .A(G140), .B(G104), .ZN(n562) );
  INV_X1 U422 ( .A(KEYINPUT91), .ZN(n561) );
  NAND2_X1 U423 ( .A1(n598), .A2(n397), .ZN(n457) );
  XNOR2_X1 U424 ( .A(n533), .B(n354), .ZN(n566) );
  NAND2_X1 U425 ( .A1(n640), .A2(n658), .ZN(n436) );
  XNOR2_X1 U426 ( .A(n504), .B(KEYINPUT83), .ZN(n505) );
  NAND2_X1 U427 ( .A1(n503), .A2(n654), .ZN(n385) );
  NOR2_X1 U428 ( .A1(n668), .A2(n667), .ZN(n672) );
  XNOR2_X1 U429 ( .A(G902), .B(KEYINPUT15), .ZN(n654) );
  NOR2_X1 U430 ( .A1(KEYINPUT75), .A2(n651), .ZN(n650) );
  AND2_X1 U431 ( .A1(n383), .A2(n362), .ZN(n681) );
  NAND2_X1 U432 ( .A1(n353), .A2(n384), .ZN(n383) );
  INV_X1 U433 ( .A(n678), .ZN(n384) );
  XNOR2_X1 U434 ( .A(n602), .B(KEYINPUT101), .ZN(n441) );
  AND2_X1 U435 ( .A1(n477), .A2(n356), .ZN(n415) );
  NOR2_X1 U436 ( .A1(n632), .A2(n627), .ZN(n677) );
  AND2_X1 U437 ( .A1(n640), .A2(n407), .ZN(n574) );
  XNOR2_X1 U438 ( .A(n588), .B(n484), .ZN(n615) );
  INV_X1 U439 ( .A(KEYINPUT19), .ZN(n484) );
  XNOR2_X1 U440 ( .A(n571), .B(n460), .ZN(n459) );
  OR2_X1 U441 ( .A1(n716), .A2(G902), .ZN(n461) );
  INV_X1 U442 ( .A(G475), .ZN(n460) );
  XNOR2_X1 U443 ( .A(n524), .B(n424), .ZN(n713) );
  XNOR2_X1 U444 ( .A(n525), .B(n425), .ZN(n424) );
  XNOR2_X1 U445 ( .A(n426), .B(n526), .ZN(n425) );
  NAND2_X1 U446 ( .A1(n352), .A2(n437), .ZN(n645) );
  NAND2_X1 U447 ( .A1(n627), .A2(n372), .ZN(n371) );
  INV_X1 U448 ( .A(KEYINPUT116), .ZN(n372) );
  AND2_X1 U449 ( .A1(n375), .A2(n374), .ZN(n373) );
  NAND2_X1 U450 ( .A1(n404), .A2(KEYINPUT116), .ZN(n374) );
  XNOR2_X1 U451 ( .A(n496), .B(G128), .ZN(n515) );
  INV_X1 U452 ( .A(G143), .ZN(n496) );
  XNOR2_X1 U453 ( .A(n499), .B(n434), .ZN(n433) );
  INV_X1 U454 ( .A(KEYINPUT4), .ZN(n434) );
  XOR2_X1 U455 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n499) );
  XNOR2_X1 U456 ( .A(n382), .B(n381), .ZN(n380) );
  INV_X1 U457 ( .A(KEYINPUT51), .ZN(n381) );
  OR2_X1 U458 ( .A1(n676), .A2(n677), .ZN(n382) );
  OR2_X1 U459 ( .A1(G237), .A2(G902), .ZN(n518) );
  INV_X1 U460 ( .A(KEYINPUT48), .ZN(n456) );
  XNOR2_X1 U461 ( .A(n491), .B(n490), .ZN(n493) );
  NAND2_X1 U462 ( .A1(n388), .A2(n390), .ZN(n387) );
  AND2_X1 U463 ( .A1(n391), .A2(KEYINPUT94), .ZN(n390) );
  AND2_X1 U464 ( .A1(n392), .A2(n630), .ZN(n388) );
  NAND2_X1 U465 ( .A1(n393), .A2(n630), .ZN(n389) );
  NAND2_X1 U466 ( .A1(n757), .A2(n399), .ZN(n395) );
  XNOR2_X1 U467 ( .A(n515), .B(n514), .ZN(n550) );
  INV_X1 U468 ( .A(G134), .ZN(n514) );
  XNOR2_X1 U469 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U470 ( .A(G122), .B(G113), .Z(n558) );
  XNOR2_X1 U471 ( .A(n550), .B(n516), .ZN(n741) );
  XOR2_X1 U472 ( .A(KEYINPUT4), .B(G131), .Z(n516) );
  XOR2_X1 U473 ( .A(G137), .B(G140), .Z(n534) );
  INV_X1 U474 ( .A(n588), .ZN(n454) );
  OR2_X1 U475 ( .A1(n684), .A2(G902), .ZN(n468) );
  XNOR2_X1 U476 ( .A(n670), .B(n442), .ZN(n621) );
  INV_X1 U477 ( .A(KEYINPUT6), .ZN(n442) );
  INV_X1 U478 ( .A(KEYINPUT23), .ZN(n535) );
  XNOR2_X1 U479 ( .A(G128), .B(G110), .ZN(n536) );
  XNOR2_X1 U480 ( .A(n566), .B(n534), .ZN(n740) );
  XNOR2_X1 U481 ( .A(G116), .B(G107), .ZN(n548) );
  XOR2_X1 U482 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n531) );
  XNOR2_X1 U483 ( .A(n483), .B(n732), .ZN(n525) );
  XNOR2_X1 U484 ( .A(n438), .B(n482), .ZN(n426) );
  INV_X1 U485 ( .A(KEYINPUT84), .ZN(n482) );
  INV_X1 U486 ( .A(n534), .ZN(n438) );
  NOR2_X1 U487 ( .A1(n437), .A2(n450), .ZN(n449) );
  NOR2_X1 U488 ( .A1(n454), .A2(n586), .ZN(n450) );
  XNOR2_X1 U489 ( .A(n600), .B(KEYINPUT107), .ZN(n455) );
  XNOR2_X1 U490 ( .A(n585), .B(KEYINPUT36), .ZN(n586) );
  INV_X1 U491 ( .A(KEYINPUT80), .ZN(n585) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n544) );
  INV_X1 U493 ( .A(KEYINPUT30), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n670), .B(n467), .ZN(n640) );
  INV_X1 U495 ( .A(KEYINPUT95), .ZN(n467) );
  XNOR2_X1 U496 ( .A(n620), .B(n488), .ZN(n639) );
  XNOR2_X1 U497 ( .A(n489), .B(KEYINPUT22), .ZN(n488) );
  INV_X1 U498 ( .A(KEYINPUT65), .ZN(n489) );
  BUF_X1 U499 ( .A(n625), .Z(n636) );
  OR2_X1 U500 ( .A1(n722), .A2(G902), .ZN(n408) );
  XNOR2_X1 U501 ( .A(n502), .B(n501), .ZN(n655) );
  NAND2_X1 U502 ( .A1(n681), .A2(n473), .ZN(n418) );
  AND2_X1 U503 ( .A1(n421), .A2(n472), .ZN(n420) );
  NAND2_X1 U504 ( .A1(n422), .A2(KEYINPUT118), .ZN(n421) );
  INV_X1 U505 ( .A(n681), .ZN(n422) );
  AND2_X1 U506 ( .A1(n441), .A2(n437), .ZN(n603) );
  XNOR2_X1 U507 ( .A(n471), .B(n469), .ZN(n751) );
  XNOR2_X1 U508 ( .A(n470), .B(KEYINPUT104), .ZN(n469) );
  INV_X1 U509 ( .A(KEYINPUT40), .ZN(n470) );
  INV_X1 U510 ( .A(KEYINPUT35), .ZN(n413) );
  NAND2_X1 U511 ( .A1(n625), .A2(n677), .ZN(n443) );
  NAND2_X1 U512 ( .A1(n412), .A2(n410), .ZN(n409) );
  INV_X1 U513 ( .A(n575), .ZN(n410) );
  INV_X1 U514 ( .A(n615), .ZN(n412) );
  AND2_X1 U515 ( .A1(n636), .A2(n403), .ZN(n689) );
  NOR2_X1 U516 ( .A1(n628), .A2(n404), .ZN(n403) );
  INV_X1 U517 ( .A(KEYINPUT60), .ZN(n401) );
  XNOR2_X1 U518 ( .A(n711), .B(n440), .ZN(n714) );
  INV_X1 U519 ( .A(n645), .ZN(n693) );
  AND2_X1 U520 ( .A1(n641), .A2(n668), .ZN(n352) );
  XOR2_X1 U521 ( .A(n359), .B(KEYINPUT52), .Z(n353) );
  XOR2_X1 U522 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n354) );
  XOR2_X1 U523 ( .A(n542), .B(n541), .Z(n355) );
  AND2_X1 U524 ( .A1(n478), .A2(n638), .ZN(n356) );
  OR2_X1 U525 ( .A1(n680), .A2(n666), .ZN(n357) );
  XOR2_X1 U526 ( .A(n558), .B(n557), .Z(n358) );
  AND2_X1 U527 ( .A1(n378), .A2(n357), .ZN(n359) );
  XOR2_X1 U528 ( .A(G104), .B(G107), .Z(n360) );
  AND2_X1 U529 ( .A1(n636), .A2(n479), .ZN(n361) );
  INV_X1 U530 ( .A(n437), .ZN(n671) );
  INV_X1 U531 ( .A(n627), .ZN(n404) );
  OR2_X1 U532 ( .A1(n680), .A2(n679), .ZN(n362) );
  AND2_X1 U533 ( .A1(n454), .A2(n586), .ZN(n363) );
  AND2_X1 U534 ( .A1(n429), .A2(n399), .ZN(n364) );
  XNOR2_X1 U535 ( .A(n443), .B(n626), .ZN(n708) );
  INV_X1 U536 ( .A(KEYINPUT34), .ZN(n479) );
  XOR2_X1 U537 ( .A(n686), .B(n685), .Z(n365) );
  XOR2_X1 U538 ( .A(n716), .B(n715), .Z(n366) );
  INV_X1 U539 ( .A(KEYINPUT94), .ZN(n399) );
  XOR2_X1 U540 ( .A(n656), .B(KEYINPUT56), .Z(n367) );
  XOR2_X1 U541 ( .A(n683), .B(n682), .Z(n368) );
  NOR2_X1 U542 ( .A1(G952), .A2(n472), .ZN(n724) );
  INV_X1 U543 ( .A(n724), .ZN(n446) );
  INV_X1 U544 ( .A(KEYINPUT118), .ZN(n473) );
  XNOR2_X1 U545 ( .A(n464), .B(G125), .ZN(n533) );
  NOR2_X1 U546 ( .A1(n674), .A2(n369), .ZN(n675) );
  OR2_X1 U547 ( .A1(n376), .A2(n371), .ZN(n370) );
  NAND2_X1 U548 ( .A1(n376), .A2(KEYINPUT116), .ZN(n375) );
  XNOR2_X1 U549 ( .A(n669), .B(n377), .ZN(n376) );
  INV_X1 U550 ( .A(KEYINPUT49), .ZN(n377) );
  NAND2_X1 U551 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U552 ( .A(n679), .ZN(n379) );
  XNOR2_X2 U553 ( .A(n385), .B(n505), .ZN(n582) );
  NAND2_X1 U554 ( .A1(n389), .A2(n387), .ZN(n648) );
  NAND2_X1 U555 ( .A1(n430), .A2(n429), .ZN(n391) );
  INV_X1 U556 ( .A(n757), .ZN(n392) );
  NAND2_X1 U557 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U558 ( .A1(n430), .A2(n364), .ZN(n394) );
  XNOR2_X1 U559 ( .A(n427), .B(n649), .ZN(n725) );
  NAND2_X1 U560 ( .A1(n405), .A2(G475), .ZN(n717) );
  NOR2_X4 U561 ( .A1(n657), .A2(n654), .ZN(n405) );
  XNOR2_X1 U562 ( .A(n396), .B(n647), .ZN(n431) );
  NAND2_X1 U563 ( .A1(n351), .A2(n646), .ZN(n396) );
  XNOR2_X1 U564 ( .A(n687), .B(n365), .ZN(n447) );
  NAND2_X1 U565 ( .A1(n637), .A2(KEYINPUT34), .ZN(n478) );
  NOR2_X1 U566 ( .A1(n760), .A2(n458), .ZN(n397) );
  NAND2_X1 U567 ( .A1(n465), .A2(n446), .ZN(n439) );
  NOR2_X2 U568 ( .A1(n639), .A2(n621), .ZN(n643) );
  XNOR2_X1 U569 ( .A(n466), .B(n655), .ZN(n465) );
  NAND2_X1 U570 ( .A1(n659), .A2(n658), .ZN(n406) );
  XNOR2_X1 U571 ( .A(n432), .B(KEYINPUT41), .ZN(n679) );
  NOR2_X2 U572 ( .A1(n754), .A2(n751), .ZN(n580) );
  XNOR2_X1 U573 ( .A(n579), .B(n578), .ZN(n754) );
  NAND2_X1 U574 ( .A1(n398), .A2(n704), .ZN(n600) );
  XNOR2_X1 U575 ( .A(n584), .B(KEYINPUT100), .ZN(n398) );
  NAND2_X1 U576 ( .A1(n447), .A2(n446), .ZN(n445) );
  XNOR2_X1 U577 ( .A(n547), .B(n546), .ZN(n607) );
  XNOR2_X1 U578 ( .A(n539), .B(n462), .ZN(n722) );
  XNOR2_X1 U579 ( .A(n402), .B(n401), .ZN(G60) );
  NAND2_X1 U580 ( .A1(n428), .A2(n446), .ZN(n402) );
  NAND2_X1 U581 ( .A1(n405), .A2(G472), .ZN(n687) );
  NAND2_X1 U582 ( .A1(n405), .A2(G210), .ZN(n466) );
  NAND2_X1 U583 ( .A1(n405), .A2(G478), .ZN(n718) );
  NAND2_X1 U584 ( .A1(n405), .A2(G469), .ZN(n711) );
  NAND2_X1 U585 ( .A1(n405), .A2(G217), .ZN(n721) );
  XNOR2_X2 U586 ( .A(n605), .B(n506), .ZN(n659) );
  INV_X1 U587 ( .A(n583), .ZN(n407) );
  OR2_X1 U588 ( .A1(n576), .A2(n575), .ZN(n589) );
  INV_X1 U589 ( .A(n646), .ZN(n753) );
  NAND2_X1 U590 ( .A1(n416), .A2(n420), .ZN(n423) );
  NAND2_X1 U591 ( .A1(n419), .A2(n417), .ZN(n416) );
  NAND2_X1 U592 ( .A1(n474), .A2(n418), .ZN(n417) );
  XNOR2_X1 U593 ( .A(n423), .B(n368), .ZN(G75) );
  NAND2_X1 U594 ( .A1(n648), .A2(n431), .ZN(n427) );
  XNOR2_X1 U595 ( .A(n445), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U596 ( .A1(n639), .A2(n640), .ZN(n641) );
  XNOR2_X1 U597 ( .A(n581), .B(n480), .ZN(n599) );
  XNOR2_X1 U598 ( .A(n717), .B(n366), .ZN(n428) );
  OR2_X1 U599 ( .A1(n592), .A2(n698), .ZN(n458) );
  NAND2_X1 U600 ( .A1(n607), .A2(n591), .ZN(n471) );
  BUF_X1 U601 ( .A(n599), .Z(n437) );
  XNOR2_X1 U602 ( .A(n510), .B(KEYINPUT71), .ZN(n483) );
  XNOR2_X1 U603 ( .A(n439), .B(n367), .ZN(G51) );
  XNOR2_X1 U604 ( .A(n657), .B(KEYINPUT78), .ZN(n474) );
  OR2_X2 U605 ( .A1(n632), .A2(n633), .ZN(n635) );
  XNOR2_X1 U606 ( .A(n624), .B(KEYINPUT74), .ZN(n632) );
  XNOR2_X1 U607 ( .A(n713), .B(n712), .ZN(n440) );
  XNOR2_X1 U608 ( .A(n512), .B(n513), .ZN(n517) );
  INV_X1 U609 ( .A(n600), .ZN(n601) );
  NOR2_X1 U610 ( .A1(n759), .A2(n608), .ZN(n609) );
  XNOR2_X1 U611 ( .A(n606), .B(KEYINPUT102), .ZN(n759) );
  INV_X1 U612 ( .A(n599), .ZN(n453) );
  XNOR2_X1 U613 ( .A(n444), .B(n650), .ZN(n653) );
  NAND2_X1 U614 ( .A1(n725), .A2(n743), .ZN(n444) );
  NAND2_X1 U615 ( .A1(n455), .A2(n363), .ZN(n451) );
  NOR2_X1 U616 ( .A1(n452), .A2(n448), .ZN(n587) );
  NAND2_X1 U617 ( .A1(n451), .A2(n449), .ZN(n448) );
  NOR2_X1 U618 ( .A1(n455), .A2(n586), .ZN(n452) );
  XNOR2_X1 U619 ( .A(n457), .B(n456), .ZN(n610) );
  NAND2_X1 U620 ( .A1(n476), .A2(n361), .ZN(n475) );
  INV_X1 U621 ( .A(n680), .ZN(n476) );
  NAND2_X1 U622 ( .A1(n680), .A2(KEYINPUT34), .ZN(n477) );
  XNOR2_X2 U623 ( .A(n635), .B(n634), .ZN(n680) );
  XNOR2_X1 U624 ( .A(n515), .B(n495), .ZN(n485) );
  XNOR2_X2 U625 ( .A(n511), .B(n486), .ZN(n731) );
  XNOR2_X1 U626 ( .A(n500), .B(n525), .ZN(n487) );
  INV_X1 U627 ( .A(KEYINPUT70), .ZN(n490) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(n565) );
  INV_X1 U629 ( .A(n710), .ZN(n608) );
  XNOR2_X1 U630 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U631 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n578) );
  XNOR2_X1 U632 ( .A(KEYINPUT55), .B(KEYINPUT81), .ZN(n502) );
  XOR2_X1 U633 ( .A(KEYINPUT3), .B(G119), .Z(n492) );
  XNOR2_X2 U634 ( .A(n493), .B(n492), .ZN(n511) );
  INV_X1 U635 ( .A(n533), .ZN(n495) );
  NAND2_X1 U636 ( .A1(G224), .A2(n472), .ZN(n498) );
  XNOR2_X1 U637 ( .A(n503), .B(KEYINPUT54), .ZN(n501) );
  INV_X1 U638 ( .A(KEYINPUT38), .ZN(n506) );
  NAND2_X1 U639 ( .A1(G210), .A2(n518), .ZN(n504) );
  BUF_X1 U640 ( .A(n582), .Z(n605) );
  INV_X1 U641 ( .A(n659), .ZN(n545) );
  XOR2_X1 U642 ( .A(G137), .B(KEYINPUT86), .Z(n508) );
  NOR2_X1 U643 ( .A1(G953), .A2(G237), .ZN(n567) );
  NAND2_X1 U644 ( .A1(n567), .A2(G210), .ZN(n507) );
  XNOR2_X1 U645 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U646 ( .A(n509), .B(KEYINPUT5), .Z(n513) );
  XNOR2_X1 U647 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U648 ( .A(n517), .B(n524), .ZN(n684) );
  NAND2_X1 U649 ( .A1(G214), .A2(n518), .ZN(n658) );
  NAND2_X1 U650 ( .A1(G234), .A2(G237), .ZN(n519) );
  XNOR2_X1 U651 ( .A(n519), .B(KEYINPUT14), .ZN(n520) );
  NAND2_X1 U652 ( .A1(n520), .A2(G952), .ZN(n678) );
  NOR2_X1 U653 ( .A1(G953), .A2(n678), .ZN(n613) );
  NAND2_X1 U654 ( .A1(n520), .A2(G902), .ZN(n611) );
  OR2_X1 U655 ( .A1(n472), .A2(n611), .ZN(n521) );
  XOR2_X1 U656 ( .A(KEYINPUT99), .B(n521), .Z(n522) );
  NOR2_X1 U657 ( .A1(G900), .A2(n522), .ZN(n523) );
  NOR2_X1 U658 ( .A1(n613), .A2(n523), .ZN(n572) );
  NAND2_X1 U659 ( .A1(G227), .A2(n472), .ZN(n526) );
  XOR2_X1 U660 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n529) );
  NAND2_X1 U661 ( .A1(G234), .A2(n654), .ZN(n527) );
  XNOR2_X1 U662 ( .A(KEYINPUT20), .B(n527), .ZN(n540) );
  NAND2_X1 U663 ( .A1(n540), .A2(G221), .ZN(n528) );
  XNOR2_X1 U664 ( .A(n529), .B(n528), .ZN(n667) );
  NAND2_X1 U665 ( .A1(G234), .A2(n472), .ZN(n530) );
  XNOR2_X1 U666 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U667 ( .A(KEYINPUT77), .B(n532), .Z(n553) );
  NAND2_X1 U668 ( .A1(G221), .A2(n553), .ZN(n539) );
  XOR2_X1 U669 ( .A(G119), .B(KEYINPUT24), .Z(n538) );
  XOR2_X1 U670 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n542) );
  NAND2_X1 U671 ( .A1(n540), .A2(G217), .ZN(n541) );
  NAND2_X1 U672 ( .A1(n581), .A2(n672), .ZN(n628) );
  NOR2_X1 U673 ( .A1(n572), .A2(n628), .ZN(n543) );
  NAND2_X1 U674 ( .A1(n544), .A2(n543), .ZN(n597) );
  XNOR2_X1 U675 ( .A(KEYINPUT79), .B(KEYINPUT39), .ZN(n546) );
  XNOR2_X1 U676 ( .A(n548), .B(KEYINPUT7), .ZN(n549) );
  XOR2_X1 U677 ( .A(n549), .B(KEYINPUT9), .Z(n552) );
  XNOR2_X1 U678 ( .A(n550), .B(G122), .ZN(n551) );
  XNOR2_X1 U679 ( .A(n552), .B(n551), .ZN(n555) );
  NAND2_X1 U680 ( .A1(G217), .A2(n553), .ZN(n554) );
  XOR2_X1 U681 ( .A(n554), .B(n555), .Z(n719) );
  NOR2_X1 U682 ( .A1(G902), .A2(n719), .ZN(n556) );
  XNOR2_X1 U683 ( .A(G478), .B(n556), .ZN(n590) );
  XNOR2_X1 U684 ( .A(KEYINPUT92), .B(KEYINPUT13), .ZN(n571) );
  XOR2_X1 U685 ( .A(KEYINPUT11), .B(KEYINPUT90), .Z(n560) );
  XNOR2_X1 U686 ( .A(KEYINPUT89), .B(KEYINPUT12), .ZN(n559) );
  XNOR2_X1 U687 ( .A(n560), .B(n559), .ZN(n564) );
  XNOR2_X1 U688 ( .A(n566), .B(n565), .ZN(n569) );
  NAND2_X1 U689 ( .A1(G214), .A2(n567), .ZN(n568) );
  XNOR2_X1 U690 ( .A(n569), .B(n568), .ZN(n570) );
  NOR2_X1 U691 ( .A1(n667), .A2(n572), .ZN(n573) );
  XOR2_X1 U692 ( .A(KEYINPUT28), .B(n574), .Z(n576) );
  XNOR2_X1 U693 ( .A(n581), .B(KEYINPUT103), .ZN(n575) );
  INV_X1 U694 ( .A(KEYINPUT105), .ZN(n577) );
  INV_X1 U695 ( .A(n590), .ZN(n593) );
  NOR2_X1 U696 ( .A1(n594), .A2(n593), .ZN(n617) );
  INV_X1 U697 ( .A(n617), .ZN(n661) );
  NOR2_X1 U698 ( .A1(n589), .A2(n679), .ZN(n579) );
  XNOR2_X1 U699 ( .A(n580), .B(KEYINPUT46), .ZN(n598) );
  XOR2_X1 U700 ( .A(KEYINPUT98), .B(n591), .Z(n701) );
  XNOR2_X1 U701 ( .A(KEYINPUT108), .B(n587), .ZN(n760) );
  NOR2_X1 U702 ( .A1(n590), .A2(n594), .ZN(n707) );
  NAND2_X1 U703 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U704 ( .A(n595), .B(KEYINPUT97), .ZN(n638) );
  NAND2_X1 U705 ( .A1(n605), .A2(n638), .ZN(n596) );
  NOR2_X1 U706 ( .A1(n597), .A2(n596), .ZN(n698) );
  NAND2_X1 U707 ( .A1(n601), .A2(n658), .ZN(n602) );
  XNOR2_X1 U708 ( .A(n603), .B(KEYINPUT43), .ZN(n604) );
  NOR2_X1 U709 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U710 ( .A1(n707), .A2(n607), .ZN(n710) );
  AND2_X2 U711 ( .A1(n610), .A2(n609), .ZN(n743) );
  OR2_X1 U712 ( .A1(n472), .A2(G898), .ZN(n737) );
  NOR2_X1 U713 ( .A1(n611), .A2(n737), .ZN(n612) );
  NOR2_X1 U714 ( .A1(n613), .A2(n612), .ZN(n614) );
  INV_X1 U715 ( .A(n667), .ZN(n618) );
  AND2_X1 U716 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U717 ( .A1(n625), .A2(n619), .ZN(n620) );
  NOR2_X1 U718 ( .A1(n671), .A2(n668), .ZN(n622) );
  NAND2_X1 U719 ( .A1(n643), .A2(n622), .ZN(n623) );
  XOR2_X1 U720 ( .A(KEYINPUT31), .B(KEYINPUT87), .Z(n626) );
  NAND2_X1 U721 ( .A1(n453), .A2(n672), .ZN(n624) );
  INV_X1 U722 ( .A(n670), .ZN(n627) );
  INV_X1 U723 ( .A(KEYINPUT72), .ZN(n631) );
  NAND2_X1 U724 ( .A1(n631), .A2(KEYINPUT44), .ZN(n630) );
  NOR2_X1 U725 ( .A1(n631), .A2(KEYINPUT44), .ZN(n647) );
  XOR2_X1 U726 ( .A(KEYINPUT96), .B(KEYINPUT33), .Z(n634) );
  INV_X1 U727 ( .A(n636), .ZN(n637) );
  AND2_X1 U728 ( .A1(n671), .A2(n668), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U730 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n649) );
  INV_X1 U731 ( .A(KEYINPUT2), .ZN(n651) );
  NAND2_X1 U732 ( .A1(KEYINPUT75), .A2(n651), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n657) );
  INV_X1 U734 ( .A(KEYINPUT121), .ZN(n656) );
  NOR2_X1 U735 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U736 ( .A1(n661), .A2(n660), .ZN(n665) );
  NOR2_X1 U737 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n666) );
  AND2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U741 ( .A(KEYINPUT50), .B(n673), .ZN(n674) );
  XOR2_X1 U742 ( .A(KEYINPUT117), .B(n675), .Z(n676) );
  XNOR2_X1 U743 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n683) );
  INV_X1 U744 ( .A(KEYINPUT53), .ZN(n682) );
  XOR2_X1 U745 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n686) );
  XNOR2_X1 U746 ( .A(n684), .B(KEYINPUT110), .ZN(n685) );
  INV_X1 U747 ( .A(n701), .ZN(n704) );
  NAND2_X1 U748 ( .A1(n704), .A2(n689), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n688), .B(G104), .ZN(G6) );
  XOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n691) );
  NAND2_X1 U751 ( .A1(n689), .A2(n707), .ZN(n690) );
  XNOR2_X1 U752 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U753 ( .A(G107), .B(n692), .ZN(G9) );
  XOR2_X1 U754 ( .A(G110), .B(n693), .Z(G12) );
  INV_X1 U755 ( .A(n707), .ZN(n694) );
  NOR2_X1 U756 ( .A1(n694), .A2(n700), .ZN(n696) );
  XNOR2_X1 U757 ( .A(KEYINPUT29), .B(KEYINPUT112), .ZN(n695) );
  XNOR2_X1 U758 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U759 ( .A(G128), .B(n697), .ZN(G30) );
  XNOR2_X1 U760 ( .A(G143), .B(n698), .ZN(n699) );
  XNOR2_X1 U761 ( .A(n699), .B(KEYINPUT113), .ZN(G45) );
  NOR2_X1 U762 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U763 ( .A(KEYINPUT114), .B(n702), .Z(n703) );
  XNOR2_X1 U764 ( .A(G146), .B(n703), .ZN(G48) );
  XOR2_X1 U765 ( .A(G113), .B(KEYINPUT115), .Z(n706) );
  NAND2_X1 U766 ( .A1(n708), .A2(n704), .ZN(n705) );
  XNOR2_X1 U767 ( .A(n706), .B(n705), .ZN(G15) );
  NAND2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U769 ( .A(n709), .B(G116), .ZN(G18) );
  XNOR2_X1 U770 ( .A(G134), .B(n710), .ZN(G36) );
  XOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  NOR2_X1 U772 ( .A1(n724), .A2(n714), .ZN(G54) );
  XOR2_X1 U773 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n715) );
  XNOR2_X1 U774 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U775 ( .A1(n724), .A2(n720), .ZN(G63) );
  XNOR2_X1 U776 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n724), .A2(n723), .ZN(G66) );
  NAND2_X1 U778 ( .A1(n725), .A2(n472), .ZN(n730) );
  NAND2_X1 U779 ( .A1(G224), .A2(G953), .ZN(n726) );
  XNOR2_X1 U780 ( .A(n726), .B(KEYINPUT61), .ZN(n727) );
  XNOR2_X1 U781 ( .A(KEYINPUT122), .B(n727), .ZN(n728) );
  NAND2_X1 U782 ( .A1(G898), .A2(n728), .ZN(n729) );
  NAND2_X1 U783 ( .A1(n730), .A2(n729), .ZN(n739) );
  XOR2_X1 U784 ( .A(G101), .B(KEYINPUT123), .Z(n735) );
  XNOR2_X1 U785 ( .A(n731), .B(n732), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n733), .B(KEYINPUT124), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U788 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U789 ( .A(n739), .B(n738), .Z(G69) );
  XNOR2_X1 U790 ( .A(KEYINPUT84), .B(n740), .ZN(n742) );
  XOR2_X1 U791 ( .A(n741), .B(n742), .Z(n745) );
  XOR2_X1 U792 ( .A(n745), .B(n743), .Z(n744) );
  NAND2_X1 U793 ( .A1(n744), .A2(n472), .ZN(n749) );
  XNOR2_X1 U794 ( .A(n745), .B(G227), .ZN(n746) );
  NOR2_X1 U795 ( .A1(n472), .A2(n746), .ZN(n747) );
  NAND2_X1 U796 ( .A1(G900), .A2(n747), .ZN(n748) );
  NAND2_X1 U797 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U798 ( .A(KEYINPUT125), .B(n750), .ZN(G72) );
  XNOR2_X1 U799 ( .A(n751), .B(G131), .ZN(n752) );
  XNOR2_X1 U800 ( .A(n752), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U801 ( .A(n753), .B(G122), .Z(G24) );
  XOR2_X1 U802 ( .A(G137), .B(n754), .Z(G39) );
  XNOR2_X1 U803 ( .A(G119), .B(n755), .ZN(n756) );
  XNOR2_X1 U804 ( .A(n756), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U805 ( .A(G101), .B(n757), .ZN(n758) );
  XNOR2_X1 U806 ( .A(n758), .B(KEYINPUT111), .ZN(G3) );
  XOR2_X1 U807 ( .A(n759), .B(G140), .Z(G42) );
  XNOR2_X1 U808 ( .A(G125), .B(KEYINPUT37), .ZN(n761) );
  XNOR2_X1 U809 ( .A(n761), .B(n760), .ZN(G27) );
endmodule

