//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1305, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G1), .B2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n206), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n208), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n211), .B(new_n220), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n222), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n247), .B(new_n253), .ZN(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n216), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n206), .A2(G116), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G97), .ZN(new_n260));
  AOI21_X1  g0060(.A(G20), .B1(G33), .B2(G283), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n258), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n257), .A2(KEYINPUT20), .A3(new_n262), .ZN(new_n266));
  INV_X1    g0066(.A(G13), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n265), .A2(new_n266), .B1(new_n268), .B2(new_n258), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n256), .A2(new_n216), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n256), .A2(new_n216), .A3(KEYINPUT70), .A4(new_n270), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n259), .A2(G1), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n273), .A2(G116), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n269), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n205), .B(G45), .C1(new_n281), .C2(KEYINPUT5), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT79), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n282), .B2(KEYINPUT79), .ZN(new_n286));
  OAI211_X1 g0086(.A(G270), .B(new_n280), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n282), .A2(KEYINPUT79), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  INV_X1    g0089(.A(new_n214), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n279), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n288), .A2(new_n283), .A3(new_n285), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n279), .B1(new_n213), .B2(new_n215), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G257), .A2(G1698), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n231), .B2(G1698), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G303), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n294), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(G200), .B1(new_n293), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT80), .B1(new_n278), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n293), .A2(new_n306), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G190), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT80), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n269), .A2(new_n307), .A3(new_n312), .A4(new_n277), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT3), .B(G33), .ZN(new_n315));
  INV_X1    g0115(.A(G1698), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(G222), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(G223), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n317), .B1(new_n228), .B2(new_n315), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n294), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G45), .ZN(new_n323));
  AOI21_X1  g0123(.A(G1), .B1(new_n281), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(new_n280), .A3(G274), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n280), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G226), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT66), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n329), .A2(new_n330), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n322), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G200), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(new_n333), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n206), .A2(G33), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT68), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT8), .B(G58), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n206), .A2(new_n259), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n270), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n345), .A2(new_n257), .B1(new_n248), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n271), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n205), .A2(G20), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(G50), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT9), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT9), .B1(new_n347), .B2(new_n350), .ZN(new_n355));
  NOR4_X1   g0155(.A1(new_n336), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n333), .A2(G179), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n333), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n351), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  NOR2_X1   g0165(.A1(G223), .A2(G1698), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n328), .B2(G1698), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n302), .A2(KEYINPUT73), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n370), .A3(G33), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n371), .A3(new_n295), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n259), .A2(new_n224), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n321), .ZN(new_n376));
  INV_X1    g0176(.A(new_n327), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G232), .B1(new_n291), .B2(new_n324), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n361), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n294), .B1(new_n372), .B2(new_n374), .ZN(new_n380));
  INV_X1    g0180(.A(G179), .ZN(new_n381));
  INV_X1    g0181(.A(G232), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n325), .B1(new_n327), .B2(new_n382), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n365), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(G169), .B1(new_n380), .B2(new_n383), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n373), .B1(new_n298), .B2(new_n367), .ZN(new_n387));
  OAI211_X1 g0187(.A(G179), .B(new_n378), .C1(new_n387), .C2(new_n294), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n388), .A3(KEYINPUT77), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n339), .B1(new_n205), .B2(G20), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n348), .A2(new_n391), .B1(new_n346), .B2(new_n339), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n214), .B(KEYINPUT64), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND3_X1   g0197(.A1(KEYINPUT74), .A2(G58), .A3(G68), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT74), .B1(G58), .B2(G68), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n206), .B1(new_n400), .B2(new_n202), .ZN(new_n401));
  INV_X1    g0201(.A(G159), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n344), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n303), .B1(new_n297), .B2(G33), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(G20), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n304), .A2(new_n206), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n405), .A2(new_n407), .B1(new_n408), .B2(new_n406), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n404), .B1(new_n409), .B2(new_n222), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n397), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT75), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n401), .B2(new_n403), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n398), .A2(new_n399), .A3(new_n201), .ZN(new_n415));
  OAI221_X1 g0215(.A(KEYINPUT75), .B1(new_n402), .B2(new_n344), .C1(new_n415), .C2(new_n206), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT7), .B1(new_n298), .B2(G20), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n371), .A2(new_n295), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(new_n406), .A3(new_n206), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(G68), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n421), .A3(KEYINPUT16), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n393), .B1(new_n412), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n390), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT18), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n410), .A2(new_n411), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n426), .A3(new_n257), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT78), .ZN(new_n428));
  AOI21_X1  g0228(.A(G200), .B1(new_n376), .B2(new_n378), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n380), .A2(G190), .A3(new_n383), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n376), .A2(new_n335), .A3(new_n378), .ZN(new_n432));
  INV_X1    g0232(.A(G200), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n380), .B2(new_n383), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(KEYINPUT78), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n427), .A2(new_n431), .A3(new_n435), .A4(new_n392), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n425), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n315), .A2(G226), .A3(new_n316), .ZN(new_n439));
  INV_X1    g0239(.A(G97), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n259), .B2(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n304), .A2(new_n382), .A3(new_n316), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n321), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT13), .ZN(new_n444));
  INV_X1    g0244(.A(new_n325), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(G238), .B2(new_n377), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n444), .B1(new_n443), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g0249(.A(G200), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n273), .A2(G68), .A3(new_n274), .A4(new_n349), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n338), .A2(G77), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n344), .A2(new_n248), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(G20), .B2(new_n222), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n397), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n455), .A2(KEYINPUT11), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n270), .A2(G68), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT12), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n455), .B2(KEYINPUT11), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n450), .A2(new_n451), .A3(new_n456), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n449), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n447), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT72), .B1(new_n463), .B2(new_n335), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT72), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n462), .A2(new_n465), .A3(G190), .A4(new_n447), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n456), .A2(new_n451), .A3(new_n459), .ZN(new_n469));
  OAI21_X1  g0269(.A(G169), .B1(new_n448), .B2(new_n449), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n470), .A2(KEYINPUT14), .B1(new_n463), .B2(new_n381), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT14), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n463), .B2(G169), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G20), .A2(G77), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT15), .B(G87), .ZN(new_n477));
  OAI221_X1 g0277(.A(new_n476), .B1(new_n477), .B2(new_n337), .C1(new_n344), .C2(new_n339), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n257), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n479), .B(KEYINPUT69), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n228), .B2(new_n346), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n273), .A2(G77), .A3(new_n274), .A4(new_n349), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n318), .A2(new_n223), .B1(new_n230), .B2(new_n315), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n304), .A2(new_n382), .A3(G1698), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n321), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n445), .B1(G244), .B2(new_n377), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G179), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n361), .B2(new_n488), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(G200), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n335), .B2(new_n488), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n483), .B2(new_n493), .ZN(new_n494));
  NOR4_X1   g0294(.A1(new_n364), .A2(new_n438), .A3(new_n475), .A4(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT21), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n265), .A2(new_n266), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n268), .A2(new_n258), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n497), .A2(new_n277), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(G169), .B1(new_n293), .B2(new_n306), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n269), .B2(new_n277), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT21), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n293), .A2(new_n306), .A3(new_n381), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n278), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n405), .A2(new_n407), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n406), .B1(new_n315), .B2(G20), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n230), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT6), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n511), .A2(new_n440), .A3(G107), .ZN(new_n512));
  XNOR2_X1  g0312(.A(G97), .B(G107), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n514), .A2(new_n206), .B1(new_n228), .B2(new_n344), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n257), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n270), .A2(G97), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n271), .A2(new_n275), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(G97), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n315), .A2(KEYINPUT4), .A3(G244), .A4(new_n316), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n315), .A2(G250), .A3(G1698), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n229), .A2(G1698), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n419), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n294), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G257), .B(new_n280), .C1(new_n284), .C2(new_n286), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n292), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G190), .ZN(new_n533));
  INV_X1    g0333(.A(new_n531), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT4), .B1(new_n298), .B2(new_n526), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n321), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n520), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G264), .B(new_n280), .C1(new_n284), .C2(new_n286), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G250), .A2(G1698), .ZN(new_n542));
  INV_X1    g0342(.A(G257), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(G1698), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n298), .A2(new_n544), .B1(G33), .B2(G294), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n541), .B(new_n292), .C1(new_n545), .C2(new_n294), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n433), .ZN(new_n547));
  INV_X1    g0347(.A(new_n544), .ZN(new_n548));
  INV_X1    g0348(.A(G294), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n419), .A2(new_n548), .B1(new_n259), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n321), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n551), .A2(new_n335), .A3(new_n292), .A4(new_n541), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n224), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n371), .A2(new_n206), .A3(new_n295), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n206), .A2(G87), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n554), .B1(new_n304), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G116), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(G20), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT23), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n206), .B2(G107), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n230), .A2(KEYINPUT23), .A3(G20), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n556), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT24), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT24), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n556), .A2(new_n558), .A3(new_n567), .A4(new_n564), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n397), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n270), .A2(G107), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n570), .B(KEYINPUT25), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n397), .A2(new_n270), .A3(new_n276), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(new_n230), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n553), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n516), .A2(new_n519), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n361), .B1(new_n529), .B2(new_n531), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n534), .A2(new_n381), .A3(new_n537), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n540), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n546), .A2(new_n361), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n551), .A2(new_n381), .A3(new_n292), .A4(new_n541), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n582), .C1(new_n569), .C2(new_n573), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n225), .B1(new_n323), .B2(G1), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n205), .A2(new_n289), .A3(G45), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n280), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(G238), .A2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n229), .B2(G1698), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n298), .A2(new_n588), .B1(G33), .B2(G116), .ZN(new_n589));
  OAI211_X1 g0389(.A(G190), .B(new_n586), .C1(new_n589), .C2(new_n294), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n371), .A3(new_n295), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n294), .B1(new_n591), .B2(new_n559), .ZN(new_n592));
  INV_X1    g0392(.A(new_n586), .ZN(new_n593));
  OAI21_X1  g0393(.A(G200), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n595));
  AOI21_X1  g0395(.A(G20), .B1(G33), .B2(G97), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT19), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT19), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(new_n206), .A3(G33), .A4(G97), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n371), .A2(new_n206), .A3(G68), .A4(new_n295), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(new_n257), .B1(new_n346), .B2(new_n477), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n348), .A2(G87), .A3(new_n276), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n590), .A2(new_n594), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n477), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n518), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n603), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n586), .B1(new_n589), .B2(new_n294), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n361), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n592), .A2(new_n593), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n381), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n583), .A2(new_n605), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n580), .A2(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n314), .A2(new_n495), .A3(new_n507), .A4(new_n615), .ZN(G372));
  AND3_X1   g0416(.A1(new_n540), .A2(new_n575), .A3(new_n579), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT82), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n608), .A2(new_n610), .A3(new_n612), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n590), .A2(new_n594), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n603), .A2(new_n604), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT81), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n603), .A2(new_n604), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n617), .A2(new_n618), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n624), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n623), .B1(new_n603), .B2(new_n604), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n620), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n613), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT82), .B1(new_n580), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n502), .A2(KEYINPUT21), .B1(new_n278), .B2(new_n504), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n501), .A3(new_n583), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n627), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n576), .A2(new_n578), .A3(new_n577), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n630), .A3(new_n613), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(KEYINPUT26), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n613), .A2(new_n605), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n579), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n613), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n635), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n495), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n363), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n421), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n415), .A2(new_n206), .B1(new_n402), .B2(new_n344), .ZN(new_n648));
  INV_X1    g0448(.A(new_n303), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n368), .A2(new_n370), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(new_n259), .ZN(new_n651));
  INV_X1    g0451(.A(new_n407), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n509), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n648), .B1(new_n653), .B2(G68), .ZN(new_n654));
  INV_X1    g0454(.A(new_n411), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n257), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n392), .B1(new_n647), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n386), .A2(new_n388), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n491), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n470), .A2(KEYINPUT14), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n463), .A2(new_n472), .A3(G169), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n664), .B(new_n665), .C1(new_n381), .C2(new_n463), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n468), .A2(new_n663), .B1(new_n469), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n437), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n358), .A2(new_n359), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n646), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n645), .A2(new_n671), .ZN(G369));
  INV_X1    g0472(.A(KEYINPUT85), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n506), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n268), .A2(new_n206), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n278), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT84), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n314), .A2(KEYINPUT85), .A3(new_n501), .A4(new_n633), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n675), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n507), .A2(new_n683), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n681), .B1(new_n569), .B2(new_n573), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n575), .A2(new_n583), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT86), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT86), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n575), .A2(new_n691), .A3(new_n583), .A4(new_n688), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n583), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n681), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n687), .A2(G330), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n681), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n690), .A2(new_n506), .A3(new_n698), .A4(new_n692), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n209), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(G116), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n595), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n703), .A2(new_n705), .A3(new_n205), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n219), .B2(new_n703), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  AOI21_X1  g0508(.A(new_n641), .B1(new_n626), .B2(new_n636), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n538), .A2(new_n361), .B1(new_n516), .B2(new_n519), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n578), .A3(new_n605), .A4(new_n613), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n613), .B1(new_n711), .B2(KEYINPUT26), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT89), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n634), .A2(new_n617), .A3(new_n626), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n619), .B1(new_n640), .B2(new_n641), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n637), .A2(KEYINPUT26), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT89), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n713), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(KEYINPUT90), .A3(new_n698), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT90), .B1(new_n719), .B2(new_n698), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT29), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n681), .B1(new_n635), .B2(new_n643), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(KEYINPUT29), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n532), .A2(new_n504), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n541), .B1(new_n545), .B2(new_n294), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT87), .B1(new_n727), .B2(new_n609), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT87), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n611), .A2(new_n729), .A3(new_n541), .A4(new_n551), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n310), .A2(G179), .A3(new_n611), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n546), .A3(new_n538), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n728), .A2(new_n504), .A3(new_n532), .A4(new_n730), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n731), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT88), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n615), .A2(new_n507), .A3(new_n314), .A4(new_n698), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n737), .A2(new_n681), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n737), .A2(KEYINPUT88), .A3(KEYINPUT31), .A4(new_n681), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n740), .A2(new_n741), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n722), .A2(new_n725), .B1(G330), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n708), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n267), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n205), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n703), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n702), .A2(new_n298), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n323), .B2(new_n219), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n323), .B2(new_n253), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n702), .A2(new_n304), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n757), .A2(G355), .B1(new_n704), .B2(new_n702), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n756), .A2(KEYINPUT91), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n216), .B1(G20), .B2(new_n361), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT91), .B1(new_n756), .B2(new_n758), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n752), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n760), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n206), .B1(new_n769), .B2(G190), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n440), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n206), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n769), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G159), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n771), .B1(new_n775), .B2(KEYINPUT32), .ZN(new_n776));
  NAND3_X1  g0576(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT93), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n335), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n776), .B1(KEYINPUT32), .B2(new_n775), .C1(new_n780), .C2(new_n248), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(G190), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(G68), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n206), .A2(new_n335), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n381), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G58), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n772), .A2(new_n785), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n228), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT92), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n433), .A2(G179), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n772), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n230), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n784), .A2(new_n793), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n315), .B1(new_n796), .B2(new_n224), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n791), .A2(new_n792), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n794), .ZN(new_n799));
  INV_X1    g0599(.A(new_n788), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G283), .A2(new_n799), .B1(new_n800), .B2(G311), .ZN(new_n801));
  INV_X1    g0601(.A(new_n796), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G303), .A2(new_n802), .B1(new_n774), .B2(G329), .ZN(new_n803));
  INV_X1    g0603(.A(new_n770), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G294), .ZN(new_n805));
  INV_X1    g0605(.A(new_n786), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n315), .B1(new_n806), .B2(G322), .ZN(new_n807));
  AND4_X1   g0607(.A1(new_n801), .A2(new_n803), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n779), .A2(G326), .ZN(new_n809));
  INV_X1    g0609(.A(new_n782), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT33), .B(G317), .Z(new_n811));
  OAI211_X1 g0611(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT94), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n783), .A2(new_n798), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n768), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n767), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n763), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n687), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G330), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n685), .B2(new_n686), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(new_n752), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n687), .A2(G330), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n819), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT95), .Z(G396));
  NAND2_X1  g0625(.A1(new_n663), .A2(new_n698), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n483), .A2(new_n493), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n698), .B1(new_n481), .B2(new_n482), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n491), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n723), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n746), .A2(G330), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n752), .B1(new_n831), .B2(new_n832), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n760), .A2(new_n761), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n752), .B1(new_n837), .B2(G77), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n224), .A2(new_n794), .B1(new_n788), .B2(new_n704), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n796), .A2(new_n230), .B1(new_n773), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n304), .B1(new_n786), .B2(new_n549), .ZN(new_n842));
  NOR4_X1   g0642(.A1(new_n839), .A2(new_n841), .A3(new_n842), .A4(new_n771), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  INV_X1    g0644(.A(G303), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n843), .B1(new_n844), .B2(new_n810), .C1(new_n845), .C2(new_n780), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n799), .A2(G68), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n248), .B2(new_n796), .C1(new_n848), .C2(new_n773), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n419), .B(new_n849), .C1(G58), .C2(new_n804), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n806), .B1(new_n800), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G137), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n810), .B2(new_n343), .C1(new_n852), .C2(new_n780), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT34), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n854), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n846), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n838), .B1(new_n858), .B2(new_n760), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n830), .B2(new_n762), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT96), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n835), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  NOR2_X1   g0663(.A1(new_n749), .A2(new_n205), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n741), .A2(new_n744), .A3(new_n738), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n460), .B1(new_n466), .B2(new_n464), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n469), .B(new_n681), .C1(new_n866), .C2(new_n666), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n469), .A2(new_n681), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n468), .A2(new_n474), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n865), .A2(new_n870), .A3(new_n830), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(KEYINPUT40), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT97), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n655), .B1(new_n417), .B2(new_n421), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n397), .ZN(new_n876));
  AOI21_X1  g0676(.A(G20), .B1(new_n371), .B2(new_n295), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n222), .B1(new_n877), .B2(new_n406), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n414), .A2(new_n416), .B1(new_n878), .B2(new_n418), .ZN(new_n879));
  OAI211_X1 g0679(.A(KEYINPUT97), .B(new_n257), .C1(new_n879), .C2(new_n655), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n422), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n392), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n386), .A2(new_n388), .A3(new_n679), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n873), .B1(new_n884), .B2(new_n436), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT98), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n390), .B2(new_n423), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n386), .A2(new_n388), .A3(KEYINPUT77), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT77), .B1(new_n386), .B2(new_n388), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(new_n657), .A3(KEYINPUT98), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT99), .B1(new_n423), .B2(new_n679), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT99), .ZN(new_n894));
  INV_X1    g0694(.A(new_n679), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n657), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n436), .A2(new_n873), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n892), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT100), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT100), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n892), .A2(new_n897), .A3(new_n898), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n885), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n882), .A2(new_n895), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n425), .B2(new_n437), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n885), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n436), .A2(new_n873), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n896), .B2(new_n893), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n901), .B1(new_n910), .B2(new_n892), .ZN(new_n911));
  AND4_X1   g0711(.A1(new_n901), .A2(new_n892), .A3(new_n897), .A4(new_n898), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n906), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n872), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n436), .A2(KEYINPUT101), .B1(new_n657), .B2(new_n658), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n897), .B(new_n917), .C1(KEYINPUT101), .C2(new_n436), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n900), .A2(new_n902), .B1(KEYINPUT37), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n897), .B1(new_n662), .B2(new_n437), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n904), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n913), .A2(KEYINPUT38), .A3(new_n914), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n871), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n916), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT103), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n495), .A2(new_n865), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(G330), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n926), .A2(new_n928), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n904), .B1(new_n903), .B2(new_n906), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n922), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n867), .A2(new_n869), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n644), .A2(new_n830), .A3(new_n698), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n937), .B2(new_n826), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n662), .B2(new_n895), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n921), .A2(new_n922), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT102), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n935), .A2(KEYINPUT39), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT102), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n921), .A2(new_n922), .A3(new_n945), .A4(new_n941), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n666), .A2(new_n469), .A3(new_n698), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n940), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n722), .A2(new_n495), .A3(new_n725), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n671), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n950), .B(new_n952), .Z(new_n953));
  AOI21_X1  g0753(.A(new_n864), .B1(new_n933), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n933), .ZN(new_n955));
  INV_X1    g0755(.A(new_n514), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT35), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT35), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n957), .A2(G116), .A3(new_n217), .A4(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT36), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n219), .A2(G77), .A3(new_n400), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n249), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(G1), .A3(new_n267), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n955), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT105), .Z(G367));
  INV_X1    g0765(.A(new_n752), .ZN(new_n966));
  INV_X1    g0766(.A(new_n764), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n702), .B2(new_n606), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n753), .A2(new_n243), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n626), .B1(new_n625), .B2(new_n698), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n619), .A2(new_n622), .A3(new_n624), .A4(new_n681), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n786), .A2(new_n343), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n770), .A2(new_n222), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n779), .C2(G143), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT113), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT113), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n782), .A2(G159), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n315), .B1(new_n796), .B2(new_n787), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n248), .A2(new_n788), .B1(new_n794), .B2(new_n228), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(G137), .C2(new_n774), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(G317), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n786), .A2(new_n845), .B1(new_n773), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n802), .A2(KEYINPUT46), .A3(G116), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n419), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n985), .B(new_n987), .C1(G97), .C2(new_n799), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n549), .B2(new_n810), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT46), .B1(new_n802), .B2(G116), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT112), .Z(new_n991));
  OAI22_X1  g0791(.A1(new_n788), .A2(new_n844), .B1(new_n770), .B2(new_n230), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT111), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(new_n840), .C2(new_n780), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n983), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT114), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  OAI221_X1 g0797(.A(new_n970), .B1(new_n818), .B2(new_n973), .C1(new_n997), .C2(new_n768), .ZN(new_n998));
  INV_X1    g0798(.A(new_n747), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n700), .A2(new_n699), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n540), .B(new_n579), .C1(new_n520), .C2(new_n698), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n636), .A2(new_n681), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1000), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1000), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n700), .A2(new_n699), .A3(new_n1004), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1004), .B1(new_n700), .B2(new_n699), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT108), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1009), .B(new_n697), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1013), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n697), .B1(new_n1023), .B2(new_n1009), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT109), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n507), .A2(new_n681), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n700), .B1(new_n696), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n821), .B(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1025), .A2(new_n1026), .A3(new_n747), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT29), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n719), .A2(new_n698), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT90), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n719), .A2(KEYINPUT90), .A3(new_n698), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n832), .B(new_n1029), .C1(new_n1036), .C2(new_n724), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1009), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n697), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n1018), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT109), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n999), .B1(new_n1030), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n703), .B(KEYINPUT41), .Z(new_n1044));
  OAI21_X1  g0844(.A(new_n750), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1005), .A2(new_n700), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(KEYINPUT42), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT106), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1002), .A2(new_n583), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n681), .B1(new_n1049), .B2(new_n579), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1046), .B2(KEYINPUT42), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n973), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT43), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1048), .A2(new_n1054), .A3(new_n1053), .A4(new_n1051), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n697), .A2(new_n1005), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n1045), .A2(KEYINPUT110), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT110), .B1(new_n1045), .B2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n998), .B1(new_n1062), .B2(new_n1063), .ZN(G387));
  NAND3_X1  g0864(.A1(new_n693), .A2(new_n695), .A3(new_n763), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n757), .A2(new_n705), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(G107), .B2(new_n209), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n240), .A2(new_n323), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n339), .A2(G50), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT50), .ZN(new_n1070));
  AOI211_X1 g0870(.A(G45), .B(new_n705), .C1(G68), .C2(G77), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n754), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1067), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n752), .B1(new_n1073), .B2(new_n967), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G159), .A2(new_n779), .B1(new_n782), .B2(new_n340), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n802), .A2(G77), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G50), .A2(new_n806), .B1(new_n800), .B2(G68), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n794), .A2(new_n440), .B1(new_n773), .B2(new_n343), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n770), .A2(new_n477), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1078), .A2(new_n419), .A3(new_n1079), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n786), .A2(new_n984), .B1(new_n788), .B2(new_n845), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT115), .Z(new_n1083));
  XOR2_X1   g0883(.A(KEYINPUT116), .B(G322), .Z(new_n1084));
  NAND2_X1  g0884(.A1(new_n779), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(new_n840), .C2(new_n810), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n796), .A2(new_n549), .B1(new_n770), .B2(new_n844), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT117), .B(KEYINPUT49), .Z(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G116), .A2(new_n799), .B1(new_n774), .B2(G326), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1092), .A2(new_n419), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1091), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1081), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1074), .B1(new_n1096), .B2(new_n760), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1029), .A2(new_n751), .B1(new_n1065), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1037), .A2(new_n703), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n747), .A2(new_n1029), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(G393));
  NAND2_X1  g0901(.A1(new_n1030), .A2(new_n1042), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n703), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1025), .A2(new_n751), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n764), .B1(new_n440), .B2(new_n209), .C1(new_n754), .C2(new_n247), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n752), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n315), .B(new_n795), .C1(G116), .C2(new_n804), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n782), .A2(G303), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n800), .A2(G294), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G283), .A2(new_n802), .B1(new_n774), .B2(new_n1084), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n779), .A2(G317), .B1(G311), .B2(new_n806), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT52), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n779), .A2(G150), .B1(G159), .B2(new_n806), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT51), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n782), .A2(G50), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G87), .A2(new_n799), .B1(new_n774), .B2(G143), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n802), .A2(G68), .B1(new_n800), .B2(new_n340), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n419), .B1(G77), .B2(new_n804), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1113), .A2(new_n1115), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1108), .B1(new_n1123), .B2(new_n760), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1004), .B2(new_n818), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1105), .A2(new_n1106), .A3(new_n1125), .ZN(G390));
  AOI22_X1  g0926(.A1(new_n723), .A2(new_n829), .B1(new_n663), .B2(new_n698), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n948), .B1(new_n1127), .B2(new_n936), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n943), .A2(new_n944), .A3(new_n946), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n949), .B1(new_n921), .B2(new_n922), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1034), .A2(new_n1035), .A3(new_n826), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n829), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1132), .B2(new_n936), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n865), .A2(G330), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(new_n830), .A3(new_n870), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n746), .A2(G330), .A3(new_n830), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1139), .A2(new_n936), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1129), .A2(new_n1133), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n752), .B1(new_n837), .B2(new_n340), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n304), .B1(new_n770), .B2(new_n228), .C1(new_n224), .C2(new_n796), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n847), .B1(new_n704), .B2(new_n786), .C1(new_n549), .C2(new_n773), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(G283), .C2(new_n779), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n810), .A2(new_n230), .B1(new_n440), .B2(new_n788), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT121), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1152), .A2(KEYINPUT122), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G128), .A2(new_n779), .B1(new_n782), .B2(G137), .ZN(new_n1154));
  INV_X1    g0954(.A(G125), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n786), .A2(new_n848), .B1(new_n773), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n800), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n796), .A2(new_n343), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n315), .B1(new_n794), .B2(new_n248), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G159), .B2(new_n804), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1154), .A2(new_n1159), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1152), .A2(KEYINPUT122), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1153), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1144), .B1(new_n1166), .B2(new_n760), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n947), .B2(new_n762), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT123), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1143), .A2(new_n750), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1127), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1139), .A2(KEYINPUT118), .A3(new_n936), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1136), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT118), .B1(new_n1139), .B2(new_n936), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1175), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n865), .A2(new_n830), .A3(G330), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT119), .B1(new_n1180), .B2(new_n936), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1140), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(KEYINPUT119), .A3(new_n936), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n1132), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n495), .A2(new_n1135), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n951), .A2(new_n671), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1103), .B1(new_n1143), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1138), .A2(new_n1142), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1174), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1129), .A2(new_n1133), .A3(new_n1141), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1136), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1189), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AND4_X1   g0996(.A1(new_n1174), .A2(new_n1196), .A3(new_n1192), .A4(new_n703), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1173), .B1(new_n1193), .B2(new_n1197), .ZN(G378));
  AOI21_X1  g0998(.A(new_n679), .B1(new_n347), .B2(new_n350), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n364), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n364), .A2(new_n1199), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n925), .A2(G330), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n925), .B2(G330), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n941), .B1(new_n934), .B2(new_n922), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n921), .A2(new_n922), .A3(new_n941), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n945), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n948), .B1(new_n1212), .B2(new_n943), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1208), .A2(new_n1209), .B1(new_n1213), .B2(new_n940), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1207), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n871), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n920), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n911), .B2(new_n912), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT38), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1216), .B1(new_n1220), .B2(new_n907), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1221), .A2(KEYINPUT40), .B1(new_n935), .B2(new_n872), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1215), .B1(new_n1222), .B2(new_n820), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n925), .A2(G330), .A3(new_n1207), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n950), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1214), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1215), .A2(new_n761), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n298), .A2(G41), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G50), .B(new_n1228), .C1(new_n259), .C2(new_n281), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n806), .A2(G107), .B1(new_n800), .B2(new_n606), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n844), .B2(new_n773), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n794), .A2(new_n787), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n975), .B(new_n1233), .C1(G77), .C2(new_n802), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G97), .A2(new_n782), .B1(new_n779), .B2(G116), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1234), .A3(new_n1228), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT58), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1229), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n788), .A2(new_n852), .ZN(new_n1239));
  INV_X1    g1039(.A(G128), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1240), .A2(new_n786), .B1(new_n796), .B2(new_n1157), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1239), .B(new_n1241), .C1(G150), .C2(new_n804), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n1155), .B2(new_n780), .C1(new_n848), .C2(new_n810), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n259), .B(new_n281), .C1(new_n794), .C2(new_n402), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G124), .B2(new_n774), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1238), .B1(new_n1237), .B2(new_n1236), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n760), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT124), .Z(new_n1251));
  AOI211_X1 g1051(.A(new_n966), .B(new_n1251), .C1(new_n248), .C2(new_n836), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1226), .A2(new_n751), .B1(new_n1227), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT57), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1214), .B2(new_n1225), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1192), .A2(new_n1188), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n703), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT57), .B1(new_n1256), .B2(new_n1226), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1253), .B1(new_n1258), .B2(new_n1259), .ZN(G375));
  INV_X1    g1060(.A(new_n1044), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1187), .A2(new_n1179), .A3(new_n1184), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1189), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n936), .A2(new_n761), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n752), .B1(new_n837), .B2(G68), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n440), .A2(new_n796), .B1(new_n786), .B2(new_n844), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n788), .A2(new_n230), .B1(new_n773), .B2(new_n845), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n304), .B1(new_n794), .B2(new_n228), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .A4(new_n1079), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n1269), .B1(new_n704), .B2(new_n810), .C1(new_n549), .C2(new_n780), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n419), .B(new_n1233), .C1(G150), .C2(new_n800), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n796), .A2(new_n402), .B1(new_n773), .B2(new_n1240), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G137), .B2(new_n806), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1271), .B(new_n1273), .C1(new_n248), .C2(new_n770), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n848), .A2(new_n780), .B1(new_n810), .B2(new_n1157), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1270), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(KEYINPUT125), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n768), .B1(new_n1276), .B2(KEYINPUT125), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1265), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1185), .A2(new_n751), .B1(new_n1264), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1263), .A2(new_n1280), .ZN(G381));
  OR4_X1    g1081(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1172), .B1(new_n1192), .B2(new_n1190), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1282), .A2(new_n1284), .A3(G381), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1045), .A2(new_n1061), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT110), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1045), .A2(new_n1061), .A3(KEYINPUT110), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n950), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n947), .A2(new_n949), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n940), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1223), .A2(new_n1224), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n751), .B1(new_n1291), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1227), .A2(new_n1252), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1187), .B1(new_n1298), .B2(new_n1185), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1254), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1103), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1297), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1285), .A2(new_n1290), .A3(new_n998), .A4(new_n1303), .ZN(G407));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n680), .A3(new_n1283), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(G407), .A2(G213), .A3(new_n1305), .ZN(G409));
  NAND3_X1  g1106(.A1(new_n1256), .A2(new_n1261), .A3(new_n1226), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1253), .A2(new_n1307), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1303), .A2(G378), .B1(new_n1283), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  INV_X1    g1110(.A(G213), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(G343), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1189), .A2(KEYINPUT60), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1262), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1187), .A2(new_n1179), .A3(new_n1184), .A4(KEYINPUT60), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n703), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(G384), .A3(new_n1280), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1316), .B1(new_n1313), .B2(new_n1262), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1280), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n862), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1319), .A2(new_n1322), .ZN(new_n1323));
  NOR4_X1   g1123(.A1(new_n1309), .A2(new_n1310), .A3(new_n1312), .A4(new_n1323), .ZN(new_n1324));
  XOR2_X1   g1124(.A(G393), .B(G396), .Z(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(G390), .B1(new_n1290), .B2(new_n998), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n998), .B(G390), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1326), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  INV_X1    g1131(.A(G390), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G387), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1333), .A2(new_n1325), .A3(new_n1328), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1330), .A2(new_n1331), .A3(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1324), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1303), .A2(G378), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1308), .A2(new_n1283), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1312), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1312), .A2(G2897), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1323), .B(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(KEYINPUT126), .B1(new_n1339), .B2(new_n1342), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1323), .B(new_n1340), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1344), .B(new_n1345), .C1(new_n1312), .C2(new_n1309), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1343), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1323), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1339), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1310), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1336), .A2(new_n1347), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1330), .A2(new_n1334), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1344), .B1(new_n1309), .B2(new_n1312), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1190), .A2(new_n1174), .A3(new_n1192), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1196), .A2(new_n1192), .A3(new_n703), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(KEYINPUT120), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1172), .B1(new_n1354), .B2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1338), .B1(G375), .B2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1312), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1358), .A2(new_n1359), .A3(new_n1360), .A4(new_n1348), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1353), .A2(new_n1361), .A3(new_n1331), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1359), .B1(new_n1339), .B2(new_n1348), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1352), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1351), .A2(new_n1364), .ZN(G405));
  INV_X1    g1165(.A(new_n1352), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(G375), .A2(new_n1283), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1348), .A2(KEYINPUT127), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1367), .A2(new_n1368), .A3(new_n1337), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT127), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1369), .A2(new_n1370), .A3(new_n1323), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1323), .A2(new_n1370), .ZN(new_n1372));
  NAND4_X1  g1172(.A1(new_n1367), .A2(new_n1368), .A3(new_n1337), .A4(new_n1372), .ZN(new_n1373));
  AND3_X1   g1173(.A1(new_n1366), .A2(new_n1371), .A3(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1366), .B1(new_n1371), .B2(new_n1373), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1374), .A2(new_n1375), .ZN(G402));
endmodule


