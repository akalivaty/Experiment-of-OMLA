

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U555 ( .A1(n615), .A2(n614), .ZN(n678) );
  AND2_X1 U556 ( .A1(n528), .A2(G2104), .ZN(n898) );
  OR2_X1 U557 ( .A1(n678), .A2(n618), .ZN(n620) );
  NOR2_X1 U558 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  NOR2_X1 U560 ( .A1(n748), .A2(n747), .ZN(n749) );
  AND2_X1 U561 ( .A1(n531), .A2(n521), .ZN(G164) );
  XNOR2_X1 U562 ( .A(n525), .B(KEYINPUT87), .ZN(n531) );
  XNOR2_X2 U563 ( .A(n527), .B(n526), .ZN(n608) );
  XOR2_X2 U564 ( .A(KEYINPUT64), .B(n522), .Z(n895) );
  AND2_X1 U565 ( .A1(n530), .A2(n529), .ZN(n521) );
  XNOR2_X1 U566 ( .A(n669), .B(KEYINPUT30), .ZN(n670) );
  XNOR2_X1 U567 ( .A(n671), .B(n670), .ZN(n672) );
  INV_X1 U568 ( .A(KEYINPUT32), .ZN(n689) );
  NAND2_X1 U569 ( .A1(n612), .A2(n768), .ZN(n613) );
  NOR2_X1 U570 ( .A1(G2104), .A2(n528), .ZN(n894) );
  NOR2_X1 U571 ( .A1(G651), .A2(n575), .ZN(n796) );
  XNOR2_X1 U572 ( .A(n764), .B(KEYINPUT40), .ZN(n765) );
  INV_X1 U573 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U574 ( .A1(G126), .A2(n894), .ZN(n524) );
  NAND2_X1 U575 ( .A1(G114), .A2(n895), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U577 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n527) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  NAND2_X1 U579 ( .A1(G138), .A2(n608), .ZN(n530) );
  NAND2_X1 U580 ( .A1(G102), .A2(n898), .ZN(n529) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n575) );
  NAND2_X1 U582 ( .A1(n796), .A2(G52), .ZN(n534) );
  XOR2_X1 U583 ( .A(KEYINPUT68), .B(G651), .Z(n535) );
  NOR2_X1 U584 ( .A1(G543), .A2(n535), .ZN(n532) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n532), .Z(n621) );
  BUF_X1 U586 ( .A(n621), .Z(n793) );
  NAND2_X1 U587 ( .A1(G64), .A2(n793), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n541) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n792) );
  NAND2_X1 U590 ( .A1(G90), .A2(n792), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n575), .A2(n535), .ZN(n797) );
  NAND2_X1 U592 ( .A1(G77), .A2(n797), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U594 ( .A(KEYINPUT71), .B(n538), .ZN(n539) );
  XNOR2_X1 U595 ( .A(KEYINPUT9), .B(n539), .ZN(n540) );
  NOR2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U597 ( .A(KEYINPUT72), .B(n542), .Z(G301) );
  INV_X1 U598 ( .A(G301), .ZN(G171) );
  NAND2_X1 U599 ( .A1(G53), .A2(n796), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT74), .B(n543), .Z(n548) );
  NAND2_X1 U601 ( .A1(G91), .A2(n792), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G78), .A2(n797), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U604 ( .A(KEYINPUT73), .B(n546), .Z(n547) );
  NOR2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G65), .A2(n793), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(G299) );
  NAND2_X1 U608 ( .A1(n796), .A2(G51), .ZN(n551) );
  XOR2_X1 U609 ( .A(KEYINPUT77), .B(n551), .Z(n553) );
  NAND2_X1 U610 ( .A1(G63), .A2(n793), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U612 ( .A(KEYINPUT6), .B(n554), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G89), .A2(n792), .ZN(n555) );
  XNOR2_X1 U614 ( .A(n555), .B(KEYINPUT4), .ZN(n556) );
  XNOR2_X1 U615 ( .A(n556), .B(KEYINPUT76), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G76), .A2(n797), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U618 ( .A(n559), .B(KEYINPUT5), .Z(n560) );
  NOR2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U620 ( .A(KEYINPUT7), .B(n562), .Z(n563) );
  XNOR2_X1 U621 ( .A(KEYINPUT78), .B(n563), .ZN(G168) );
  NAND2_X1 U622 ( .A1(G88), .A2(n792), .ZN(n565) );
  NAND2_X1 U623 ( .A1(G50), .A2(n796), .ZN(n564) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n797), .A2(G75), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT82), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G62), .A2(n793), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U629 ( .A1(n570), .A2(n569), .ZN(G166) );
  INV_X1 U630 ( .A(G166), .ZN(G303) );
  XOR2_X1 U631 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U632 ( .A1(G49), .A2(n796), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U635 ( .A1(n793), .A2(n573), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT79), .B(n574), .Z(n577) );
  NAND2_X1 U637 ( .A1(n575), .A2(G87), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n577), .A2(n576), .ZN(G288) );
  NAND2_X1 U639 ( .A1(n792), .A2(G86), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G61), .A2(n793), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U642 ( .A(KEYINPUT80), .B(n580), .ZN(n584) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n582) );
  NAND2_X1 U644 ( .A1(n797), .A2(G73), .ZN(n581) );
  XOR2_X1 U645 ( .A(n582), .B(n581), .Z(n583) );
  NOR2_X1 U646 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n796), .A2(G48), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(G305) );
  NAND2_X1 U649 ( .A1(n793), .A2(G60), .ZN(n587) );
  XNOR2_X1 U650 ( .A(n587), .B(KEYINPUT70), .ZN(n590) );
  NAND2_X1 U651 ( .A1(G85), .A2(n792), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT67), .B(n588), .Z(n589) );
  NAND2_X1 U653 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U654 ( .A1(G72), .A2(n797), .ZN(n591) );
  XNOR2_X1 U655 ( .A(KEYINPUT69), .B(n591), .ZN(n592) );
  NOR2_X1 U656 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U657 ( .A1(n796), .A2(G47), .ZN(n594) );
  NAND2_X1 U658 ( .A1(n595), .A2(n594), .ZN(G290) );
  XNOR2_X1 U659 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  NAND2_X1 U660 ( .A1(G140), .A2(n608), .ZN(n597) );
  NAND2_X1 U661 ( .A1(G104), .A2(n898), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U663 ( .A(KEYINPUT34), .B(n598), .ZN(n604) );
  NAND2_X1 U664 ( .A1(G128), .A2(n894), .ZN(n600) );
  NAND2_X1 U665 ( .A1(G116), .A2(n895), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U667 ( .A(KEYINPUT35), .B(n601), .ZN(n602) );
  XNOR2_X1 U668 ( .A(KEYINPUT89), .B(n602), .ZN(n603) );
  NOR2_X1 U669 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U670 ( .A(KEYINPUT36), .B(n605), .ZN(n907) );
  NOR2_X1 U671 ( .A1(n758), .A2(n907), .ZN(n930) );
  NOR2_X1 U672 ( .A1(G164), .A2(G1384), .ZN(n615) );
  NAND2_X1 U673 ( .A1(G101), .A2(n898), .ZN(n606) );
  XOR2_X1 U674 ( .A(KEYINPUT23), .B(n606), .Z(n770) );
  AND2_X1 U675 ( .A1(n770), .A2(G40), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n894), .A2(G125), .ZN(n767) );
  AND2_X1 U677 ( .A1(n607), .A2(n767), .ZN(n612) );
  NAND2_X1 U678 ( .A1(n608), .A2(G137), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G113), .A2(n895), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U681 ( .A(KEYINPUT66), .B(n611), .Z(n768) );
  NOR2_X1 U682 ( .A1(n615), .A2(n613), .ZN(n760) );
  NAND2_X1 U683 ( .A1(n930), .A2(n760), .ZN(n756) );
  XOR2_X1 U684 ( .A(KEYINPUT92), .B(n613), .Z(n614) );
  XNOR2_X1 U685 ( .A(G2078), .B(KEYINPUT25), .ZN(n951) );
  NOR2_X1 U686 ( .A1(n678), .A2(n951), .ZN(n617) );
  AND2_X1 U687 ( .A1(n678), .A2(G1961), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n673) );
  NAND2_X1 U689 ( .A1(G171), .A2(n673), .ZN(n667) );
  INV_X1 U690 ( .A(KEYINPUT29), .ZN(n665) );
  INV_X1 U691 ( .A(G1996), .ZN(n618) );
  INV_X1 U692 ( .A(KEYINPUT26), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n620), .B(n619), .ZN(n633) );
  AND2_X1 U694 ( .A1(n678), .A2(G1341), .ZN(n631) );
  NAND2_X1 U695 ( .A1(n621), .A2(G56), .ZN(n622) );
  XOR2_X1 U696 ( .A(KEYINPUT14), .B(n622), .Z(n628) );
  NAND2_X1 U697 ( .A1(n792), .A2(G81), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(KEYINPUT12), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G68), .A2(n797), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U701 ( .A(KEYINPUT13), .B(n626), .Z(n627) );
  NOR2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n796), .A2(G43), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n972) );
  OR2_X1 U705 ( .A1(n631), .A2(n972), .ZN(n632) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n643) );
  NAND2_X1 U707 ( .A1(G54), .A2(n796), .ZN(n640) );
  NAND2_X1 U708 ( .A1(G66), .A2(n793), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G79), .A2(n797), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G92), .A2(n792), .ZN(n636) );
  XNOR2_X1 U712 ( .A(KEYINPUT75), .B(n636), .ZN(n637) );
  NOR2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(KEYINPUT15), .ZN(n973) );
  NOR2_X1 U716 ( .A1(n643), .A2(n973), .ZN(n642) );
  XOR2_X1 U717 ( .A(n642), .B(KEYINPUT96), .Z(n650) );
  NAND2_X1 U718 ( .A1(n643), .A2(n973), .ZN(n648) );
  NAND2_X1 U719 ( .A1(G1348), .A2(n678), .ZN(n645) );
  INV_X1 U720 ( .A(n678), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n653), .A2(G2067), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U723 ( .A(KEYINPUT95), .B(n646), .Z(n647) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(n657) );
  XOR2_X1 U726 ( .A(KEYINPUT93), .B(KEYINPUT27), .Z(n652) );
  NAND2_X1 U727 ( .A1(G2072), .A2(n653), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(n655) );
  INV_X1 U729 ( .A(G1956), .ZN(n981) );
  NOR2_X1 U730 ( .A1(n653), .A2(n981), .ZN(n654) );
  NOR2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n659) );
  INV_X1 U732 ( .A(G299), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n657), .A2(n656), .ZN(n663) );
  NOR2_X1 U735 ( .A1(n659), .A2(n658), .ZN(n661) );
  XOR2_X1 U736 ( .A(KEYINPUT28), .B(KEYINPUT94), .Z(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U738 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n667), .A2(n666), .ZN(n692) );
  NAND2_X1 U741 ( .A1(G8), .A2(n678), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n677), .A2(G1966), .ZN(n697) );
  NOR2_X1 U743 ( .A1(G2084), .A2(n678), .ZN(n693) );
  NOR2_X1 U744 ( .A1(n697), .A2(n693), .ZN(n668) );
  NAND2_X1 U745 ( .A1(n668), .A2(G8), .ZN(n671) );
  INV_X1 U746 ( .A(KEYINPUT97), .ZN(n669) );
  NOR2_X1 U747 ( .A1(n672), .A2(G168), .ZN(n675) );
  NOR2_X1 U748 ( .A1(n673), .A2(G171), .ZN(n674) );
  XOR2_X1 U749 ( .A(KEYINPUT31), .B(n676), .Z(n691) );
  INV_X1 U750 ( .A(G8), .ZN(n683) );
  NOR2_X1 U751 ( .A1(G1971), .A2(n677), .ZN(n680) );
  NOR2_X1 U752 ( .A1(G2090), .A2(n678), .ZN(n679) );
  NOR2_X1 U753 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U754 ( .A1(n681), .A2(G303), .ZN(n682) );
  OR2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n685) );
  AND2_X1 U756 ( .A1(n691), .A2(n685), .ZN(n684) );
  NAND2_X1 U757 ( .A1(n692), .A2(n684), .ZN(n688) );
  INV_X1 U758 ( .A(n685), .ZN(n686) );
  OR2_X1 U759 ( .A1(n686), .A2(G286), .ZN(n687) );
  NAND2_X1 U760 ( .A1(n688), .A2(n687), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n690), .B(n689), .ZN(n699) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U763 ( .A1(G8), .A2(n693), .ZN(n694) );
  NAND2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n714) );
  NOR2_X1 U767 ( .A1(G288), .A2(G1976), .ZN(n700) );
  XNOR2_X1 U768 ( .A(n700), .B(KEYINPUT98), .ZN(n987) );
  NOR2_X1 U769 ( .A1(G1971), .A2(G303), .ZN(n701) );
  XOR2_X1 U770 ( .A(n701), .B(KEYINPUT99), .Z(n702) );
  NOR2_X1 U771 ( .A1(n987), .A2(n702), .ZN(n703) );
  XOR2_X1 U772 ( .A(KEYINPUT100), .B(n703), .Z(n704) );
  NOR2_X1 U773 ( .A1(n714), .A2(n704), .ZN(n707) );
  NAND2_X1 U774 ( .A1(G1976), .A2(G288), .ZN(n985) );
  NOR2_X1 U775 ( .A1(KEYINPUT101), .A2(n677), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n985), .A2(n705), .ZN(n706) );
  NOR2_X1 U777 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U778 ( .A1(KEYINPUT33), .A2(n708), .ZN(n712) );
  XOR2_X1 U779 ( .A(n987), .B(KEYINPUT101), .Z(n709) );
  NAND2_X1 U780 ( .A1(n709), .A2(KEYINPUT33), .ZN(n710) );
  NOR2_X1 U781 ( .A1(n677), .A2(n710), .ZN(n711) );
  NOR2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U783 ( .A(G1981), .B(G305), .Z(n991) );
  NAND2_X1 U784 ( .A1(n713), .A2(n991), .ZN(n720) );
  INV_X1 U785 ( .A(n714), .ZN(n717) );
  NOR2_X1 U786 ( .A1(G2090), .A2(G303), .ZN(n715) );
  NAND2_X1 U787 ( .A1(G8), .A2(n715), .ZN(n716) );
  NAND2_X1 U788 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U789 ( .A1(n718), .A2(n677), .ZN(n719) );
  NAND2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U791 ( .A(n721), .B(KEYINPUT102), .ZN(n725) );
  NOR2_X1 U792 ( .A1(G1981), .A2(G305), .ZN(n722) );
  XOR2_X1 U793 ( .A(n722), .B(KEYINPUT24), .Z(n723) );
  NOR2_X1 U794 ( .A1(n677), .A2(n723), .ZN(n724) );
  NOR2_X1 U795 ( .A1(n725), .A2(n724), .ZN(n748) );
  NOR2_X1 U796 ( .A1(G1986), .A2(G290), .ZN(n751) );
  INV_X1 U797 ( .A(n751), .ZN(n984) );
  NAND2_X1 U798 ( .A1(G1986), .A2(G290), .ZN(n979) );
  NAND2_X1 U799 ( .A1(n984), .A2(n979), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n726), .A2(n760), .ZN(n727) );
  XNOR2_X1 U801 ( .A(n727), .B(KEYINPUT88), .ZN(n746) );
  NAND2_X1 U802 ( .A1(G119), .A2(n894), .ZN(n729) );
  NAND2_X1 U803 ( .A1(G95), .A2(n898), .ZN(n728) );
  NAND2_X1 U804 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U805 ( .A1(n895), .A2(G107), .ZN(n730) );
  XOR2_X1 U806 ( .A(KEYINPUT90), .B(n730), .Z(n731) );
  NOR2_X1 U807 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U808 ( .A1(n608), .A2(G131), .ZN(n733) );
  NAND2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n889) );
  NAND2_X1 U810 ( .A1(G1991), .A2(n889), .ZN(n744) );
  NAND2_X1 U811 ( .A1(G105), .A2(n898), .ZN(n735) );
  XOR2_X1 U812 ( .A(KEYINPUT38), .B(n735), .Z(n740) );
  NAND2_X1 U813 ( .A1(G129), .A2(n894), .ZN(n737) );
  NAND2_X1 U814 ( .A1(G117), .A2(n895), .ZN(n736) );
  NAND2_X1 U815 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U816 ( .A(KEYINPUT91), .B(n738), .Z(n739) );
  NOR2_X1 U817 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U818 ( .A1(n608), .A2(G141), .ZN(n741) );
  NAND2_X1 U819 ( .A1(n742), .A2(n741), .ZN(n885) );
  NAND2_X1 U820 ( .A1(G1996), .A2(n885), .ZN(n743) );
  NAND2_X1 U821 ( .A1(n744), .A2(n743), .ZN(n929) );
  NAND2_X1 U822 ( .A1(n929), .A2(n760), .ZN(n745) );
  NAND2_X1 U823 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U824 ( .A1(n756), .A2(n749), .ZN(n763) );
  NOR2_X1 U825 ( .A1(G1996), .A2(n885), .ZN(n750) );
  XOR2_X1 U826 ( .A(KEYINPUT103), .B(n750), .Z(n938) );
  NOR2_X1 U827 ( .A1(G1991), .A2(n889), .ZN(n928) );
  NOR2_X1 U828 ( .A1(n751), .A2(n928), .ZN(n752) );
  NOR2_X1 U829 ( .A1(n929), .A2(n752), .ZN(n753) );
  NOR2_X1 U830 ( .A1(n938), .A2(n753), .ZN(n754) );
  XNOR2_X1 U831 ( .A(n754), .B(KEYINPUT39), .ZN(n755) );
  XNOR2_X1 U832 ( .A(n755), .B(KEYINPUT104), .ZN(n757) );
  NAND2_X1 U833 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U834 ( .A1(n758), .A2(n907), .ZN(n945) );
  NAND2_X1 U835 ( .A1(n759), .A2(n945), .ZN(n761) );
  NAND2_X1 U836 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U837 ( .A1(n763), .A2(n762), .ZN(n766) );
  INV_X1 U838 ( .A(KEYINPUT105), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n766), .B(n765), .ZN(G329) );
  AND2_X1 U840 ( .A1(n768), .A2(n767), .ZN(n769) );
  AND2_X1 U841 ( .A1(n770), .A2(n769), .ZN(G160) );
  INV_X1 U842 ( .A(G96), .ZN(G221) );
  AND2_X1 U843 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U844 ( .A(G132), .ZN(G219) );
  INV_X1 U845 ( .A(G82), .ZN(G220) );
  INV_X1 U846 ( .A(G57), .ZN(G237) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n771) );
  XOR2_X1 U848 ( .A(n771), .B(KEYINPUT10), .Z(n922) );
  NAND2_X1 U849 ( .A1(n922), .A2(G567), .ZN(n772) );
  XOR2_X1 U850 ( .A(KEYINPUT11), .B(n772), .Z(G234) );
  INV_X1 U851 ( .A(G860), .ZN(n777) );
  OR2_X1 U852 ( .A1(n972), .A2(n777), .ZN(G153) );
  NAND2_X1 U853 ( .A1(G301), .A2(G868), .ZN(n774) );
  OR2_X1 U854 ( .A1(n973), .A2(G868), .ZN(n773) );
  NAND2_X1 U855 ( .A1(n774), .A2(n773), .ZN(G284) );
  NAND2_X1 U856 ( .A1(G868), .A2(G286), .ZN(n776) );
  INV_X1 U857 ( .A(G868), .ZN(n812) );
  NAND2_X1 U858 ( .A1(G299), .A2(n812), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n776), .A2(n775), .ZN(G297) );
  NAND2_X1 U860 ( .A1(n777), .A2(G559), .ZN(n778) );
  NAND2_X1 U861 ( .A1(n778), .A2(n973), .ZN(n779) );
  XNOR2_X1 U862 ( .A(n779), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U863 ( .A1(G868), .A2(n972), .ZN(n782) );
  NAND2_X1 U864 ( .A1(G868), .A2(n973), .ZN(n780) );
  NOR2_X1 U865 ( .A1(G559), .A2(n780), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(G282) );
  NAND2_X1 U867 ( .A1(n894), .A2(G123), .ZN(n783) );
  XNOR2_X1 U868 ( .A(n783), .B(KEYINPUT18), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G99), .A2(n898), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U871 ( .A1(n608), .A2(G135), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G111), .A2(n895), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n927) );
  XNOR2_X1 U875 ( .A(n927), .B(G2096), .ZN(n790) );
  INV_X1 U876 ( .A(G2100), .ZN(n858) );
  NAND2_X1 U877 ( .A1(n790), .A2(n858), .ZN(G156) );
  NAND2_X1 U878 ( .A1(n973), .A2(G559), .ZN(n809) );
  XNOR2_X1 U879 ( .A(n972), .B(n809), .ZN(n791) );
  NOR2_X1 U880 ( .A1(n791), .A2(G860), .ZN(n802) );
  NAND2_X1 U881 ( .A1(n792), .A2(G93), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G67), .A2(n793), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n801) );
  NAND2_X1 U884 ( .A1(n796), .A2(G55), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G80), .A2(n797), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n800) );
  OR2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n811) );
  XOR2_X1 U888 ( .A(n802), .B(n811), .Z(G145) );
  XOR2_X1 U889 ( .A(G299), .B(n972), .Z(n805) );
  XOR2_X1 U890 ( .A(KEYINPUT19), .B(n811), .Z(n803) );
  XNOR2_X1 U891 ( .A(n803), .B(G290), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n805), .B(n804), .ZN(n806) );
  XOR2_X1 U893 ( .A(G303), .B(n806), .Z(n807) );
  XNOR2_X1 U894 ( .A(n807), .B(G288), .ZN(n808) );
  XNOR2_X1 U895 ( .A(G305), .B(n808), .ZN(n910) );
  XNOR2_X1 U896 ( .A(n809), .B(n910), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n810), .A2(G868), .ZN(n814) );
  NAND2_X1 U898 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U899 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U900 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XOR2_X1 U901 ( .A(KEYINPUT20), .B(n815), .Z(n816) );
  NAND2_X1 U902 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U903 ( .A(n817), .B(KEYINPUT84), .ZN(n819) );
  XOR2_X1 U904 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n818) );
  XNOR2_X1 U905 ( .A(n819), .B(n818), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n820), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U908 ( .A1(G69), .A2(G120), .ZN(n821) );
  NOR2_X1 U909 ( .A1(G237), .A2(n821), .ZN(n822) );
  NAND2_X1 U910 ( .A1(G108), .A2(n822), .ZN(n845) );
  NAND2_X1 U911 ( .A1(G567), .A2(n845), .ZN(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT86), .B(n823), .Z(n829) );
  NOR2_X1 U913 ( .A1(G220), .A2(G219), .ZN(n824) );
  XOR2_X1 U914 ( .A(KEYINPUT22), .B(n824), .Z(n825) );
  NOR2_X1 U915 ( .A1(G218), .A2(n825), .ZN(n826) );
  XNOR2_X1 U916 ( .A(n826), .B(KEYINPUT85), .ZN(n827) );
  OR2_X1 U917 ( .A1(G221), .A2(n827), .ZN(n846) );
  AND2_X1 U918 ( .A1(n846), .A2(G2106), .ZN(n828) );
  NOR2_X1 U919 ( .A1(n829), .A2(n828), .ZN(G319) );
  INV_X1 U920 ( .A(G319), .ZN(n831) );
  NAND2_X1 U921 ( .A1(G661), .A2(G483), .ZN(n830) );
  NOR2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n844) );
  NAND2_X1 U923 ( .A1(n844), .A2(G36), .ZN(G176) );
  XNOR2_X1 U924 ( .A(G2454), .B(G2451), .ZN(n840) );
  XNOR2_X1 U925 ( .A(G2430), .B(G2446), .ZN(n838) );
  XOR2_X1 U926 ( .A(G2435), .B(G2427), .Z(n833) );
  XNOR2_X1 U927 ( .A(KEYINPUT106), .B(G2438), .ZN(n832) );
  XNOR2_X1 U928 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U929 ( .A(n834), .B(G2443), .Z(n836) );
  XNOR2_X1 U930 ( .A(G1341), .B(G1348), .ZN(n835) );
  XNOR2_X1 U931 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U932 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U933 ( .A(n840), .B(n839), .ZN(n841) );
  NAND2_X1 U934 ( .A1(n841), .A2(G14), .ZN(n917) );
  XNOR2_X1 U935 ( .A(KEYINPUT107), .B(n917), .ZN(G401) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n922), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n842) );
  NAND2_X1 U938 ( .A1(G661), .A2(n842), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U940 ( .A1(n844), .A2(n843), .ZN(G188) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  NOR2_X1 U944 ( .A1(n846), .A2(n845), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G1961), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1981), .B(G1966), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n849), .B(KEYINPUT111), .Z(n851) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U952 ( .A(G1986), .B(G1976), .Z(n853) );
  XOR2_X1 U953 ( .A(n981), .B(G1971), .Z(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U956 ( .A(G2474), .B(KEYINPUT110), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(G229) );
  XNOR2_X1 U958 ( .A(n858), .B(KEYINPUT109), .ZN(n860) );
  XNOR2_X1 U959 ( .A(G2678), .B(KEYINPUT43), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2067), .Z(n862) );
  XNOR2_X1 U962 ( .A(G2090), .B(G2072), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U965 ( .A(KEYINPUT108), .B(G2096), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n868) );
  XOR2_X1 U967 ( .A(G2078), .B(G2084), .Z(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(G227) );
  NAND2_X1 U969 ( .A1(n894), .A2(G124), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G100), .A2(n898), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n608), .A2(G136), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G112), .A2(n895), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U976 ( .A1(n875), .A2(n874), .ZN(G162) );
  NAND2_X1 U977 ( .A1(G139), .A2(n608), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G103), .A2(n898), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G115), .A2(n895), .ZN(n878) );
  XOR2_X1 U981 ( .A(KEYINPUT113), .B(n878), .Z(n880) );
  NAND2_X1 U982 ( .A1(n894), .A2(G127), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n923) );
  XOR2_X1 U986 ( .A(G164), .B(n923), .Z(n884) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n893) );
  XOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n887) );
  XNOR2_X1 U989 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U990 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U991 ( .A(G162), .B(n888), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n889), .B(n927), .ZN(n890) );
  XNOR2_X1 U993 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U994 ( .A(n893), .B(n892), .Z(n906) );
  NAND2_X1 U995 ( .A1(G130), .A2(n894), .ZN(n897) );
  NAND2_X1 U996 ( .A1(G118), .A2(n895), .ZN(n896) );
  NAND2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n903) );
  NAND2_X1 U998 ( .A1(G142), .A2(n608), .ZN(n900) );
  NAND2_X1 U999 ( .A1(G106), .A2(n898), .ZN(n899) );
  NAND2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1001 ( .A(KEYINPUT45), .B(n901), .Z(n902) );
  NOR2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(G160), .B(n904), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n908), .B(n907), .Z(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G395) );
  XNOR2_X1 U1007 ( .A(n910), .B(KEYINPUT115), .ZN(n912) );
  XOR2_X1 U1008 ( .A(G171), .B(n973), .Z(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n913), .B(G286), .Z(n914) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n917), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  INV_X1 U1021 ( .A(n922), .ZN(G223) );
  INV_X1 U1022 ( .A(KEYINPUT55), .ZN(n970) );
  XOR2_X1 U1023 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n948) );
  XOR2_X1 U1024 ( .A(G2072), .B(n923), .Z(n925) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n926), .Z(n944) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(G2084), .B(G160), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT117), .B(n933), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1034 ( .A(KEYINPUT118), .B(n936), .Z(n941) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(KEYINPUT51), .B(n939), .ZN(n940) );
  NOR2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(KEYINPUT119), .B(n942), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n948), .B(n947), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n970), .A2(n949), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1045 ( .A(G27), .B(n951), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(G1996), .B(G32), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G26), .B(G2067), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1050 ( .A(KEYINPUT121), .B(G2072), .Z(n956) );
  XNOR2_X1 U1051 ( .A(G33), .B(n956), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1053 ( .A(KEYINPUT122), .B(n959), .Z(n961) );
  XNOR2_X1 U1054 ( .A(G1991), .B(G25), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(G28), .A2(n962), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n963), .B(KEYINPUT53), .ZN(n966) );
  XOR2_X1 U1058 ( .A(G2084), .B(G34), .Z(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(n964), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(G35), .B(G2090), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n970), .B(n969), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(G29), .A2(n971), .ZN(n1027) );
  INV_X1 U1065 ( .A(G16), .ZN(n1023) );
  XOR2_X1 U1066 ( .A(n1023), .B(KEYINPUT56), .Z(n999) );
  XOR2_X1 U1067 ( .A(n972), .B(G1341), .Z(n976) );
  XOR2_X1 U1068 ( .A(n973), .B(KEYINPUT123), .Z(n974) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n974), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n978) );
  XOR2_X1 U1071 ( .A(G1961), .B(G171), .Z(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n997) );
  XOR2_X1 U1073 ( .A(G303), .B(G1971), .Z(n980) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n983) );
  XOR2_X1 U1075 ( .A(n981), .B(G299), .Z(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(KEYINPUT124), .B(n990), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1083 ( .A(KEYINPUT57), .B(n993), .Z(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1025) );
  XNOR2_X1 U1087 ( .A(G1966), .B(KEYINPUT126), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(G21), .ZN(n1007) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(G1986), .B(G24), .Z(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1018) );
  XOR2_X1 U1096 ( .A(G1981), .B(G6), .Z(n1009) );
  XOR2_X1 U1097 ( .A(G1956), .B(G20), .Z(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(G1341), .B(G19), .Z(n1013) );
  XOR2_X1 U1100 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n1010) );
  XNOR2_X1 U1101 ( .A(G4), .B(n1010), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(n1011), .B(G1348), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(n1016), .B(KEYINPUT60), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G5), .B(G1961), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(G11), .A2(n1028), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1117 ( .A(G150), .ZN(G311) );
endmodule

