//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  NOR2_X1   g0019(.A1(new_n209), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT0), .ZN(new_n222));
  INV_X1    g0022(.A(new_n201), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n207), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n222), .B(new_n228), .C1(new_n217), .C2(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n219), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G68), .ZN(new_n242));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n207), .A3(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n226), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n206), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n249), .A2(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n254), .A2(new_n256), .B1(G50), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n203), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g0065(.A(KEYINPUT8), .B(G58), .Z(new_n266));
  NAND2_X1  g0066(.A1(new_n207), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT67), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n265), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n252), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n260), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1698), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G222), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n277), .ZN(new_n281));
  INV_X1    g0081(.A(G223), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(G1698), .ZN(new_n283));
  OAI221_X1 g0083(.A(new_n279), .B1(new_n280), .B2(new_n281), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n226), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT66), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n285), .B2(new_n226), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(KEYINPUT66), .A3(G1), .A4(G13), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G226), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n293), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n289), .A2(new_n295), .A3(G274), .A4(new_n291), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n287), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G179), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  AOI211_X1 g0099(.A(new_n273), .B(new_n298), .C1(new_n299), .C2(new_n297), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n273), .A2(KEYINPUT9), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n272), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(new_n297), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G190), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT68), .B(G200), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n297), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n304), .A2(new_n305), .A3(new_n307), .A4(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n307), .A2(new_n310), .A3(new_n301), .A4(new_n303), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n300), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n289), .A2(G238), .A3(new_n293), .A4(new_n291), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G97), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  MUX2_X1   g0117(.A(G226), .B(G232), .S(G1698), .Z(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n281), .ZN(new_n319));
  INV_X1    g0119(.A(new_n286), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n296), .B(new_n315), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT74), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n328));
  INV_X1    g0128(.A(G179), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n326), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n324), .A3(new_n325), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT74), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n319), .A2(new_n320), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n335), .A2(new_n336), .A3(new_n296), .A4(new_n315), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n299), .B1(new_n337), .B2(new_n322), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT73), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT73), .B(KEYINPUT14), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n334), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n269), .A2(G77), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n243), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT72), .B1(new_n250), .B2(new_n243), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT12), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n253), .A2(G68), .A3(new_n255), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT11), .B1(new_n347), .B2(new_n252), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n344), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n337), .B2(new_n322), .ZN(new_n358));
  XOR2_X1   g0158(.A(new_n358), .B(KEYINPUT70), .Z(new_n359));
  INV_X1    g0159(.A(G190), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n328), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n355), .B1(new_n326), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n278), .A2(G232), .ZN(new_n364));
  INV_X1    g0164(.A(G107), .ZN(new_n365));
  INV_X1    g0165(.A(G238), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n364), .B1(new_n365), .B2(new_n281), .C1(new_n366), .C2(new_n283), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n286), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n292), .A2(G244), .A3(new_n293), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n369), .A2(new_n296), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n299), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n296), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n286), .B2(new_n367), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n372), .A2(KEYINPUT69), .B1(new_n329), .B2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT69), .A4(new_n329), .ZN(new_n376));
  INV_X1    g0176(.A(new_n266), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n377), .A2(new_n264), .B1(new_n207), .B2(new_n280), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n267), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n252), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n253), .A2(G77), .A3(new_n255), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n381), .B(new_n382), .C1(G77), .C2(new_n258), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n371), .A2(new_n309), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n374), .B2(G190), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n314), .A2(new_n356), .A3(new_n363), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT77), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n266), .A2(new_n255), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n253), .B1(new_n250), .B2(new_n377), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n276), .A2(new_n207), .A3(new_n277), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT75), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n277), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n398), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT75), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(G68), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G58), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n243), .ZN(new_n404));
  OAI21_X1  g0204(.A(G20), .B1(new_n404), .B2(new_n201), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n263), .A2(G159), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n396), .A2(new_n398), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n407), .B1(new_n412), .B2(G68), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n271), .B1(new_n413), .B2(KEYINPUT16), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n393), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n289), .A2(G232), .A3(new_n293), .A4(new_n291), .ZN(new_n416));
  INV_X1    g0216(.A(G87), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n275), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(G223), .A2(G1698), .ZN(new_n419));
  INV_X1    g0219(.A(G226), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(G1698), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n418), .B1(new_n421), .B2(new_n281), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n416), .B(new_n296), .C1(new_n422), .C2(new_n320), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n357), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(G1698), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G223), .B2(G1698), .ZN(new_n426));
  AND2_X1   g0226(.A1(KEYINPUT3), .A2(G33), .ZN(new_n427));
  NOR2_X1   g0227(.A1(KEYINPUT3), .A2(G33), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n426), .A2(new_n429), .B1(new_n275), .B2(new_n417), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n286), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n360), .A2(KEYINPUT76), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n360), .A2(KEYINPUT76), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n431), .A2(new_n416), .A3(new_n296), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n424), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT17), .B1(new_n415), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT16), .B1(new_n402), .B2(new_n408), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT7), .B1(new_n429), .B2(new_n207), .ZN(new_n439));
  OAI21_X1  g0239(.A(G68), .B1(new_n439), .B2(new_n400), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n252), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n392), .B(new_n436), .C1(new_n438), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n390), .B1(new_n437), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n392), .B1(new_n438), .B2(new_n442), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n423), .A2(G169), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n329), .B2(new_n423), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n448), .B1(new_n447), .B2(new_n450), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n415), .A2(KEYINPUT17), .A3(new_n436), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n443), .A2(new_n444), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(KEYINPUT77), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n446), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n389), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(G257), .B(G1698), .C1(new_n427), .C2(new_n428), .ZN(new_n459));
  INV_X1    g0259(.A(G1698), .ZN(new_n460));
  OAI211_X1 g0260(.A(G250), .B(new_n460), .C1(new_n427), .C2(new_n428), .ZN(new_n461));
  INV_X1    g0261(.A(G294), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n459), .B(new_n461), .C1(new_n275), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n286), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT86), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT86), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n466), .A3(new_n286), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n206), .A2(G45), .ZN(new_n468));
  OR2_X1    g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NAND2_X1  g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n471), .A2(G274), .A3(new_n289), .A4(new_n291), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  INV_X1    g0274(.A(new_n470), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n477), .A2(new_n289), .A3(G264), .A4(new_n291), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n465), .A2(new_n360), .A3(new_n467), .A4(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n464), .A2(new_n472), .A3(new_n478), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n357), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g0283(.A(KEYINPUT82), .B(KEYINPUT24), .Z(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT23), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(new_n365), .A3(G20), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n486), .A2(new_n488), .A3(new_n489), .A4(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n207), .B1(new_n427), .B2(new_n428), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n417), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n417), .B1(KEYINPUT81), .B2(KEYINPUT22), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n496), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n281), .A2(new_n499), .A3(new_n207), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n485), .B1(new_n494), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n491), .A2(new_n493), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(new_n484), .A3(new_n498), .A4(new_n501), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n252), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n207), .A2(G107), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n257), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(KEYINPUT84), .A3(KEYINPUT25), .ZN(new_n509));
  OR2_X1    g0309(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n510));
  NAND2_X1  g0310(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n257), .A2(new_n507), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n275), .A2(G1), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n250), .A2(new_n252), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n509), .B(new_n512), .C1(new_n515), .C2(new_n365), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n483), .A2(new_n506), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT85), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n504), .A2(new_n498), .A3(new_n501), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n271), .B1(new_n521), .B2(new_n485), .ZN(new_n522));
  AOI211_X1 g0322(.A(new_n520), .B(new_n516), .C1(new_n522), .C2(new_n505), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT85), .B1(new_n506), .B2(new_n517), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n465), .A2(new_n467), .A3(new_n479), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n526), .A2(new_n299), .B1(new_n329), .B2(new_n481), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n519), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n399), .A2(G107), .A3(new_n401), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  INV_X1    g0330(.A(G97), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n365), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n365), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n529), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n252), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT78), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT78), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n541), .A3(new_n252), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G283), .ZN(new_n544));
  OAI211_X1 g0344(.A(G250), .B(G1698), .C1(new_n427), .C2(new_n428), .ZN(new_n545));
  OAI211_X1 g0345(.A(G244), .B(new_n460), .C1(new_n427), .C2(new_n428), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT4), .B1(new_n278), .B2(G244), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n286), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n477), .A2(new_n289), .A3(G257), .A4(new_n291), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n472), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n357), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n552), .A3(G190), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT79), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n550), .A2(new_n552), .A3(KEYINPUT79), .A4(G190), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n258), .A2(G97), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n514), .B2(G97), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n543), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n541), .B1(new_n538), .B2(new_n252), .ZN(new_n562));
  AOI211_X1 g0362(.A(KEYINPUT78), .B(new_n271), .C1(new_n529), .C2(new_n537), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(G169), .B1(new_n550), .B2(new_n552), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n550), .A2(new_n552), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n565), .B1(new_n567), .B2(new_n329), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n281), .A2(G264), .A3(G1698), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n281), .A2(G257), .A3(new_n460), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n429), .A2(G303), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n286), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n292), .A2(G270), .A3(new_n477), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n472), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n514), .A2(G116), .ZN(new_n579));
  INV_X1    g0379(.A(G116), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n250), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n544), .B(new_n207), .C1(G33), .C2(new_n531), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(G20), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n252), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT20), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n579), .B(new_n581), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n578), .B(new_n589), .C1(new_n434), .C2(new_n577), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n577), .A2(G169), .A3(new_n588), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n577), .A2(new_n329), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n588), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n577), .A2(KEYINPUT21), .A3(G169), .A4(new_n588), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n590), .A2(new_n593), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(G244), .B(G1698), .C1(new_n427), .C2(new_n428), .ZN(new_n598));
  OAI211_X1 g0398(.A(G238), .B(new_n460), .C1(new_n427), .C2(new_n428), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G33), .A2(G116), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n286), .ZN(new_n602));
  AOI21_X1  g0402(.A(G250), .B1(new_n206), .B2(G45), .ZN(new_n603));
  INV_X1    g0403(.A(G274), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n604), .B2(new_n474), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n292), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n299), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n207), .B(G68), .C1(new_n427), .C2(new_n428), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n267), .B2(new_n531), .ZN(new_n611));
  AOI21_X1  g0411(.A(G20), .B1(new_n317), .B2(KEYINPUT19), .ZN(new_n612));
  NOR3_X1   g0412(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n609), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n252), .ZN(new_n615));
  INV_X1    g0415(.A(new_n379), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT80), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT80), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n379), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n514), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n379), .A2(new_n250), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n615), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n602), .A2(new_n606), .A3(new_n329), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n608), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n607), .A2(new_n360), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n614), .A2(new_n252), .B1(new_n250), .B2(new_n379), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n514), .A2(G87), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n286), .A2(new_n601), .B1(new_n292), .B2(new_n605), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n308), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n624), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n597), .A2(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n458), .A2(new_n528), .A3(new_n570), .A4(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n624), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n625), .B1(new_n629), .B2(KEYINPUT87), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(new_n627), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n308), .B1(new_n602), .B2(new_n606), .ZN(new_n636));
  OR3_X1    g0436(.A1(new_n635), .A2(new_n636), .A3(KEYINPUT87), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n561), .A2(new_n569), .A3(new_n638), .A4(new_n518), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n506), .A2(new_n517), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n527), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT26), .B1(new_n569), .B2(new_n630), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n638), .A2(new_n645), .A3(new_n564), .A4(new_n568), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n646), .A3(new_n624), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n458), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n363), .A2(new_n385), .B1(new_n344), .B2(new_n355), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n446), .A2(new_n456), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n453), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n311), .A2(new_n313), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n300), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(KEYINPUT91), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n257), .A2(new_n207), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n588), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT88), .Z(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n640), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n664), .A2(KEYINPUT89), .B1(new_n597), .B2(new_n663), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n664), .A2(KEYINPUT89), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g0468(.A(KEYINPUT90), .B(G330), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n655), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(KEYINPUT91), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n525), .ZN(new_n674));
  INV_X1    g0474(.A(new_n661), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n528), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n641), .A2(new_n520), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n506), .A2(KEYINPUT85), .A3(new_n517), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n527), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n676), .B1(new_n679), .B2(new_n675), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n640), .A2(new_n675), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n528), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n527), .A2(new_n641), .A3(new_n675), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n220), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n613), .A2(new_n580), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n689), .A2(new_n690), .A3(new_n206), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n225), .B2(new_n689), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT28), .Z(new_n693));
  AOI21_X1  g0493(.A(new_n640), .B1(new_n525), .B2(new_n527), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT94), .B1(new_n639), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n640), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n679), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT94), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n634), .A2(new_n637), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n699), .A2(new_n518), .A3(new_n624), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n570), .A2(new_n697), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n565), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(G179), .B2(new_n566), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n543), .B2(new_n560), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n645), .B1(new_n704), .B2(new_n638), .ZN(new_n705));
  AOI21_X1  g0505(.A(G169), .B1(new_n602), .B2(new_n606), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n329), .B2(new_n628), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n635), .A2(new_n636), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n628), .A2(G190), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n707), .A2(new_n622), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n564), .A3(new_n645), .A4(new_n568), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n624), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n695), .A2(new_n701), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n675), .B1(new_n643), .B2(new_n647), .ZN(new_n716));
  XNOR2_X1  g0516(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n628), .A2(new_n464), .A3(new_n478), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n594), .A2(new_n567), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT30), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n628), .A2(G179), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n577), .A3(new_n566), .A4(new_n481), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT92), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n675), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n570), .A2(new_n528), .A3(new_n631), .A4(new_n675), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n661), .A2(KEYINPUT31), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n722), .B2(new_n724), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n671), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n719), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n693), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(new_n689), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n249), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n206), .B1(new_n736), .B2(G45), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n739), .B(new_n673), .C1(new_n669), .C2(new_n668), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n688), .A2(new_n429), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n741), .A2(G355), .B1(new_n580), .B2(new_n688), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n688), .A2(new_n281), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G45), .B2(new_n224), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n247), .A2(new_n473), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT95), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n226), .B1(G20), .B2(new_n299), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n746), .B2(KEYINPUT95), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n738), .B1(new_n747), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n207), .A2(new_n329), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G190), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n207), .A2(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n757), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n281), .B(new_n760), .C1(G329), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n309), .A2(new_n761), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  INV_X1    g0568(.A(G303), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n765), .A2(new_n360), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n764), .B1(new_n767), .B2(new_n768), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n756), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n434), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G326), .ZN(new_n776));
  INV_X1    g0576(.A(new_n434), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n207), .A2(new_n329), .A3(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G322), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n775), .A2(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n773), .A2(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT33), .B(G317), .Z(new_n784));
  NOR3_X1   g0584(.A1(new_n360), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n207), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n783), .A2(new_n784), .B1(new_n462), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n772), .A2(new_n781), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n767), .A2(new_n365), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n429), .B(new_n789), .C1(G87), .C2(new_n770), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT96), .ZN(new_n791));
  INV_X1    g0591(.A(new_n779), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G58), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n762), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n796), .A2(KEYINPUT32), .B1(new_n782), .B2(G68), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n786), .A2(new_n531), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G50), .B2(new_n774), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT32), .ZN(new_n800));
  INV_X1    g0600(.A(new_n758), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n795), .A2(new_n800), .B1(new_n801), .B2(G77), .ZN(new_n802));
  AND4_X1   g0602(.A1(new_n793), .A2(new_n797), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n788), .B1(new_n791), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n751), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n755), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n668), .B2(new_n750), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n740), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  INV_X1    g0609(.A(KEYINPUT99), .ZN(new_n810));
  INV_X1    g0610(.A(new_n384), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n372), .A2(KEYINPUT69), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n371), .A2(G179), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n387), .A2(new_n386), .B1(new_n383), .B2(new_n661), .ZN(new_n815));
  OAI21_X1  g0615(.A(KEYINPUT99), .B1(new_n375), .B2(new_n384), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n675), .B(new_n817), .C1(new_n643), .C2(new_n647), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n817), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n385), .A2(new_n661), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n819), .B1(new_n716), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n731), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n739), .B1(new_n825), .B2(new_n731), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(new_n748), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n805), .A2(new_n749), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n739), .B1(G77), .B2(new_n830), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n779), .A2(new_n462), .B1(new_n783), .B2(new_n768), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n798), .B(new_n832), .C1(G303), .C2(new_n774), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n429), .B1(new_n762), .B2(new_n759), .C1(new_n580), .C2(new_n758), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(G87), .B2(new_n766), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n835), .C1(new_n365), .C2(new_n771), .ZN(new_n836));
  XNOR2_X1  g0636(.A(KEYINPUT97), .B(G143), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n792), .A2(new_n838), .B1(G137), .B2(new_n774), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n839), .B1(new_n262), .B2(new_n783), .C1(new_n794), .C2(new_n758), .ZN(new_n840));
  XNOR2_X1  g0640(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n281), .B1(new_n762), .B2(new_n843), .C1(new_n786), .C2(new_n403), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n767), .A2(new_n243), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n844), .B(new_n845), .C1(G50), .C2(new_n770), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n840), .A2(new_n841), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n836), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n831), .B1(new_n849), .B2(new_n751), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n827), .A2(new_n828), .B1(new_n829), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G384));
  OR2_X1    g0652(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n853), .A2(G116), .A3(new_n227), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT36), .Z(new_n856));
  OR3_X1    g0656(.A1(new_n224), .A2(new_n280), .A3(new_n404), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n206), .B(G13), .C1(new_n857), .C2(new_n242), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n715), .A2(new_n458), .A3(new_n718), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n653), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT103), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n814), .A2(new_n816), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n675), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n818), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n341), .B1(new_n338), .B2(new_n342), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n331), .B2(new_n333), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT100), .B1(new_n867), .B2(new_n354), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT100), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n344), .A2(new_n869), .A3(new_n355), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT101), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n354), .B2(new_n675), .ZN(new_n872));
  OAI211_X1 g0672(.A(KEYINPUT101), .B(new_n661), .C1(new_n352), .C2(new_n353), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n359), .B2(new_n362), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n868), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n363), .A2(new_n867), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n355), .A3(new_n661), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n865), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n447), .A2(new_n450), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n659), .B(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n447), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n882), .A2(new_n884), .A3(new_n885), .A4(new_n443), .ZN(new_n886));
  INV_X1    g0686(.A(new_n450), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n414), .B1(KEYINPUT16), .B2(new_n413), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n887), .A2(new_n659), .B1(new_n888), .B2(new_n392), .ZN(new_n889));
  INV_X1    g0689(.A(new_n443), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n659), .B1(new_n888), .B2(new_n392), .ZN(new_n892));
  AOI221_X4 g0692(.A(new_n881), .B1(new_n886), .B2(new_n891), .C1(new_n457), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n457), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n886), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n880), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n453), .A2(new_n883), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n896), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n882), .A2(KEYINPUT18), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n447), .A2(new_n450), .A3(new_n448), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n454), .A2(new_n455), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n447), .B(new_n883), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n882), .A2(new_n884), .A3(new_n443), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n886), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n881), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n902), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n661), .B1(new_n868), .B2(new_n870), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n903), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n900), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n862), .B(new_n919), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n876), .A2(new_n878), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n823), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n726), .A2(KEYINPUT31), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n728), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n922), .A2(KEYINPUT40), .A3(new_n914), .A4(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n879), .B(new_n822), .C1(new_n728), .C2(new_n923), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(new_n897), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n924), .A2(new_n458), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n931), .A2(new_n932), .A3(new_n669), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n920), .A2(new_n933), .B1(new_n206), .B2(new_n736), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n920), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n859), .B1(new_n934), .B2(new_n935), .ZN(G367));
  NAND2_X1  g0736(.A1(new_n743), .A2(new_n237), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n753), .B1(new_n688), .B2(new_n616), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n738), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n750), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n635), .A2(new_n661), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n638), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n624), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n770), .A2(G116), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT46), .ZN(new_n945));
  INV_X1    g0745(.A(new_n786), .ZN(new_n946));
  AOI22_X1  g0746(.A1(G107), .A2(new_n946), .B1(new_n782), .B2(G294), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n792), .A2(G303), .B1(G311), .B2(new_n774), .ZN(new_n948));
  INV_X1    g0748(.A(G317), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n429), .B1(new_n762), .B2(new_n949), .C1(new_n768), .C2(new_n758), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G97), .B2(new_n766), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n945), .A2(new_n947), .A3(new_n948), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT108), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n774), .A2(new_n838), .B1(new_n782), .B2(G159), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n243), .B2(new_n786), .C1(new_n262), .C2(new_n779), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n766), .A2(G77), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n281), .B1(new_n758), .B2(new_n202), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G137), .B2(new_n763), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(new_n771), .C2(new_n403), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n953), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT47), .Z(new_n961));
  OAI221_X1 g0761(.A(new_n939), .B1(new_n940), .B2(new_n943), .C1(new_n961), .C2(new_n805), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n564), .A2(new_n661), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n570), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n569), .B2(new_n675), .ZN(new_n965));
  INV_X1    g0765(.A(new_n684), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT42), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n569), .B1(new_n964), .B2(new_n679), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n675), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(KEYINPUT42), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT105), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n673), .A2(new_n680), .A3(new_n965), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT104), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n975), .A2(new_n977), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n979), .A2(new_n980), .B1(KEYINPUT43), .B2(new_n943), .ZN(new_n981));
  INV_X1    g0781(.A(new_n980), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n983), .A3(new_n978), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n737), .B(KEYINPUT107), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n686), .A2(new_n965), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n686), .A2(new_n965), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(new_n681), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n684), .B1(new_n680), .B2(new_n683), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n673), .A2(KEYINPUT106), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n673), .A2(KEYINPUT106), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n994), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n733), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n689), .B(KEYINPUT41), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n986), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n962), .B1(new_n985), .B2(new_n1003), .ZN(G387));
  INV_X1    g0804(.A(new_n743), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n266), .A2(new_n202), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT50), .Z(new_n1007));
  AOI211_X1 g0807(.A(G45), .B(new_n690), .C1(G68), .C2(G77), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n473), .B2(new_n234), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n741), .A2(new_n690), .B1(new_n365), .B2(new_n688), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(KEYINPUT109), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n752), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT109), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n739), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n775), .A2(new_n794), .B1(new_n783), .B2(new_n377), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G50), .B2(new_n792), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n281), .B1(new_n762), .B2(new_n262), .C1(new_n243), .C2(new_n758), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G97), .B2(new_n766), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n617), .A2(new_n946), .A3(new_n619), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n770), .A2(G77), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n782), .A2(G311), .B1(new_n801), .B2(G303), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n779), .B2(new_n949), .C1(new_n780), .C2(new_n775), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n770), .A2(G294), .B1(G283), .B2(new_n946), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n429), .B1(new_n776), .B2(new_n762), .C1(new_n767), .C2(new_n580), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1022), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1015), .B1(new_n1035), .B2(new_n751), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n680), .B2(new_n940), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT110), .Z(new_n1038));
  INV_X1    g0838(.A(new_n999), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1038), .B1(new_n1039), .B2(new_n986), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n733), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n997), .A2(new_n998), .A3(new_n733), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n689), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1040), .B1(new_n1041), .B2(new_n1043), .ZN(G393));
  NAND2_X1  g0844(.A1(new_n992), .A2(new_n986), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n429), .B1(new_n763), .B2(new_n838), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n767), .B2(new_n417), .C1(new_n243), .C2(new_n771), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT111), .Z(new_n1048));
  OAI22_X1  g0848(.A1(new_n775), .A2(new_n262), .B1(new_n779), .B2(new_n794), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT51), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n782), .A2(G50), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n786), .A2(new_n280), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n266), .B2(new_n801), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n429), .B1(new_n762), .B2(new_n780), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1055), .B(new_n789), .C1(G283), .C2(new_n770), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n946), .A2(G116), .B1(new_n801), .B2(G294), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n769), .B2(new_n783), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT112), .Z(new_n1059));
  OAI22_X1  g0859(.A1(new_n775), .A2(new_n949), .B1(new_n779), .B2(new_n759), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1056), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n805), .B1(new_n1054), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1005), .A2(new_n241), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n753), .B(new_n1064), .C1(G97), .C2(new_n688), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1063), .A2(new_n738), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n965), .B2(new_n940), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n689), .B1(new_n993), .B2(new_n1042), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n992), .B1(new_n1039), .B2(new_n733), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1045), .B(new_n1067), .C1(new_n1068), .C2(new_n1069), .ZN(G390));
  OAI211_X1 g0870(.A(new_n458), .B(G330), .C1(new_n728), .C2(new_n923), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n860), .A3(new_n653), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT114), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n860), .A3(KEYINPUT114), .A4(new_n653), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n714), .A2(new_n675), .A3(new_n817), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n671), .B(new_n822), .C1(new_n728), .C2(new_n730), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n864), .B(new_n1076), .C1(new_n1077), .C2(new_n921), .ZN(new_n1078));
  OAI21_X1  g0878(.A(G330), .B1(new_n728), .B2(new_n923), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT115), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(KEYINPUT115), .B(G330), .C1(new_n728), .C2(new_n923), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n822), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1078), .B1(new_n1083), .B2(new_n921), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n924), .A2(G330), .A3(new_n822), .A4(new_n879), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1077), .A2(new_n921), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1085), .A2(new_n1086), .B1(new_n818), .B2(new_n864), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1074), .B(new_n1075), .C1(new_n1084), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1085), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n868), .A2(new_n870), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n675), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n903), .A2(new_n916), .B1(new_n880), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT38), .B1(new_n908), .B2(new_n911), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n893), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1076), .A2(new_n864), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n1095), .B2(new_n879), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1089), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n879), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1094), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n893), .A2(new_n896), .A3(new_n915), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT39), .B1(new_n902), .B2(new_n913), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n818), .A2(new_n864), .B1(new_n876), .B2(new_n878), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1101), .A2(new_n1102), .B1(new_n917), .B2(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1077), .A2(new_n921), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1100), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1097), .A2(new_n1106), .A3(KEYINPUT113), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT113), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1100), .A2(new_n1104), .A3(new_n1108), .A4(new_n1105), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1088), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(KEYINPUT116), .B1(new_n1110), .B2(new_n735), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT116), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1112), .B(new_n689), .C1(new_n1113), .C2(new_n1088), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT117), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT117), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1107), .A2(new_n1117), .A3(new_n1109), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1088), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1111), .A2(new_n1114), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(G125), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n281), .B1(new_n762), .B2(new_n1121), .C1(new_n758), .C2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G159), .A2(new_n946), .B1(new_n782), .B2(G137), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n775), .C1(new_n843), .C2(new_n779), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1123), .B(new_n1126), .C1(G50), .C2(new_n766), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n770), .A2(G150), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT53), .Z(new_n1129));
  OAI22_X1  g0929(.A1(new_n779), .A2(new_n580), .B1(new_n783), .B2(new_n365), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1052), .B(new_n1130), .C1(G283), .C2(new_n774), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n429), .B1(new_n762), .B2(new_n462), .C1(new_n531), .C2(new_n758), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1132), .B(new_n845), .C1(G87), .C2(new_n770), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1127), .A2(new_n1129), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n739), .B1(new_n266), .B2(new_n830), .C1(new_n1134), .C2(new_n805), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT118), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n903), .A2(new_n916), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n748), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1115), .B2(new_n986), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1120), .A2(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT121), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n925), .A2(new_n928), .A3(G330), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n273), .A2(new_n659), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n314), .B(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n919), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n925), .A2(new_n928), .A3(G330), .A4(new_n1147), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1142), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n919), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(KEYINPUT121), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT122), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1110), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1141), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1110), .A2(new_n1161), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1141), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n735), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1154), .A2(new_n1158), .A3(new_n986), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n739), .B1(G50), .B2(new_n830), .ZN(new_n1169));
  OR3_X1    g0969(.A1(new_n779), .A2(KEYINPUT119), .A3(new_n365), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n617), .A2(new_n619), .A3(new_n801), .ZN(new_n1171));
  OAI21_X1  g0971(.A(KEYINPUT119), .B1(new_n779), .B2(new_n365), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n766), .A2(G58), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1021), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n281), .A2(G41), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n768), .B2(new_n762), .C1(new_n243), .C2(new_n786), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n775), .A2(new_n580), .B1(new_n783), .B2(new_n531), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1173), .A2(new_n1175), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT58), .Z(new_n1180));
  OAI22_X1  g0980(.A1(new_n783), .A2(new_n843), .B1(new_n262), .B2(new_n786), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G125), .B2(new_n774), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n792), .A2(G128), .B1(G137), .B2(new_n801), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(new_n771), .C2(new_n1122), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n766), .A2(G159), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G33), .B(G41), .C1(new_n763), .C2(G124), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1180), .B1(new_n1185), .B2(new_n1189), .C1(new_n1176), .C2(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT120), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n805), .B1(new_n1191), .B2(KEYINPUT120), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1169), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1147), .B2(new_n749), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1168), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1167), .A2(new_n1196), .ZN(G375));
  NOR2_X1   g0997(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n921), .A2(new_n748), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n739), .B1(G68), .B2(new_n830), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n792), .A2(G137), .B1(G50), .B2(new_n946), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n843), .B2(new_n775), .C1(new_n783), .C2(new_n1122), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n281), .B1(new_n762), .B2(new_n1125), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G150), .B2(new_n801), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1174), .B(new_n1205), .C1(new_n771), .C2(new_n794), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n792), .A2(G283), .B1(G294), .B2(new_n774), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n580), .B2(new_n783), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n770), .A2(G97), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n429), .B1(new_n758), .B2(new_n365), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G303), .B2(new_n763), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n956), .A2(new_n1209), .A3(new_n1020), .A4(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1203), .A2(new_n1206), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1201), .B1(new_n1213), .B2(new_n751), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1199), .A2(new_n986), .B1(new_n1200), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1198), .A2(new_n1160), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n1002), .A3(new_n1088), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(G381));
  INV_X1    g1018(.A(KEYINPUT124), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G378), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1120), .A2(KEYINPUT124), .A3(new_n1139), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(new_n1167), .A3(new_n1196), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(G390), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n851), .ZN(new_n1226));
  OR4_X1    g1026(.A1(G396), .A2(new_n1226), .A3(G387), .A4(G393), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(G381), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1228), .A2(KEYINPUT123), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(KEYINPUT123), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1224), .B1(new_n1229), .B2(new_n1230), .ZN(G407));
  OAI211_X1 g1031(.A(G407), .B(G213), .C1(G343), .C2(new_n1223), .ZN(G409));
  OAI211_X1 g1032(.A(new_n962), .B(G390), .C1(new_n985), .C2(new_n1003), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT126), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(G393), .B(G396), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(new_n1225), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1233), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(KEYINPUT126), .A3(new_n1233), .A4(new_n1236), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1088), .A2(KEYINPUT60), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1245), .A2(new_n1216), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n689), .B1(new_n1245), .B2(new_n1216), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1215), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(new_n851), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n851), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n660), .A2(G213), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(G2897), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1251), .B(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1164), .A2(new_n1002), .A3(new_n1158), .A4(new_n1154), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n986), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1195), .A3(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1220), .A2(new_n1221), .A3(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1167), .A2(G378), .A3(new_n1196), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1253), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1253), .B(new_n1251), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1244), .B1(new_n1256), .B2(new_n1262), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1251), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1252), .A3(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1243), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(KEYINPUT125), .B1(new_n1263), .B2(KEYINPUT63), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT125), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1268), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1252), .A4(new_n1267), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1242), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1244), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT127), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1275), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1270), .B1(new_n1281), .B2(new_n1282), .ZN(G405));
  NAND2_X1  g1083(.A1(new_n1222), .A2(G375), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1284), .A2(new_n1261), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1285), .A2(new_n1251), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1251), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1286), .A2(new_n1243), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1243), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G402));
endmodule


