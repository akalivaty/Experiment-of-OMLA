//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040;
  XNOR2_X1  g000(.A(KEYINPUT11), .B(G169gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(G113gat), .B(G141gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(G1gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G1gat), .B2(new_n208), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G8gat), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n211), .B(new_n214), .C1(G1gat), .C2(new_n208), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT98), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT98), .B1(new_n213), .B2(new_n215), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  XOR2_X1   g020(.A(G43gat), .B(G50gat), .Z(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n221), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT96), .B(G29gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G36gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT97), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n226), .A2(G36gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT97), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n223), .A2(new_n225), .A3(new_n228), .A4(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n224), .B1(new_n229), .B2(new_n220), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n233), .B1(new_n232), .B2(new_n234), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n218), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n213), .A2(new_n215), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n234), .B2(new_n232), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT99), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n238), .A2(KEYINPUT99), .A3(new_n241), .A4(new_n242), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT100), .B(KEYINPUT18), .Z(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n238), .A2(KEYINPUT18), .A3(new_n241), .A4(new_n242), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n239), .A2(new_n234), .A3(new_n232), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n242), .B(KEYINPUT13), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT95), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n207), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI211_X1 g057(.A(KEYINPUT95), .B(new_n206), .C1(new_n248), .C2(new_n254), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G127gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT71), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G127gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n266), .A3(G134gat), .ZN(new_n267));
  INV_X1    g066(.A(G134gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G113gat), .B(G120gat), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n267), .B(new_n269), .C1(KEYINPUT1), .C2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G120gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G113gat), .ZN(new_n273));
  INV_X1    g072(.A(G113gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G120gat), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT1), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277));
  NAND2_X1  g076(.A1(G127gat), .A2(G134gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(G127gat), .A2(G134gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n269), .A2(KEYINPUT72), .A3(new_n278), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n271), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(G183gat), .B(G190gat), .C1(KEYINPUT68), .C2(KEYINPUT24), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n288), .B(new_n289), .C1(G183gat), .C2(G190gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n290), .A2(new_n293), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT25), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NOR3_X1   g098(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n285), .A2(KEYINPUT24), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n287), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n292), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n294), .B(KEYINPUT66), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT25), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI22_X1  g106(.A1(KEYINPUT67), .A2(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n297), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT27), .B(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT28), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n318));
  NOR4_X1   g117(.A1(new_n318), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT26), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT69), .B1(new_n291), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n319), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n285), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT70), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n291), .A2(new_n320), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n318), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n291), .A2(KEYINPUT69), .A3(new_n320), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n329), .A2(new_n323), .A3(new_n322), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n332), .A3(new_n285), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n317), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n284), .B1(new_n310), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n302), .A2(new_n303), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT65), .ZN(new_n338));
  INV_X1    g137(.A(G183gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n312), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n298), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n293), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n294), .B(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n336), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n345), .A2(new_n308), .B1(KEYINPUT25), .B2(new_n296), .ZN(new_n346));
  INV_X1    g145(.A(new_n284), .ZN(new_n347));
  INV_X1    g146(.A(new_n317), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n325), .A2(KEYINPUT70), .A3(new_n326), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n332), .B1(new_n331), .B2(new_n285), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT64), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT32), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT33), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G15gat), .B(G43gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n356), .B(KEYINPUT32), .C1(new_n358), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT34), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n335), .A2(new_n352), .A3(KEYINPUT73), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT73), .B1(new_n335), .B2(new_n352), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n367), .B1(new_n370), .B2(new_n353), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n335), .A2(new_n352), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(new_n367), .A3(new_n354), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT74), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT34), .B1(new_n335), .B2(new_n352), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n354), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n366), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  AND4_X1   g178(.A1(new_n376), .A2(new_n372), .A3(new_n367), .A4(new_n354), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n376), .B1(new_n375), .B2(new_n354), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT73), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n335), .A2(new_n352), .A3(KEYINPUT73), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n353), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT34), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n382), .A2(new_n387), .A3(new_n365), .A4(new_n363), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT75), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n379), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n366), .B(KEYINPUT75), .C1(new_n371), .C2(new_n378), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(KEYINPUT36), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT36), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n379), .A2(new_n388), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G8gat), .B(G36gat), .ZN(new_n396));
  INV_X1    g195(.A(G64gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n346), .B2(new_n351), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n310), .B2(new_n334), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n406));
  NOR2_X1   g205(.A1(KEYINPUT76), .A2(G204gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(KEYINPUT76), .A2(G204gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(G197gat), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G197gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n409), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n407), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT77), .B(G218gat), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT22), .B1(new_n415), .B2(G211gat), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT78), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G218gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT77), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT77), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G218gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n421), .A3(G211gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT22), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n410), .A4(new_n413), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G211gat), .B(G218gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n406), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n430), .B1(new_n417), .B2(new_n426), .ZN(new_n433));
  INV_X1    g232(.A(new_n431), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT79), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n405), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n401), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n310), .B2(new_n334), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n433), .A2(new_n434), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT29), .B1(new_n346), .B2(new_n351), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n439), .B(new_n441), .C1(new_n442), .C2(new_n438), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n400), .B1(new_n437), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n439), .B1(new_n442), .B2(new_n438), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n432), .B2(new_n435), .ZN(new_n447));
  INV_X1    g246(.A(new_n400), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n443), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n447), .A2(new_n451), .A3(new_n448), .A4(new_n443), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT0), .B(G57gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(G85gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G1gat), .B(G29gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g257(.A(G155gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT83), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT83), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G155gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n462), .A3(G162gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(KEYINPUT84), .A3(KEYINPUT2), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G155gat), .B(G162gat), .ZN(new_n466));
  INV_X1    g265(.A(G141gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  INV_X1    g267(.A(G148gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(G148gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n466), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT84), .B1(new_n463), .B2(KEYINPUT2), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n465), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G162gat), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT2), .B1(new_n459), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT81), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n469), .A2(G141gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(KEYINPUT81), .B(KEYINPUT2), .C1(new_n459), .C2(new_n478), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n466), .A2(KEYINPUT80), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n466), .A2(KEYINPUT80), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT3), .B1(new_n477), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n463), .A2(KEYINPUT2), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(G155gat), .B(G162gat), .Z(new_n493));
  INV_X1    g292(.A(new_n471), .ZN(new_n494));
  NOR2_X1   g293(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n495));
  OAI21_X1  g294(.A(G141gat), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n493), .B1(new_n473), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n492), .A2(new_n497), .A3(new_n464), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n485), .A2(new_n487), .A3(new_n486), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT3), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n489), .A2(new_n347), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT85), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n489), .A2(new_n504), .A3(new_n347), .A4(new_n501), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n498), .A2(new_n284), .A3(new_n499), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g307(.A1(G225gat), .A2(G233gat), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n477), .A2(new_n488), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(KEYINPUT4), .A3(new_n284), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n506), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n512), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n347), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n507), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n510), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(KEYINPUT5), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n520));
  OR2_X1    g319(.A1(KEYINPUT86), .A2(KEYINPUT4), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n507), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(KEYINPUT86), .A2(KEYINPUT4), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n523), .B(KEYINPUT87), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n524), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n503), .B2(new_n505), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n520), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n527), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n526), .B1(new_n507), .B2(new_n521), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND4_X1   g333(.A1(new_n520), .A2(new_n506), .A3(new_n534), .A4(new_n530), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n458), .B(new_n519), .C1(new_n531), .C2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n519), .B1(new_n531), .B2(new_n535), .ZN(new_n539));
  INV_X1    g338(.A(new_n458), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n500), .B1(new_n498), .B2(new_n499), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n504), .B1(new_n545), .B2(new_n347), .ZN(new_n546));
  INV_X1    g345(.A(new_n505), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n534), .B(new_n530), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT88), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n506), .A2(new_n520), .A3(new_n534), .A4(new_n530), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n551), .A2(KEYINPUT89), .A3(new_n458), .A4(new_n519), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n538), .A2(new_n541), .A3(new_n542), .A4(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n458), .B1(new_n551), .B2(new_n519), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT6), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n454), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(G228gat), .ZN(new_n557));
  INV_X1    g356(.A(G233gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n403), .B1(new_n433), .B2(new_n434), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n512), .B1(new_n561), .B2(new_n500), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n501), .A2(new_n403), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n440), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n432), .B2(new_n435), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n559), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n561), .A2(new_n500), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n515), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n429), .A2(new_n406), .A3(new_n431), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT79), .B1(new_n433), .B2(new_n434), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n571), .A2(new_n572), .B1(new_n403), .B2(new_n501), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n573), .B2(KEYINPUT90), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n565), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(G22gat), .ZN(new_n576));
  INV_X1    g375(.A(G22gat), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(new_n565), .C1(new_n568), .C2(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G78gat), .B(G106gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT31), .ZN(new_n581));
  INV_X1    g380(.A(G50gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n562), .B1(new_n566), .B2(new_n567), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n560), .B1(new_n573), .B2(KEYINPUT90), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n562), .A2(new_n564), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n585), .A2(new_n586), .B1(new_n587), .B2(new_n560), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT91), .B1(new_n588), .B2(new_n577), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n579), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n576), .B(new_n578), .C1(KEYINPUT91), .C2(new_n583), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n395), .B1(new_n556), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT40), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT93), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n509), .B1(new_n506), .B2(new_n534), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n540), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n516), .A2(new_n509), .A3(new_n507), .ZN(new_n601));
  OAI211_X1 g400(.A(KEYINPUT39), .B(new_n601), .C1(new_n529), .C2(new_n509), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n597), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n453), .A2(new_n554), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(new_n597), .A3(new_n602), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n604), .A2(new_n605), .B1(new_n591), .B2(new_n590), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n607), .B(new_n443), .C1(new_n405), .C2(new_n436), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n400), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n447), .B2(new_n443), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT38), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT94), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n613), .B(KEYINPUT38), .C1(new_n609), .C2(new_n610), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n614), .A2(new_n449), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n553), .A2(new_n555), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n609), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n446), .A2(new_n441), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n619), .B(KEYINPUT37), .C1(new_n446), .C2(new_n436), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n606), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n395), .B(KEYINPUT92), .C1(new_n556), .C2(new_n592), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n595), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n553), .A2(new_n555), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n590), .A2(new_n591), .B1(new_n390), .B2(new_n391), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n453), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT35), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT35), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n379), .A2(new_n388), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n590), .B2(new_n591), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n556), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n262), .B1(new_n625), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636));
  INV_X1    g435(.A(G211gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n397), .A2(G57gat), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT101), .B(G57gat), .Z(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n640), .B2(new_n397), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G71gat), .A2(G78gat), .ZN(new_n644));
  OR2_X1    g443(.A1(G71gat), .A2(G78gat), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT9), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(KEYINPUT102), .B(new_n639), .C1(new_n640), .C2(new_n397), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n643), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G57gat), .B(G64gat), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n644), .B(new_n645), .C1(new_n650), .C2(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT21), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n239), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G183gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(G231gat), .A2(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n638), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  INV_X1    g460(.A(new_n638), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n652), .A2(new_n653), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n660), .A2(new_n663), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n237), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n235), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  INV_X1    g473(.A(G85gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n675), .B2(new_n399), .ZN(new_n676));
  NAND3_X1  g475(.A1(KEYINPUT103), .A2(G85gat), .A3(G92gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(KEYINPUT7), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G99gat), .A2(G106gat), .ZN(new_n679));
  AOI22_X1  g478(.A1(KEYINPUT8), .A2(new_n679), .B1(new_n675), .B2(new_n399), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT7), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n674), .B(new_n681), .C1(new_n675), .C2(new_n399), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n678), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(G99gat), .B(G106gat), .Z(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n684), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n686), .A2(new_n680), .A3(new_n678), .A4(new_n682), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(KEYINPUT104), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n683), .A2(new_n689), .A3(new_n684), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n673), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n232), .A2(new_n234), .ZN(new_n696));
  AND2_X1   g495(.A1(G232gat), .A2(G233gat), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n691), .A2(new_n696), .B1(KEYINPUT41), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n673), .A2(KEYINPUT105), .A3(new_n692), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(G134gat), .B(G162gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n697), .A2(KEYINPUT41), .ZN(new_n703));
  XNOR2_X1  g502(.A(G190gat), .B(G218gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n700), .A2(new_n701), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n700), .A2(new_n701), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(G230gat), .A2(G233gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n691), .A2(new_n652), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n685), .A2(new_n687), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n649), .A2(new_n714), .A3(new_n651), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT10), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n691), .A2(KEYINPUT10), .A3(new_n651), .A4(new_n649), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n712), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n712), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n713), .A2(new_n720), .A3(new_n715), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(G176gat), .B(G204gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT106), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G120gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(new_n469), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n722), .B(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n671), .A2(new_n711), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n635), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n626), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT107), .B(G1gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1324gat));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n453), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n209), .A2(new_n214), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n209), .A2(new_n214), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n734), .A2(KEYINPUT42), .A3(new_n736), .A4(new_n737), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n740), .B(new_n741), .C1(new_n214), .C2(new_n734), .ZN(G1325gat));
  INV_X1    g541(.A(new_n730), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n392), .A2(KEYINPUT108), .A3(new_n394), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT108), .B1(new_n392), .B2(new_n394), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n743), .A2(G15gat), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n631), .ZN(new_n749));
  AOI21_X1  g548(.A(G15gat), .B1(new_n743), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n748), .A2(new_n750), .ZN(G1326gat));
  NOR2_X1   g550(.A1(new_n730), .A2(new_n592), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT43), .B(G22gat), .Z(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1327gat));
  INV_X1    g553(.A(new_n711), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n625), .B2(new_n634), .ZN(new_n756));
  INV_X1    g555(.A(new_n671), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n757), .A2(new_n262), .A3(new_n728), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n626), .A2(new_n226), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT45), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n392), .A2(new_n394), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n392), .A2(KEYINPUT108), .A3(new_n394), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n765), .B(new_n766), .C1(new_n556), .C2(new_n592), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n453), .A2(new_n603), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n541), .A3(new_n605), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n592), .ZN(new_n770));
  AND4_X1   g569(.A1(new_n553), .A2(new_n555), .A3(new_n612), .A4(new_n615), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n621), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n630), .B1(new_n556), .B2(new_n627), .ZN(new_n773));
  AND4_X1   g572(.A1(new_n630), .A2(new_n626), .A3(new_n453), .A4(new_n632), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n767), .A2(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT44), .B1(new_n775), .B2(new_n711), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(KEYINPUT44), .B2(new_n756), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n758), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n226), .B1(new_n778), .B2(new_n626), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n779), .ZN(G1328gat));
  INV_X1    g579(.A(G36gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n759), .A2(new_n781), .A3(new_n454), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(KEYINPUT46), .ZN(new_n783));
  OAI21_X1  g582(.A(G36gat), .B1(new_n778), .B2(new_n453), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(KEYINPUT46), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(G1329gat));
  NAND2_X1  g585(.A1(new_n759), .A2(new_n749), .ZN(new_n787));
  INV_X1    g586(.A(G43gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n777), .A2(G43gat), .A3(new_n747), .A4(new_n758), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT47), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1330gat));
  INV_X1    g594(.A(new_n592), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n777), .A2(KEYINPUT109), .A3(new_n796), .A4(new_n758), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n625), .A2(new_n634), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(KEYINPUT44), .A3(new_n711), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n775), .A2(new_n711), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n799), .A2(new_n802), .A3(new_n796), .A4(new_n758), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n797), .A2(new_n805), .A3(G50gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n759), .A2(new_n582), .A3(new_n796), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT48), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n803), .A2(G50gat), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n807), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n806), .A2(new_n808), .B1(new_n810), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g610(.A1(new_n757), .A2(new_n755), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n261), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n775), .A2(new_n728), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n553), .A2(new_n555), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(new_n640), .ZN(G1332gat));
  INV_X1    g616(.A(new_n814), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n453), .ZN(new_n819));
  NOR2_X1   g618(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n820));
  AND2_X1   g619(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n822), .B1(new_n819), .B2(new_n820), .ZN(G1333gat));
  NAND3_X1  g622(.A1(new_n814), .A2(G71gat), .A3(new_n747), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n814), .A2(KEYINPUT110), .A3(G71gat), .A4(new_n747), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(G71gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n818), .B2(new_n631), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT50), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n833), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(G1334gat));
  NAND2_X1  g634(.A1(new_n814), .A2(new_n796), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g636(.A1(new_n757), .A2(new_n261), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n728), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n777), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(new_n675), .A3(new_n626), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n843));
  AND4_X1   g642(.A1(new_n843), .A2(new_n775), .A3(new_n711), .A4(new_n838), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n796), .B1(new_n815), .B2(new_n454), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n746), .A3(new_n623), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n755), .B1(new_n846), .B2(new_n634), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n843), .B1(new_n847), .B2(new_n838), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n815), .A3(new_n728), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n842), .B1(new_n675), .B2(new_n850), .ZN(G1336gat));
  NAND3_X1  g650(.A1(new_n775), .A2(new_n711), .A3(new_n838), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT51), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n847), .A2(new_n843), .A3(new_n838), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n454), .A3(new_n728), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n399), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n453), .A2(new_n399), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n841), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n856), .B(KEYINPUT52), .C1(new_n841), .C2(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1337gat));
  OAI21_X1  g662(.A(G99gat), .B1(new_n841), .B2(new_n746), .ZN(new_n864));
  INV_X1    g663(.A(G99gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n865), .A3(new_n728), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n631), .B2(new_n866), .ZN(G1338gat));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n592), .A2(G106gat), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n849), .A2(new_n868), .A3(new_n728), .A4(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n799), .A2(new_n802), .A3(new_n796), .A4(new_n840), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT111), .B(G106gat), .Z(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n728), .A3(new_n854), .A4(new_n869), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT112), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT53), .ZN(new_n877));
  XNOR2_X1  g676(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(G1339gat));
  NAND3_X1  g679(.A1(new_n248), .A2(new_n206), .A3(new_n254), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n251), .A2(new_n252), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n242), .B1(new_n238), .B2(new_n241), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n205), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n726), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n722), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT10), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n690), .A2(new_n688), .B1(new_n649), .B2(new_n651), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n649), .A2(new_n714), .A3(new_n651), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n720), .B1(new_n891), .B2(new_n717), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n726), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n720), .A3(new_n717), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n719), .A2(KEYINPUT54), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n887), .B1(new_n898), .B2(KEYINPUT55), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT55), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AND4_X1   g700(.A1(new_n711), .A2(new_n885), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n899), .B(new_n901), .C1(new_n257), .C2(new_n259), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n728), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n711), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n671), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n729), .A2(new_n262), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n908), .A2(new_n815), .A3(new_n453), .A4(new_n632), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT114), .ZN(new_n910));
  OAI21_X1  g709(.A(G113gat), .B1(new_n910), .B2(new_n262), .ZN(new_n911));
  INV_X1    g710(.A(new_n908), .ZN(new_n912));
  INV_X1    g711(.A(new_n627), .ZN(new_n913));
  NOR4_X1   g712(.A1(new_n912), .A2(new_n626), .A3(new_n454), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n274), .A3(new_n261), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n915), .ZN(G1340gat));
  OAI21_X1  g715(.A(G120gat), .B1(new_n910), .B2(new_n727), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n272), .A3(new_n728), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1341gat));
  AND2_X1   g718(.A1(new_n264), .A2(new_n266), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n914), .B2(new_n757), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n910), .A2(new_n671), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n920), .ZN(G1342gat));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n268), .A3(new_n711), .ZN(new_n924));
  XOR2_X1   g723(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G134gat), .B1(new_n910), .B2(new_n755), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1343gat));
  NAND2_X1  g727(.A1(new_n897), .A2(KEYINPUT116), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n894), .A2(new_n896), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n929), .A2(new_n900), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n899), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(new_n899), .A3(KEYINPUT117), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n261), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n711), .B1(new_n937), .B2(new_n904), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n671), .B1(new_n938), .B2(new_n902), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n592), .B1(new_n939), .B2(new_n907), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT57), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n746), .A2(new_n815), .A3(new_n453), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n592), .B1(new_n906), .B2(new_n907), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n941), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n467), .B1(new_n947), .B2(new_n261), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n908), .A2(new_n796), .ZN(new_n949));
  NOR4_X1   g748(.A1(new_n949), .A2(G141gat), .A3(new_n262), .A4(new_n943), .ZN(new_n950));
  XNOR2_X1  g749(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OR3_X1    g751(.A1(new_n948), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n948), .B2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1344gat));
  NOR2_X1   g754(.A1(new_n912), .A2(new_n626), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n494), .A2(new_n495), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n747), .A2(new_n957), .A3(new_n592), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n956), .A2(new_n453), .A3(new_n728), .A4(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n945), .B(new_n728), .C1(new_n940), .C2(new_n941), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT59), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n960), .A2(new_n961), .A3(new_n957), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n261), .A2(new_n936), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT117), .B1(new_n932), .B2(new_n899), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n904), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n755), .ZN(new_n966));
  INV_X1    g765(.A(new_n902), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n757), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n907), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n941), .B(new_n796), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n949), .A2(KEYINPUT57), .ZN(new_n971));
  INV_X1    g770(.A(new_n943), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n970), .A2(new_n971), .A3(new_n728), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n961), .B1(new_n973), .B2(G148gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n959), .B1(new_n962), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT119), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT119), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n977), .B(new_n959), .C1(new_n962), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1345gat));
  NOR2_X1   g778(.A1(new_n949), .A2(new_n943), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n757), .ZN(new_n981));
  XOR2_X1   g780(.A(new_n981), .B(KEYINPUT120), .Z(new_n982));
  NAND2_X1  g781(.A1(new_n460), .A2(new_n462), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n671), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g783(.A(new_n984), .B(KEYINPUT121), .Z(new_n985));
  AOI22_X1  g784(.A1(new_n982), .A2(new_n983), .B1(new_n947), .B2(new_n985), .ZN(G1346gat));
  AOI21_X1  g785(.A(G162gat), .B1(new_n980), .B2(new_n711), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n942), .A2(new_n946), .A3(new_n755), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n987), .B1(new_n988), .B2(G162gat), .ZN(G1347gat));
  NAND3_X1  g788(.A1(new_n908), .A2(new_n626), .A3(new_n454), .ZN(new_n990));
  NOR4_X1   g789(.A1(new_n990), .A2(G169gat), .A3(new_n262), .A4(new_n913), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT122), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n908), .A2(new_n626), .A3(new_n454), .A4(new_n632), .ZN(new_n993));
  OAI21_X1  g792(.A(G169gat), .B1(new_n993), .B2(new_n262), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(G1348gat));
  NOR2_X1   g794(.A1(new_n990), .A2(new_n913), .ZN(new_n996));
  AOI21_X1  g795(.A(G176gat), .B1(new_n996), .B2(new_n728), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n993), .A2(new_n727), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n997), .B1(new_n998), .B2(G176gat), .ZN(G1349gat));
  NAND3_X1  g798(.A1(new_n996), .A2(new_n311), .A3(new_n757), .ZN(new_n1000));
  OAI21_X1  g799(.A(G183gat), .B1(new_n993), .B2(new_n671), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1002), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g802(.A(G190gat), .B1(new_n993), .B2(new_n755), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT61), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n996), .A2(new_n312), .A3(new_n711), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(G1351gat));
  NAND3_X1  g806(.A1(new_n746), .A2(new_n626), .A3(new_n454), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n949), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1009), .A2(KEYINPUT123), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT123), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1011), .B1(new_n949), .B2(new_n1008), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1010), .A2(new_n261), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(new_n411), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n970), .A2(new_n971), .ZN(new_n1015));
  INV_X1    g814(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g815(.A(KEYINPUT124), .ZN(new_n1017));
  XNOR2_X1  g816(.A(new_n1008), .B(new_n1017), .ZN(new_n1018));
  NOR3_X1   g817(.A1(new_n1018), .A2(new_n411), .A3(new_n262), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g820(.A(new_n1021), .B(KEYINPUT125), .ZN(G1352gat));
  NAND2_X1  g821(.A1(new_n1016), .A2(new_n728), .ZN(new_n1023));
  OAI21_X1  g822(.A(G204gat), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1024));
  NOR4_X1   g823(.A1(new_n949), .A2(G204gat), .A3(new_n727), .A4(new_n1008), .ZN(new_n1025));
  XNOR2_X1  g824(.A(new_n1025), .B(KEYINPUT62), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1024), .A2(new_n1026), .ZN(G1353gat));
  OR3_X1    g826(.A1(new_n1015), .A2(new_n671), .A3(new_n1008), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1028), .A2(G211gat), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1029), .A2(KEYINPUT63), .ZN(new_n1030));
  NAND4_X1  g829(.A1(new_n1010), .A2(new_n637), .A3(new_n757), .A4(new_n1012), .ZN(new_n1031));
  XNOR2_X1  g830(.A(new_n1031), .B(KEYINPUT126), .ZN(new_n1032));
  INV_X1    g831(.A(KEYINPUT63), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1028), .A2(new_n1033), .A3(G211gat), .ZN(new_n1034));
  NAND3_X1  g833(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(G1354gat));
  NAND3_X1  g834(.A1(new_n1010), .A2(new_n711), .A3(new_n1012), .ZN(new_n1036));
  AND3_X1   g835(.A1(new_n1036), .A2(KEYINPUT127), .A3(new_n418), .ZN(new_n1037));
  AOI21_X1  g836(.A(KEYINPUT127), .B1(new_n1036), .B2(new_n418), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n711), .A2(new_n415), .ZN(new_n1039));
  NOR3_X1   g838(.A1(new_n1015), .A2(new_n1018), .A3(new_n1039), .ZN(new_n1040));
  NOR3_X1   g839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(G1355gat));
endmodule


