//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT11), .B(G169gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G1gat), .ZN(new_n210));
  INV_X1    g009(.A(G22gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G15gat), .ZN(new_n212));
  INV_X1    g011(.A(G15gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G22gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT86), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(new_n210), .A3(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n207), .B(KEYINPUT86), .C1(new_n208), .C2(G1gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT87), .B(G8gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n216), .A2(new_n217), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT87), .A2(G8gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G43gat), .A2(G50gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G43gat), .A2(G50gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT83), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G43gat), .ZN(new_n226));
  INV_X1    g025(.A(G50gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229));
  NAND2_X1  g028(.A1(G43gat), .A2(G50gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n225), .A2(new_n231), .A3(KEYINPUT15), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n233), .A3(new_n230), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT14), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(G29gat), .B2(G36gat), .ZN(new_n236));
  INV_X1    g035(.A(G29gat), .ZN(new_n237));
  INV_X1    g036(.A(G36gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT14), .ZN(new_n239));
  NAND2_X1  g038(.A1(G29gat), .A2(G36gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n234), .A2(new_n236), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT84), .B1(new_n232), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n236), .A3(new_n240), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(KEYINPUT15), .A3(new_n225), .A4(new_n231), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n231), .A3(KEYINPUT15), .ZN(new_n245));
  INV_X1    g044(.A(new_n243), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .A4(new_n234), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n242), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n222), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G229gat), .A2(G233gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n242), .A2(KEYINPUT17), .A3(new_n244), .A4(new_n248), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT88), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n258));
  NAND2_X1  g057(.A1(new_n248), .A2(new_n244), .ZN(new_n259));
  AND4_X1   g058(.A1(new_n236), .A2(new_n234), .A3(new_n239), .A4(new_n240), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n247), .B1(new_n260), .B2(new_n245), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n221), .B1(new_n216), .B2(new_n217), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n250), .B(new_n254), .C1(new_n257), .C2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n248), .A2(new_n244), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n242), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(KEYINPUT89), .A3(new_n250), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n251), .B(KEYINPUT13), .Z(new_n271));
  OR3_X1    g070(.A1(new_n222), .A2(new_n249), .A3(KEYINPUT89), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n250), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n268), .A2(new_n256), .A3(KEYINPUT17), .A4(new_n242), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n255), .A2(KEYINPUT88), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n222), .B1(new_n249), .B2(new_n258), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT18), .B1(new_n280), .B2(new_n251), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n206), .B1(new_n274), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n251), .B(new_n250), .C1(new_n257), .C2(new_n266), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n253), .ZN(new_n284));
  INV_X1    g083(.A(new_n206), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n284), .A2(new_n273), .A3(new_n267), .A4(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G141gat), .B(G148gat), .Z(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT75), .ZN(new_n289));
  XNOR2_X1  g088(.A(G141gat), .B(G148gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT75), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT2), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G155gat), .B(G162gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n294), .A2(KEYINPUT76), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(KEYINPUT76), .ZN(new_n298));
  INV_X1    g097(.A(G155gat), .ZN(new_n299));
  INV_X1    g098(.A(G162gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT2), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n297), .A2(new_n288), .A3(new_n298), .A4(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT22), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT72), .B(G211gat), .ZN(new_n306));
  INV_X1    g105(.A(G218gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(G211gat), .B(G218gat), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n310), .B2(new_n311), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n304), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n303), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n310), .A2(new_n311), .ZN(new_n318));
  INV_X1    g117(.A(new_n312), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n296), .A2(new_n316), .A3(new_n302), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(KEYINPUT29), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G228gat), .ZN(new_n327));
  INV_X1    g126(.A(G233gat), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n317), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n296), .A2(new_n302), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT29), .B1(new_n320), .B2(new_n321), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(KEYINPUT3), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n327), .A2(new_n328), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n313), .A2(new_n314), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(KEYINPUT29), .B2(new_n324), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n211), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n329), .A2(new_n336), .A3(new_n211), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(G50gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT80), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n343), .B(KEYINPUT31), .Z(new_n344));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n337), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n338), .A2(new_n345), .A3(new_n339), .A4(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G169gat), .ZN(new_n350));
  INV_X1    g149(.A(G176gat), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT26), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(new_n350), .B2(new_n351), .ZN(new_n353));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT26), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT66), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT27), .B(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT65), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT28), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT28), .B1(new_n360), .B2(new_n363), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n358), .B(new_n359), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT64), .B1(new_n350), .B2(new_n351), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT23), .ZN(new_n369));
  OR2_X1    g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(KEYINPUT24), .A3(new_n354), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n354), .A2(KEYINPUT24), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(G169gat), .B2(G176gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n369), .A2(KEYINPUT25), .A3(new_n371), .A4(new_n373), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(G127gat), .A2(G134gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(G127gat), .A2(G134gat), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT1), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G113gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G120gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT69), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT68), .B(G120gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(new_n382), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n381), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT67), .B(G134gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G127gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G113gat), .B(G120gat), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n389), .B(new_n379), .C1(KEYINPUT1), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n367), .A2(new_n378), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT70), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n367), .A2(new_n378), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n392), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT70), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n367), .A2(new_n378), .A3(new_n399), .A4(new_n393), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n395), .A2(new_n397), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT34), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT32), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n400), .A3(new_n397), .ZN(new_n404));
  INV_X1    g203(.A(new_n398), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT33), .B1(new_n404), .B2(new_n405), .ZN(new_n407));
  XOR2_X1   g206(.A(G15gat), .B(G43gat), .Z(new_n408));
  XNOR2_X1  g207(.A(G71gat), .B(G99gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n406), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  AOI221_X4 g211(.A(new_n403), .B1(KEYINPUT33), .B2(new_n410), .C1(new_n404), .C2(new_n405), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n402), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT71), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(KEYINPUT71), .B(new_n402), .C1(new_n412), .C2(new_n413), .ZN(new_n417));
  INV_X1    g216(.A(new_n402), .ZN(new_n418));
  INV_X1    g217(.A(new_n406), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n405), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n422), .A3(new_n410), .ZN(new_n423));
  INV_X1    g222(.A(new_n413), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n418), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n349), .A2(new_n416), .A3(new_n417), .A4(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT0), .ZN(new_n428));
  XNOR2_X1  g227(.A(G57gat), .B(G85gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n330), .A2(new_n392), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n296), .A2(new_n302), .A3(new_n387), .A4(new_n391), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n330), .A2(KEYINPUT77), .A3(new_n392), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n431), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(new_n323), .A3(new_n392), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n434), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n303), .A2(new_n393), .A3(KEYINPUT4), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .A4(new_n438), .ZN(new_n445));
  INV_X1    g244(.A(new_n438), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n435), .A2(KEYINPUT78), .A3(new_n446), .A4(new_n436), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n439), .A2(KEYINPUT5), .A3(new_n445), .A4(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT79), .B1(new_n445), .B2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT5), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n452), .B2(new_n439), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n430), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n450), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n449), .A3(new_n439), .ZN(new_n457));
  INV_X1    g256(.A(new_n430), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n456), .A2(KEYINPUT6), .A3(new_n457), .A4(new_n458), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n396), .A2(KEYINPUT74), .ZN(new_n463));
  INV_X1    g262(.A(G226gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n328), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n367), .A2(new_n378), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n465), .A2(KEYINPUT29), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n396), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n334), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n367), .A2(new_n378), .A3(new_n465), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n463), .A2(new_n467), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(new_n469), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n471), .B1(new_n475), .B2(new_n334), .ZN(new_n476));
  XNOR2_X1  g275(.A(G8gat), .B(G36gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n477), .B(new_n478), .Z(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OR3_X1    g279(.A1(new_n476), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n367), .A2(new_n466), .A3(new_n378), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n466), .B1(new_n367), .B2(new_n378), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n469), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n334), .B1(new_n484), .B2(new_n472), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n471), .A3(new_n479), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n468), .A2(new_n334), .A3(new_n470), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n480), .B1(new_n488), .B2(new_n485), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(KEYINPUT30), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n462), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT35), .B1(new_n426), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n414), .A2(new_n425), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n348), .B2(new_n347), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n460), .A2(new_n461), .B1(new_n481), .B2(new_n490), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n414), .A2(new_n425), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n416), .A2(new_n417), .A3(new_n425), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n502), .B2(KEYINPUT36), .ZN(new_n503));
  INV_X1    g302(.A(new_n349), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n492), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n476), .A2(new_n480), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n468), .A2(new_n322), .A3(new_n470), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n507), .A2(KEYINPUT37), .ZN(new_n508));
  INV_X1    g307(.A(new_n484), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n334), .B1(new_n509), .B2(new_n473), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT38), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n480), .A2(KEYINPUT37), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n489), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n506), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n480), .B1(new_n476), .B2(KEYINPUT37), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n486), .B2(new_n471), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT38), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n514), .A2(new_n460), .A3(new_n461), .A4(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT40), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n444), .A2(new_n443), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n438), .B1(new_n521), .B2(new_n441), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT39), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n458), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n441), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n444), .A2(new_n443), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n446), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n437), .A2(new_n438), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT39), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n520), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI211_X1 g331(.A(KEYINPUT82), .B(KEYINPUT40), .C1(new_n524), .C2(new_n529), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(new_n481), .A3(new_n490), .A4(new_n459), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n535), .A3(new_n349), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n503), .A2(new_n505), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n287), .B1(new_n499), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(KEYINPUT41), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT93), .ZN(new_n541));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G190gat), .B(G218gat), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  INV_X1    g351(.A(G92gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n548), .A2(new_n551), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G99gat), .B(G106gat), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559));
  AOI22_X1  g358(.A1(KEYINPUT8), .A2(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n560));
  XNOR2_X1  g359(.A(G99gat), .B(G106gat), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n560), .A2(new_n561), .A3(new_n551), .A4(new_n555), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  OR3_X1    g362(.A1(new_n556), .A2(new_n559), .A3(new_n557), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n249), .B2(new_n258), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n278), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n259), .B2(new_n261), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n539), .A2(KEYINPUT41), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n546), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n545), .B(new_n570), .C1(new_n278), .C2(new_n566), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n544), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n565), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n262), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n576), .B1(new_n277), .B2(new_n276), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n545), .B1(new_n577), .B2(new_n570), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n567), .A2(new_n546), .A3(new_n571), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n543), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(new_n299), .ZN(new_n583));
  XNOR2_X1  g382(.A(G183gat), .B(G211gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G57gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(G64gat), .ZN(new_n588));
  INV_X1    g387(.A(G64gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(G57gat), .ZN(new_n590));
  OAI22_X1  g389(.A1(new_n588), .A2(new_n590), .B1(KEYINPUT90), .B2(KEYINPUT9), .ZN(new_n591));
  INV_X1    g390(.A(G71gat), .ZN(new_n592));
  INV_X1    g391(.A(G78gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OR3_X1    g393(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT90), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT90), .B1(new_n592), .B2(new_n593), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n591), .A2(new_n594), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT9), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n592), .B2(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n587), .A2(KEYINPUT91), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G57gat), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n600), .A2(new_n602), .A3(G64gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(new_n587), .B2(G64gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n589), .A2(KEYINPUT92), .A3(G57gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n599), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n597), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G127gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n609), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n222), .B1(KEYINPUT21), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n615), .A2(new_n617), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n586), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n615), .A2(new_n617), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(new_n618), .A3(new_n585), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n581), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT95), .Z(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n563), .A2(new_n564), .B1(new_n608), .B2(new_n597), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n558), .A2(new_n562), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n630), .A2(new_n608), .A3(new_n597), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n628), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n565), .A2(new_n616), .A3(KEYINPUT10), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n627), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n627), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n629), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n635), .A2(new_n637), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n625), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n538), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n462), .B(KEYINPUT96), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(new_n210), .ZN(G1324gat));
  NOR2_X1   g449(.A1(new_n647), .A2(new_n491), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(G8gat), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n651), .ZN(new_n655));
  MUX2_X1   g454(.A(new_n653), .B(new_n655), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g455(.A(G15gat), .B1(new_n647), .B2(new_n503), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n414), .A2(new_n425), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n213), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n657), .B1(new_n647), .B2(new_n660), .ZN(G1326gat));
  NAND3_X1  g460(.A1(new_n538), .A2(new_n504), .A3(new_n646), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT97), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  INV_X1    g464(.A(new_n648), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n621), .A2(new_n623), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n645), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n581), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT98), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n538), .A2(new_n237), .A3(new_n666), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n503), .A2(new_n505), .A3(new_n536), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n417), .A2(new_n425), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n423), .A2(new_n424), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT71), .B1(new_n676), .B2(new_n402), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n497), .A3(new_n349), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n679), .A2(KEYINPUT35), .B1(new_n497), .B2(new_n496), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n581), .B1(new_n674), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n499), .A2(new_n537), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(KEYINPUT44), .A3(new_n581), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n645), .B(KEYINPUT99), .Z(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(new_n287), .A3(new_n667), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n683), .A2(new_n685), .A3(new_n666), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G29gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1328gat));
  NAND2_X1  g491(.A1(new_n538), .A2(new_n671), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n693), .A2(G36gat), .A3(new_n491), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT46), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n683), .A2(new_n685), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n687), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(new_n491), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G36gat), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n698), .A2(new_n696), .A3(new_n491), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n695), .B1(new_n700), .B2(new_n701), .ZN(G1329gat));
  NOR3_X1   g501(.A1(new_n693), .A2(G43gat), .A3(new_n658), .ZN(new_n703));
  INV_X1    g502(.A(new_n503), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n683), .A2(new_n685), .A3(new_n704), .A4(new_n687), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(G43gat), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1330gat));
  NAND3_X1  g507(.A1(new_n697), .A2(new_n504), .A3(new_n687), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G50gat), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n538), .A2(new_n227), .A3(new_n504), .A4(new_n671), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT48), .B1(new_n711), .B2(KEYINPUT104), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(KEYINPUT104), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n711), .B(KEYINPUT103), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n715), .B1(new_n709), .B2(G50gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n716), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g516(.A(new_n686), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n282), .A2(new_n286), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n718), .A2(new_n625), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n684), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n648), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT105), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n600), .A2(new_n602), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1332gat));
  XNOR2_X1  g524(.A(new_n721), .B(KEYINPUT106), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n491), .B(KEYINPUT107), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n727), .B1(new_n726), .B2(new_n729), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n730), .A2(new_n731), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n726), .A2(new_n729), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT108), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(new_n737), .ZN(G1333gat));
  NAND3_X1  g537(.A1(new_n726), .A2(G71gat), .A3(new_n704), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n592), .B1(new_n721), .B2(new_n658), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n739), .A2(KEYINPUT50), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT50), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n504), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g544(.A1(new_n667), .A2(new_n719), .A3(new_n669), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n683), .A2(new_n685), .A3(new_n666), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G85gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n668), .A2(new_n287), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n681), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n581), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n499), .B2(new_n537), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n667), .A2(new_n719), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(KEYINPUT51), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n751), .A2(KEYINPUT109), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT51), .B1(new_n753), .B2(new_n754), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n648), .A2(G85gat), .A3(new_n669), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n748), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(KEYINPUT110), .B(new_n748), .C1(new_n760), .C2(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1336gat));
  INV_X1    g566(.A(new_n728), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n683), .A2(new_n685), .A3(new_n768), .A4(new_n746), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT52), .B1(new_n769), .B2(G92gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n553), .A3(new_n686), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n760), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n491), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n683), .A2(new_n685), .A3(new_n773), .A4(new_n746), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n771), .B(KEYINPUT111), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n681), .A2(new_n749), .A3(new_n750), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n757), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT112), .B1(new_n779), .B2(KEYINPUT52), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  AOI211_X1 g581(.A(new_n781), .B(new_n782), .C1(new_n775), .C2(new_n778), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n772), .B1(new_n780), .B2(new_n783), .ZN(G1337gat));
  NAND3_X1  g583(.A1(new_n697), .A2(new_n704), .A3(new_n746), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G99gat), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n658), .A2(G99gat), .A3(new_n669), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n760), .B2(new_n787), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n697), .A2(new_n504), .A3(new_n746), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n349), .A2(new_n718), .A3(G106gat), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT113), .Z(new_n794));
  AND3_X1   g593(.A1(new_n756), .A2(new_n759), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n751), .A2(new_n755), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n789), .A2(G106gat), .B1(new_n796), .B2(new_n794), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n792), .A2(new_n795), .B1(new_n797), .B2(new_n798), .ZN(G1339gat));
  AND3_X1   g598(.A1(new_n624), .A2(new_n287), .A3(new_n669), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n274), .A2(new_n281), .A3(new_n206), .ZN(new_n802));
  INV_X1    g601(.A(new_n205), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n266), .B1(new_n277), .B2(new_n276), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n252), .B1(new_n804), .B2(new_n275), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n270), .A2(new_n272), .ZN(new_n806));
  INV_X1    g605(.A(new_n271), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n803), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n801), .B1(new_n802), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI211_X1 g611(.A(new_n811), .B(new_n641), .C1(new_n634), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n632), .A2(new_n633), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(new_n636), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n632), .A2(KEYINPUT115), .A3(new_n627), .A4(new_n633), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n632), .A2(new_n627), .A3(new_n633), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n813), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n644), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n641), .B1(new_n634), .B2(new_n812), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT55), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n805), .A2(new_n808), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n205), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n286), .A2(new_n827), .A3(KEYINPUT116), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n810), .A2(new_n825), .A3(new_n581), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n274), .A2(new_n281), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n809), .B1(new_n830), .B2(new_n285), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n825), .A2(new_n719), .B1(new_n831), .B2(new_n645), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n829), .B1(new_n832), .B2(new_n581), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n800), .B1(new_n833), .B2(new_n668), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n504), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n835), .A2(new_n659), .A3(new_n666), .A4(new_n728), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n836), .A2(new_n382), .A3(new_n287), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n648), .A2(new_n426), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n825), .A2(new_n719), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n286), .A2(new_n827), .A3(new_n645), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n581), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n828), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n635), .A2(new_n637), .A3(new_n641), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n843), .B1(new_n813), .B2(new_n820), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n820), .A2(new_n823), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n811), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n581), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT116), .B1(new_n286), .B2(new_n827), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n842), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n668), .B1(new_n841), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n800), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n838), .A2(new_n728), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n853), .A2(new_n287), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n837), .B1(new_n382), .B2(new_n854), .ZN(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n836), .B2(new_n718), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n669), .A2(new_n385), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n853), .B2(new_n857), .ZN(G1341gat));
  NOR3_X1   g657(.A1(new_n836), .A2(new_n614), .A3(new_n668), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT117), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n614), .B1(new_n853), .B2(new_n668), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(KEYINPUT117), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1342gat));
  NOR3_X1   g663(.A1(new_n773), .A2(new_n388), .A3(new_n752), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n838), .A2(new_n852), .A3(new_n865), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n836), .B2(new_n752), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT118), .ZN(G1343gat));
  AOI21_X1  g670(.A(new_n349), .B1(new_n850), .B2(new_n851), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n666), .A2(new_n503), .A3(new_n728), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n719), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n666), .A2(new_n872), .A3(new_n503), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n768), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n287), .A2(G141gat), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n877), .A2(G141gat), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g681(.A(G148gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(new_n883), .A3(new_n645), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n669), .B1(new_n875), .B2(KEYINPUT119), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n872), .B2(KEYINPUT57), .ZN(new_n888));
  NOR4_X1   g687(.A1(new_n834), .A2(KEYINPUT120), .A3(new_n873), .A4(new_n349), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n349), .B1(new_n852), .B2(KEYINPUT121), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n834), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT57), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI221_X1 g693(.A(new_n886), .B1(KEYINPUT119), .B2(new_n875), .C1(new_n890), .C2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n885), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT59), .B(new_n883), .C1(new_n876), .C2(new_n645), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n884), .B1(new_n896), .B2(new_n897), .ZN(G1345gat));
  INV_X1    g697(.A(new_n876), .ZN(new_n899));
  OAI21_X1  g698(.A(G155gat), .B1(new_n899), .B2(new_n668), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n879), .A2(new_n299), .A3(new_n667), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n899), .B2(new_n752), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n491), .A2(new_n300), .A3(new_n581), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n878), .B2(new_n904), .ZN(G1347gat));
  NAND4_X1  g704(.A1(new_n835), .A2(new_n773), .A3(new_n659), .A4(new_n648), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT122), .Z(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n719), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n908), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT123), .B1(new_n908), .B2(G169gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n666), .A2(new_n834), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n728), .A2(new_n426), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n719), .A2(new_n350), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n909), .A2(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G1348gat));
  NAND3_X1  g714(.A1(new_n907), .A2(G176gat), .A3(new_n686), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n916), .A2(KEYINPUT124), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(KEYINPUT124), .ZN(new_n918));
  INV_X1    g717(.A(new_n913), .ZN(new_n919));
  AOI21_X1  g718(.A(G176gat), .B1(new_n919), .B2(new_n645), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(G1349gat));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT122), .ZN(new_n922));
  OAI21_X1  g721(.A(G183gat), .B1(new_n922), .B2(new_n668), .ZN(new_n923));
  OR3_X1    g722(.A1(new_n913), .A2(new_n362), .A3(new_n668), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(KEYINPUT125), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n925), .B(new_n927), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n919), .A2(new_n363), .A3(new_n581), .ZN(new_n929));
  OAI21_X1  g728(.A(G190gat), .B1(new_n922), .B2(new_n752), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  NOR3_X1   g732(.A1(new_n704), .A2(new_n349), .A3(new_n728), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n911), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n935), .A2(G197gat), .A3(new_n287), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT126), .Z(new_n937));
  NAND3_X1  g736(.A1(new_n648), .A2(new_n773), .A3(new_n503), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n844), .A2(new_n846), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n840), .B1(new_n287), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n752), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n667), .B1(new_n941), .B2(new_n829), .ZN(new_n942));
  OAI211_X1 g741(.A(KEYINPUT57), .B(new_n504), .C1(new_n942), .C2(new_n800), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT120), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n872), .A2(new_n887), .A3(KEYINPUT57), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n504), .B1(new_n834), .B2(new_n892), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n942), .A2(KEYINPUT121), .A3(new_n800), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n873), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n938), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n287), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n952), .ZN(G1352gat));
  NOR3_X1   g752(.A1(new_n935), .A2(G204gat), .A3(new_n669), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT62), .ZN(new_n955));
  OAI21_X1  g754(.A(G204gat), .B1(new_n951), .B2(new_n718), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1353gat));
  INV_X1    g756(.A(new_n935), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n306), .A3(new_n667), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n960));
  INV_X1    g759(.A(G211gat), .ZN(new_n961));
  AOI211_X1 g760(.A(new_n960), .B(new_n961), .C1(new_n950), .C2(new_n667), .ZN(new_n962));
  INV_X1    g761(.A(new_n938), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n667), .B(new_n963), .C1(new_n890), .C2(new_n894), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n959), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n968), .B(new_n959), .C1(new_n962), .C2(new_n965), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1354gat));
  OAI21_X1  g769(.A(G218gat), .B1(new_n951), .B2(new_n752), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n958), .A2(new_n307), .A3(new_n581), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1355gat));
endmodule


