

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732;

  INV_X1 U373 ( .A(G953), .ZN(n719) );
  XNOR2_X2 U374 ( .A(n584), .B(KEYINPUT22), .ZN(n589) );
  NOR2_X1 U375 ( .A1(n728), .A2(n732), .ZN(n548) );
  NOR2_X1 U376 ( .A1(n659), .A2(n660), .ZN(n598) );
  INV_X1 U377 ( .A(G125), .ZN(n458) );
  OR2_X1 U378 ( .A1(n656), .A2(n655), .ZN(n374) );
  AND2_X1 U379 ( .A1(n718), .A2(n711), .ZN(n656) );
  AND2_X1 U380 ( .A1(n610), .A2(n360), .ZN(n412) );
  XNOR2_X1 U381 ( .A(n419), .B(n418), .ZN(n729) );
  XNOR2_X1 U382 ( .A(n504), .B(n391), .ZN(n665) );
  AND2_X1 U383 ( .A1(n617), .A2(n500), .ZN(n465) );
  XNOR2_X1 U384 ( .A(n422), .B(n518), .ZN(n705) );
  XNOR2_X1 U385 ( .A(n470), .B(n428), .ZN(n716) );
  OR2_X2 U386 ( .A1(n589), .A2(n585), .ZN(n588) );
  NOR2_X1 U387 ( .A1(n589), .A2(n416), .ZN(n419) );
  XNOR2_X1 U388 ( .A(n424), .B(n705), .ZN(n617) );
  XNOR2_X1 U389 ( .A(n591), .B(KEYINPUT33), .ZN(n684) );
  AND2_X1 U390 ( .A1(n598), .A2(n523), .ZN(n591) );
  XNOR2_X1 U391 ( .A(n507), .B(n390), .ZN(n664) );
  INV_X1 U392 ( .A(KEYINPUT21), .ZN(n390) );
  INV_X1 U393 ( .A(n523), .ZN(n417) );
  XNOR2_X1 U394 ( .A(n484), .B(n483), .ZN(n556) );
  XNOR2_X1 U395 ( .A(n503), .B(KEYINPUT25), .ZN(n391) );
  NOR2_X1 U396 ( .A1(n650), .A2(n564), .ZN(n565) );
  AND2_X1 U397 ( .A1(n382), .A2(n380), .ZN(n435) );
  NAND2_X1 U398 ( .A1(n381), .A2(KEYINPUT81), .ZN(n380) );
  AND2_X1 U399 ( .A1(n353), .A2(n609), .ZN(n360) );
  XNOR2_X1 U400 ( .A(n454), .B(G134), .ZN(n485) );
  XNOR2_X1 U401 ( .A(n459), .B(n443), .ZN(n410) );
  XNOR2_X1 U402 ( .A(n442), .B(n409), .ZN(n408) );
  XNOR2_X1 U403 ( .A(G101), .B(G107), .ZN(n442) );
  XNOR2_X1 U404 ( .A(G146), .B(G104), .ZN(n409) );
  AND2_X1 U405 ( .A1(n528), .A2(n664), .ZN(n437) );
  NAND2_X1 U406 ( .A1(n585), .A2(n536), .ZN(n366) );
  INV_X1 U407 ( .A(KEYINPUT30), .ZN(n365) );
  XNOR2_X1 U408 ( .A(KEYINPUT3), .B(G119), .ZN(n460) );
  XOR2_X1 U409 ( .A(G101), .B(G116), .Z(n461) );
  XOR2_X1 U410 ( .A(G122), .B(G107), .Z(n490) );
  XNOR2_X1 U411 ( .A(n716), .B(n364), .ZN(n482) );
  XNOR2_X1 U412 ( .A(n471), .B(G143), .ZN(n364) );
  NOR2_X1 U413 ( .A1(n557), .A2(n677), .ZN(n532) );
  NOR2_X1 U414 ( .A1(n590), .A2(n684), .ZN(n592) );
  NAND2_X2 U415 ( .A1(n401), .A2(n398), .ZN(n540) );
  AND2_X1 U416 ( .A1(n403), .A2(n402), .ZN(n401) );
  NAND2_X1 U417 ( .A1(G469), .A2(n400), .ZN(n399) );
  XNOR2_X1 U418 ( .A(n663), .B(n356), .ZN(n523) );
  AND2_X1 U419 ( .A1(n680), .A2(n664), .ZN(n420) );
  XNOR2_X1 U420 ( .A(n427), .B(n425), .ZN(n702) );
  XNOR2_X1 U421 ( .A(n426), .B(n498), .ZN(n425) );
  XNOR2_X1 U422 ( .A(n716), .B(n385), .ZN(n427) );
  INV_X1 U423 ( .A(KEYINPUT125), .ZN(n393) );
  NAND2_X1 U424 ( .A1(n613), .A2(n657), .ZN(n615) );
  XNOR2_X1 U425 ( .A(n374), .B(KEYINPUT78), .ZN(n441) );
  INV_X1 U426 ( .A(n642), .ZN(n384) );
  XNOR2_X1 U427 ( .A(n550), .B(KEYINPUT103), .ZN(n597) );
  NOR2_X1 U428 ( .A1(n566), .A2(n435), .ZN(n434) );
  INV_X1 U429 ( .A(n597), .ZN(n676) );
  XNOR2_X1 U430 ( .A(KEYINPUT4), .B(KEYINPUT86), .ZN(n455) );
  XNOR2_X1 U431 ( .A(n415), .B(n413), .ZN(n453) );
  XNOR2_X1 U432 ( .A(KEYINPUT76), .B(KEYINPUT18), .ZN(n415) );
  NOR2_X1 U433 ( .A1(n414), .A2(G953), .ZN(n413) );
  INV_X1 U434 ( .A(G224), .ZN(n414) );
  NAND2_X1 U435 ( .A1(n362), .A2(n361), .ZN(n572) );
  INV_X1 U436 ( .A(n652), .ZN(n361) );
  XNOR2_X1 U437 ( .A(n432), .B(n363), .ZN(n362) );
  INV_X1 U438 ( .A(KEYINPUT48), .ZN(n363) );
  XNOR2_X1 U439 ( .A(n387), .B(n386), .ZN(n496) );
  INV_X1 U440 ( .A(KEYINPUT8), .ZN(n386) );
  NAND2_X1 U441 ( .A1(n719), .A2(G234), .ZN(n387) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n508) );
  OR2_X1 U443 ( .A1(G237), .A2(G902), .ZN(n468) );
  XNOR2_X1 U444 ( .A(n388), .B(KEYINPUT69), .ZN(n541) );
  OR2_X1 U445 ( .A1(n665), .A2(n389), .ZN(n388) );
  INV_X1 U446 ( .A(G902), .ZN(n400) );
  NAND2_X1 U447 ( .A1(n404), .A2(G902), .ZN(n402) );
  XOR2_X1 U448 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n502) );
  NOR2_X1 U449 ( .A1(G953), .A2(G237), .ZN(n517) );
  XNOR2_X1 U450 ( .A(n485), .B(n448), .ZN(n516) );
  XNOR2_X1 U451 ( .A(G137), .B(G131), .ZN(n447) );
  XNOR2_X1 U452 ( .A(G113), .B(G146), .ZN(n513) );
  XOR2_X1 U453 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n514) );
  NOR2_X2 U454 ( .A1(n572), .A2(n730), .ZN(n718) );
  XNOR2_X1 U455 ( .A(n411), .B(KEYINPUT45), .ZN(n711) );
  XNOR2_X1 U456 ( .A(n429), .B(KEYINPUT10), .ZN(n428) );
  INV_X1 U457 ( .A(G140), .ZN(n429) );
  XNOR2_X1 U458 ( .A(n499), .B(n497), .ZN(n426) );
  XOR2_X1 U459 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n499) );
  XNOR2_X1 U460 ( .A(G902), .B(KEYINPUT15), .ZN(n500) );
  XNOR2_X1 U461 ( .A(n410), .B(n408), .ZN(n446) );
  XNOR2_X1 U462 ( .A(n368), .B(KEYINPUT89), .ZN(n690) );
  AND2_X1 U463 ( .A1(n510), .A2(G952), .ZN(n368) );
  XNOR2_X1 U464 ( .A(n537), .B(KEYINPUT112), .ZN(n538) );
  XNOR2_X1 U465 ( .A(n366), .B(n365), .ZN(n376) );
  NOR2_X1 U466 ( .A1(n540), .A2(n436), .ZN(n529) );
  XNOR2_X1 U467 ( .A(n663), .B(n530), .ZN(n585) );
  NAND2_X1 U468 ( .A1(n701), .A2(G472), .ZN(n397) );
  INV_X1 U469 ( .A(n490), .ZN(n423) );
  XNOR2_X1 U470 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U471 ( .A(n373), .B(n372), .ZN(n562) );
  INV_X1 U472 ( .A(KEYINPUT36), .ZN(n372) );
  NOR2_X1 U473 ( .A1(n561), .A2(n551), .ZN(n373) );
  XNOR2_X1 U474 ( .A(n405), .B(KEYINPUT35), .ZN(n727) );
  INV_X1 U475 ( .A(n593), .ZN(n406) );
  INV_X1 U476 ( .A(KEYINPUT32), .ZN(n418) );
  NAND2_X1 U477 ( .A1(n354), .A2(n417), .ZN(n416) );
  OR2_X1 U478 ( .A1(n556), .A2(n549), .ZN(n647) );
  NOR2_X1 U479 ( .A1(n540), .A2(n660), .ZN(n601) );
  NAND2_X1 U480 ( .A1(n659), .A2(n605), .ZN(n632) );
  XNOR2_X1 U481 ( .A(n394), .B(n392), .ZN(n703) );
  NAND2_X1 U482 ( .A1(n701), .A2(G217), .ZN(n394) );
  INV_X1 U483 ( .A(KEYINPUT124), .ZN(n377) );
  INV_X1 U484 ( .A(KEYINPUT53), .ZN(n370) );
  XOR2_X1 U485 ( .A(n459), .B(n470), .Z(n352) );
  AND2_X1 U486 ( .A1(n606), .A2(n632), .ZN(n353) );
  NOR2_X1 U487 ( .A1(n665), .A2(n659), .ZN(n354) );
  INV_X1 U488 ( .A(G469), .ZN(n404) );
  NOR2_X1 U489 ( .A1(n589), .A2(n523), .ZN(n355) );
  XOR2_X1 U490 ( .A(KEYINPUT6), .B(KEYINPUT104), .Z(n356) );
  XOR2_X1 U491 ( .A(n631), .B(KEYINPUT62), .Z(n357) );
  NOR2_X1 U492 ( .A1(G952), .A2(n719), .ZN(n704) );
  XOR2_X1 U493 ( .A(n623), .B(KEYINPUT83), .Z(n358) );
  XNOR2_X2 U494 ( .A(n465), .B(n464), .ZN(n551) );
  XNOR2_X2 U495 ( .A(n359), .B(n583), .ZN(n590) );
  NAND2_X1 U496 ( .A1(n580), .A2(n581), .ZN(n359) );
  XNOR2_X1 U497 ( .A(n463), .B(n423), .ZN(n422) );
  NAND2_X1 U498 ( .A1(n466), .A2(n404), .ZN(n403) );
  XNOR2_X1 U499 ( .A(n717), .B(n450), .ZN(n466) );
  NOR2_X1 U500 ( .A1(n727), .A2(KEYINPUT44), .ZN(n594) );
  NAND2_X1 U501 ( .A1(n367), .A2(n544), .ZN(n545) );
  XNOR2_X1 U502 ( .A(n542), .B(n543), .ZN(n367) );
  NAND2_X1 U503 ( .A1(n528), .A2(n664), .ZN(n389) );
  XNOR2_X1 U504 ( .A(n369), .B(n630), .ZN(G60) );
  NAND2_X1 U505 ( .A1(n628), .A2(n629), .ZN(n369) );
  XNOR2_X1 U506 ( .A(n371), .B(n370), .ZN(G75) );
  NAND2_X1 U507 ( .A1(n697), .A2(n440), .ZN(n371) );
  NAND2_X1 U508 ( .A1(n541), .A2(n523), .ZN(n524) );
  INV_X1 U509 ( .A(n590), .ZN(n421) );
  XNOR2_X1 U510 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U511 ( .A(n375), .B(n457), .ZN(n424) );
  XNOR2_X1 U512 ( .A(n352), .B(n456), .ZN(n375) );
  NAND2_X1 U513 ( .A1(n376), .A2(n531), .ZN(n557) );
  XNOR2_X2 U514 ( .A(n521), .B(n522), .ZN(n663) );
  XNOR2_X1 U515 ( .A(n378), .B(n377), .ZN(G54) );
  NAND2_X1 U516 ( .A1(n430), .A2(n629), .ZN(n378) );
  XNOR2_X1 U517 ( .A(n379), .B(n358), .ZN(G51) );
  NAND2_X1 U518 ( .A1(n622), .A2(n629), .ZN(n379) );
  XNOR2_X1 U519 ( .A(n548), .B(KEYINPUT46), .ZN(n433) );
  INV_X1 U520 ( .A(n383), .ZN(n381) );
  XNOR2_X1 U521 ( .A(n383), .B(KEYINPUT47), .ZN(n382) );
  NAND2_X1 U522 ( .A1(n384), .A2(n676), .ZN(n383) );
  NAND2_X1 U523 ( .A1(n496), .A2(G221), .ZN(n385) );
  XNOR2_X1 U524 ( .A(n702), .B(n393), .ZN(n392) );
  NOR2_X4 U525 ( .A1(n615), .A2(n614), .ZN(n701) );
  XNOR2_X1 U526 ( .A(n395), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U527 ( .A1(n396), .A2(n629), .ZN(n395) );
  XNOR2_X1 U528 ( .A(n397), .B(n357), .ZN(n396) );
  OR2_X1 U529 ( .A1(n466), .A2(n399), .ZN(n398) );
  XNOR2_X2 U530 ( .A(n540), .B(n467), .ZN(n659) );
  NAND2_X1 U531 ( .A1(n407), .A2(n406), .ZN(n405) );
  XNOR2_X1 U532 ( .A(n592), .B(KEYINPUT34), .ZN(n407) );
  XNOR2_X1 U533 ( .A(n446), .B(n445), .ZN(n450) );
  NAND2_X1 U534 ( .A1(n611), .A2(n412), .ZN(n411) );
  NAND2_X1 U535 ( .A1(n729), .A2(n639), .ZN(n607) );
  NAND2_X1 U536 ( .A1(n421), .A2(n420), .ZN(n584) );
  XNOR2_X2 U537 ( .A(n458), .B(G146), .ZN(n470) );
  XNOR2_X1 U538 ( .A(n431), .B(n616), .ZN(n430) );
  NAND2_X1 U539 ( .A1(n701), .A2(G469), .ZN(n431) );
  NAND2_X1 U540 ( .A1(n434), .A2(n433), .ZN(n432) );
  NAND2_X1 U541 ( .A1(n665), .A2(n437), .ZN(n436) );
  NAND2_X1 U542 ( .A1(n665), .A2(n664), .ZN(n660) );
  AND2_X1 U543 ( .A1(n517), .A2(G210), .ZN(n438) );
  OR2_X1 U544 ( .A1(G953), .A2(n695), .ZN(n439) );
  NOR2_X1 U545 ( .A1(n696), .A2(n439), .ZN(n440) );
  XNOR2_X1 U546 ( .A(n447), .B(KEYINPUT4), .ZN(n448) );
  INV_X1 U547 ( .A(KEYINPUT75), .ZN(n444) );
  INV_X1 U548 ( .A(n684), .ZN(n693) );
  XNOR2_X1 U549 ( .A(n444), .B(G140), .ZN(n445) );
  XNOR2_X1 U550 ( .A(n518), .B(n438), .ZN(n519) );
  XNOR2_X1 U551 ( .A(n582), .B(KEYINPUT0), .ZN(n583) );
  XNOR2_X1 U552 ( .A(n520), .B(n519), .ZN(n631) );
  XNOR2_X1 U553 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U554 ( .A(n539), .B(n538), .ZN(n694) );
  XOR2_X1 U555 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n452) );
  XOR2_X2 U556 ( .A(KEYINPUT70), .B(G110), .Z(n459) );
  NAND2_X1 U557 ( .A1(G227), .A2(n719), .ZN(n443) );
  XNOR2_X2 U558 ( .A(G143), .B(G128), .ZN(n454) );
  INV_X1 U559 ( .A(n516), .ZN(n449) );
  XOR2_X1 U560 ( .A(KEYINPUT90), .B(n449), .Z(n717) );
  XNOR2_X1 U561 ( .A(n466), .B(KEYINPUT123), .ZN(n451) );
  XNOR2_X1 U562 ( .A(n452), .B(n451), .ZN(n616) );
  INV_X1 U563 ( .A(n500), .ZN(n613) );
  XOR2_X1 U564 ( .A(n453), .B(KEYINPUT17), .Z(n457) );
  XOR2_X1 U565 ( .A(n454), .B(n455), .Z(n456) );
  XNOR2_X1 U566 ( .A(n461), .B(n460), .ZN(n518) );
  XOR2_X2 U567 ( .A(G113), .B(G104), .Z(n478) );
  XOR2_X1 U568 ( .A(KEYINPUT72), .B(KEYINPUT16), .Z(n462) );
  XNOR2_X1 U569 ( .A(n478), .B(n462), .ZN(n463) );
  AND2_X1 U570 ( .A1(G210), .A2(n468), .ZN(n464) );
  INV_X1 U571 ( .A(n551), .ZN(n560) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(KEYINPUT65), .Z(n467) );
  INV_X1 U573 ( .A(n659), .ZN(n586) );
  NAND2_X1 U574 ( .A1(G214), .A2(n468), .ZN(n469) );
  XNOR2_X1 U575 ( .A(KEYINPUT88), .B(n469), .ZN(n536) );
  NAND2_X1 U576 ( .A1(n517), .A2(G214), .ZN(n471) );
  XOR2_X1 U577 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n473) );
  XNOR2_X1 U578 ( .A(G131), .B(KEYINPUT95), .ZN(n472) );
  XNOR2_X1 U579 ( .A(n473), .B(n472), .ZN(n477) );
  XOR2_X1 U580 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n475) );
  XNOR2_X1 U581 ( .A(KEYINPUT96), .B(KEYINPUT99), .ZN(n474) );
  XNOR2_X1 U582 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U583 ( .A(n477), .B(n476), .Z(n480) );
  XNOR2_X1 U584 ( .A(G122), .B(n478), .ZN(n479) );
  XNOR2_X1 U585 ( .A(n482), .B(n481), .ZN(n625) );
  NOR2_X1 U586 ( .A1(G902), .A2(n625), .ZN(n484) );
  XNOR2_X1 U587 ( .A(KEYINPUT13), .B(G475), .ZN(n483) );
  INV_X1 U588 ( .A(n485), .ZN(n489) );
  XOR2_X1 U589 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n487) );
  XNOR2_X1 U590 ( .A(G116), .B(KEYINPUT101), .ZN(n486) );
  XNOR2_X1 U591 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U592 ( .A(n489), .B(n488), .Z(n494) );
  XOR2_X1 U593 ( .A(n490), .B(KEYINPUT100), .Z(n492) );
  NAND2_X1 U594 ( .A1(G217), .A2(n496), .ZN(n491) );
  XNOR2_X1 U595 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U596 ( .A(n494), .B(n493), .ZN(n699) );
  NOR2_X1 U597 ( .A1(G902), .A2(n699), .ZN(n495) );
  XNOR2_X1 U598 ( .A(G478), .B(n495), .ZN(n549) );
  NAND2_X1 U599 ( .A1(n556), .A2(n549), .ZN(n644) );
  XOR2_X1 U600 ( .A(G137), .B(G128), .Z(n498) );
  XNOR2_X1 U601 ( .A(G119), .B(G110), .ZN(n497) );
  NOR2_X1 U602 ( .A1(n702), .A2(G902), .ZN(n504) );
  NAND2_X1 U603 ( .A1(G234), .A2(n500), .ZN(n501) );
  XNOR2_X1 U604 ( .A(n502), .B(n501), .ZN(n505) );
  NAND2_X1 U605 ( .A1(G217), .A2(n505), .ZN(n503) );
  NAND2_X1 U606 ( .A1(n505), .A2(G221), .ZN(n506) );
  XNOR2_X1 U607 ( .A(n506), .B(KEYINPUT92), .ZN(n507) );
  XNOR2_X1 U608 ( .A(n508), .B(KEYINPUT14), .ZN(n509) );
  XOR2_X1 U609 ( .A(KEYINPUT73), .B(n509), .Z(n510) );
  OR2_X1 U610 ( .A1(n690), .A2(G953), .ZN(n578) );
  NAND2_X1 U611 ( .A1(G902), .A2(n510), .ZN(n576) );
  NOR2_X1 U612 ( .A1(G900), .A2(n576), .ZN(n511) );
  NAND2_X1 U613 ( .A1(G953), .A2(n511), .ZN(n512) );
  NAND2_X1 U614 ( .A1(n578), .A2(n512), .ZN(n528) );
  XNOR2_X1 U615 ( .A(KEYINPUT71), .B(G472), .ZN(n522) );
  XNOR2_X1 U616 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U617 ( .A(n516), .B(n515), .ZN(n520) );
  NOR2_X1 U618 ( .A1(G902), .A2(n631), .ZN(n521) );
  NOR2_X1 U619 ( .A1(n644), .A2(n524), .ZN(n525) );
  NAND2_X1 U620 ( .A1(n536), .A2(n525), .ZN(n561) );
  NOR2_X1 U621 ( .A1(n586), .A2(n561), .ZN(n526) );
  XNOR2_X1 U622 ( .A(n526), .B(KEYINPUT43), .ZN(n527) );
  NOR2_X1 U623 ( .A1(n560), .A2(n527), .ZN(n652) );
  XNOR2_X1 U624 ( .A(KEYINPUT74), .B(n529), .ZN(n531) );
  INV_X1 U625 ( .A(KEYINPUT105), .ZN(n530) );
  XOR2_X1 U626 ( .A(n551), .B(KEYINPUT38), .Z(n677) );
  XNOR2_X1 U627 ( .A(n532), .B(KEYINPUT39), .ZN(n567) );
  NOR2_X1 U628 ( .A1(n644), .A2(n567), .ZN(n535) );
  XOR2_X1 U629 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n533) );
  XNOR2_X1 U630 ( .A(KEYINPUT110), .B(n533), .ZN(n534) );
  XNOR2_X1 U631 ( .A(n535), .B(n534), .ZN(n728) );
  INV_X1 U632 ( .A(n536), .ZN(n678) );
  NOR2_X1 U633 ( .A1(n678), .A2(n677), .ZN(n675) );
  INV_X1 U634 ( .A(n549), .ZN(n555) );
  NOR2_X1 U635 ( .A1(n556), .A2(n555), .ZN(n680) );
  NAND2_X1 U636 ( .A1(n675), .A2(n680), .ZN(n539) );
  XOR2_X1 U637 ( .A(KEYINPUT113), .B(KEYINPUT41), .Z(n537) );
  XNOR2_X1 U638 ( .A(n540), .B(KEYINPUT107), .ZN(n544) );
  XOR2_X1 U639 ( .A(KEYINPUT28), .B(KEYINPUT108), .Z(n543) );
  NAND2_X1 U640 ( .A1(n585), .A2(n541), .ZN(n542) );
  XNOR2_X1 U641 ( .A(n545), .B(KEYINPUT109), .ZN(n554) );
  NAND2_X1 U642 ( .A1(n694), .A2(n554), .ZN(n547) );
  INV_X1 U643 ( .A(KEYINPUT42), .ZN(n546) );
  XNOR2_X1 U644 ( .A(n547), .B(n546), .ZN(n732) );
  XNOR2_X1 U645 ( .A(KEYINPUT102), .B(n647), .ZN(n568) );
  NAND2_X1 U646 ( .A1(n644), .A2(n568), .ZN(n550) );
  NOR2_X1 U647 ( .A1(n551), .A2(n678), .ZN(n553) );
  XOR2_X1 U648 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n552) );
  XNOR2_X1 U649 ( .A(n553), .B(n552), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n554), .A2(n580), .ZN(n642) );
  NAND2_X1 U651 ( .A1(n556), .A2(n555), .ZN(n593) );
  NOR2_X1 U652 ( .A1(n557), .A2(n593), .ZN(n558) );
  NAND2_X1 U653 ( .A1(n560), .A2(n558), .ZN(n559) );
  XNOR2_X1 U654 ( .A(KEYINPUT106), .B(n559), .ZN(n731) );
  NOR2_X1 U655 ( .A1(n659), .A2(n562), .ZN(n650) );
  NAND2_X1 U656 ( .A1(KEYINPUT81), .A2(n597), .ZN(n563) );
  NOR2_X1 U657 ( .A1(n642), .A2(n563), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n731), .A2(n565), .ZN(n566) );
  OR2_X1 U659 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U660 ( .A(n569), .B(KEYINPUT114), .Z(n730) );
  INV_X1 U661 ( .A(KEYINPUT2), .ZN(n654) );
  NOR2_X1 U662 ( .A1(KEYINPUT77), .A2(n654), .ZN(n570) );
  NAND2_X1 U663 ( .A1(n718), .A2(n570), .ZN(n575) );
  NOR2_X1 U664 ( .A1(n730), .A2(n654), .ZN(n571) );
  NOR2_X1 U665 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U666 ( .A1(KEYINPUT77), .A2(n573), .ZN(n574) );
  NAND2_X1 U667 ( .A1(n575), .A2(n574), .ZN(n612) );
  INV_X1 U668 ( .A(n576), .ZN(n577) );
  NOR2_X1 U669 ( .A1(G898), .A2(n719), .ZN(n707) );
  NAND2_X1 U670 ( .A1(n577), .A2(n707), .ZN(n579) );
  NAND2_X1 U671 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U672 ( .A(KEYINPUT67), .B(KEYINPUT85), .ZN(n582) );
  OR2_X1 U673 ( .A1(n586), .A2(n665), .ZN(n587) );
  OR2_X1 U674 ( .A1(n588), .A2(n587), .ZN(n639) );
  XOR2_X1 U675 ( .A(n607), .B(KEYINPUT84), .Z(n596) );
  XNOR2_X1 U676 ( .A(n594), .B(KEYINPUT68), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n611) );
  XOR2_X1 U678 ( .A(KEYINPUT81), .B(n676), .Z(n604) );
  NAND2_X1 U679 ( .A1(n663), .A2(n598), .ZN(n670) );
  NOR2_X1 U680 ( .A1(n670), .A2(n590), .ZN(n599) );
  XNOR2_X1 U681 ( .A(n599), .B(KEYINPUT31), .ZN(n646) );
  NOR2_X1 U682 ( .A1(n663), .A2(n590), .ZN(n600) );
  NAND2_X1 U683 ( .A1(n601), .A2(n600), .ZN(n634) );
  NAND2_X1 U684 ( .A1(n646), .A2(n634), .ZN(n602) );
  XNOR2_X1 U685 ( .A(KEYINPUT94), .B(n602), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n606) );
  AND2_X1 U687 ( .A1(n665), .A2(n355), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n607), .A2(KEYINPUT44), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT64), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n727), .A2(KEYINPUT44), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n612), .A2(n711), .ZN(n657) );
  NOR2_X1 U692 ( .A1(n656), .A2(KEYINPUT2), .ZN(n614) );
  INV_X1 U693 ( .A(n704), .ZN(n629) );
  NAND2_X1 U694 ( .A1(n701), .A2(G210), .ZN(n621) );
  XNOR2_X1 U695 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n617), .B(KEYINPUT79), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n621), .B(n620), .ZN(n622) );
  INV_X1 U699 ( .A(KEYINPUT56), .ZN(n623) );
  INV_X1 U700 ( .A(KEYINPUT60), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n701), .A2(G475), .ZN(n627) );
  XOR2_X1 U702 ( .A(KEYINPUT59), .B(KEYINPUT87), .Z(n624) );
  XNOR2_X1 U703 ( .A(G101), .B(n632), .ZN(G3) );
  NOR2_X1 U704 ( .A1(n644), .A2(n634), .ZN(n633) );
  XOR2_X1 U705 ( .A(G104), .B(n633), .Z(G6) );
  NOR2_X1 U706 ( .A1(n647), .A2(n634), .ZN(n636) );
  XNOR2_X1 U707 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U709 ( .A(G107), .B(n637), .ZN(G9) );
  XOR2_X1 U710 ( .A(G110), .B(KEYINPUT115), .Z(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(G12) );
  XOR2_X1 U712 ( .A(G128), .B(KEYINPUT29), .Z(n641) );
  OR2_X1 U713 ( .A1(n647), .A2(n642), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G30) );
  NOR2_X1 U715 ( .A1(n644), .A2(n642), .ZN(n643) );
  XOR2_X1 U716 ( .A(G146), .B(n643), .Z(G48) );
  NOR2_X1 U717 ( .A1(n644), .A2(n646), .ZN(n645) );
  XOR2_X1 U718 ( .A(G113), .B(n645), .Z(G15) );
  NOR2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U720 ( .A(KEYINPUT116), .B(n648), .Z(n649) );
  XNOR2_X1 U721 ( .A(G116), .B(n649), .ZN(G18) );
  XNOR2_X1 U722 ( .A(G125), .B(n650), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n651), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U724 ( .A(G140), .B(n652), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(KEYINPUT117), .ZN(G42) );
  XOR2_X1 U726 ( .A(KEYINPUT80), .B(n654), .Z(n655) );
  NAND2_X1 U727 ( .A1(n657), .A2(n441), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n658), .B(KEYINPUT82), .ZN(n697) );
  XNOR2_X1 U729 ( .A(KEYINPUT52), .B(KEYINPUT121), .ZN(n689) );
  AND2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U731 ( .A(n661), .B(KEYINPUT50), .ZN(n662) );
  NOR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n669) );
  XOR2_X1 U733 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n667) );
  OR2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n671) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT51), .ZN(n673) );
  XNOR2_X1 U739 ( .A(n673), .B(KEYINPUT119), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n674), .A2(n694), .ZN(n687) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n683) );
  NAND2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U743 ( .A(KEYINPUT120), .B(n679), .ZN(n681) );
  NAND2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U746 ( .A1(n685), .A2(n693), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U748 ( .A(n689), .B(n688), .ZN(n691) );
  NOR2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U750 ( .A(KEYINPUT122), .B(n692), .ZN(n696) );
  AND2_X1 U751 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U752 ( .A1(G478), .A2(n701), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U754 ( .A1(n704), .A2(n700), .ZN(G63) );
  NOR2_X1 U755 ( .A1(n704), .A2(n703), .ZN(G66) );
  XOR2_X1 U756 ( .A(n705), .B(G110), .Z(n706) );
  NOR2_X1 U757 ( .A1(n707), .A2(n706), .ZN(n715) );
  NAND2_X1 U758 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n708), .B(KEYINPUT126), .ZN(n709) );
  XNOR2_X1 U760 ( .A(KEYINPUT61), .B(n709), .ZN(n710) );
  NAND2_X1 U761 ( .A1(G898), .A2(n710), .ZN(n713) );
  NAND2_X1 U762 ( .A1(n711), .A2(n719), .ZN(n712) );
  NAND2_X1 U763 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(G69) );
  XOR2_X1 U765 ( .A(n717), .B(n716), .Z(n721) );
  XOR2_X1 U766 ( .A(n718), .B(n721), .Z(n720) );
  NAND2_X1 U767 ( .A1(n720), .A2(n719), .ZN(n725) );
  XNOR2_X1 U768 ( .A(G227), .B(n721), .ZN(n722) );
  NAND2_X1 U769 ( .A1(n722), .A2(G900), .ZN(n723) );
  NAND2_X1 U770 ( .A1(G953), .A2(n723), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U772 ( .A(KEYINPUT127), .B(n726), .Z(G72) );
  XOR2_X1 U773 ( .A(G122), .B(n727), .Z(G24) );
  XOR2_X1 U774 ( .A(n728), .B(G131), .Z(G33) );
  XNOR2_X1 U775 ( .A(G119), .B(n729), .ZN(G21) );
  XOR2_X1 U776 ( .A(G134), .B(n730), .Z(G36) );
  XNOR2_X1 U777 ( .A(G143), .B(n731), .ZN(G45) );
  XOR2_X1 U778 ( .A(n732), .B(G137), .Z(G39) );
endmodule

