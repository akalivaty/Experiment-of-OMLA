//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n459), .B1(new_n448), .B2(new_n455), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT70), .B(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(new_n469), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n471), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OAI21_X1  g060(.A(G2104), .B1(new_n469), .B2(G112), .ZN(new_n486));
  NOR2_X1   g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT72), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n467), .A2(new_n482), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n486), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT71), .B1(new_n475), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n467), .A2(new_n493), .A3(new_n478), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(G136), .B2(new_n495), .ZN(G162));
  OAI21_X1  g071(.A(G138), .B1(new_n473), .B2(new_n474), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n497), .B2(new_n482), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n467), .A2(new_n469), .A3(new_n499), .A4(G138), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G126), .B(G2105), .C1(new_n473), .C2(new_n474), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n517), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n512), .B1(new_n526), .B2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(new_n516), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n520), .A2(new_n519), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n514), .A2(new_n515), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n534), .A2(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(new_n516), .A2(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n542), .B2(new_n523), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n511), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n543), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  INV_X1    g122(.A(new_n523), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT75), .B(G81), .Z(new_n549));
  AOI22_X1  g124(.A1(new_n548), .A2(new_n549), .B1(G43), .B2(new_n516), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n509), .A2(G56), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n511), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n550), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n554), .A2(new_n551), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n523), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n536), .A2(new_n509), .A3(KEYINPUT79), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n565), .A2(G91), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n565), .A2(KEYINPUT80), .A3(G91), .A4(new_n566), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(KEYINPUT81), .B(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n535), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n569), .A2(new_n570), .B1(G651), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g149(.A(KEYINPUT77), .B(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n516), .A2(G53), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n577));
  OAI211_X1 g152(.A(G53), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  INV_X1    g155(.A(new_n578), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n575), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n577), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n574), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  NAND3_X1  g160(.A1(new_n565), .A2(G87), .A3(new_n566), .ZN(new_n586));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n535), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n516), .B2(G49), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n535), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G48), .B2(new_n516), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n565), .A2(G86), .A3(new_n566), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n516), .A2(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n523), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n511), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n599), .A2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n565), .A2(G92), .A3(new_n566), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT10), .Z(new_n605));
  INV_X1    g180(.A(G54), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n532), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n516), .A2(KEYINPUT82), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n535), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n608), .A2(new_n609), .B1(G651), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n603), .B1(new_n615), .B2(G868), .ZN(G284));
  XOR2_X1   g191(.A(G284), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  INV_X1    g198(.A(new_n557), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n614), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n625), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n495), .A2(G135), .ZN(new_n630));
  INV_X1    g205(.A(new_n489), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G123), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n469), .A2(new_n633), .A3(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n469), .B2(G111), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(G2104), .A3(new_n636), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n630), .B(new_n632), .C1(new_n634), .C2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n467), .A2(new_n470), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT13), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n639), .A2(new_n640), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT86), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2430), .Z(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n653), .B(new_n657), .Z(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n660), .A2(new_n661), .A3(G14), .ZN(G401));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT87), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT88), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT89), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  INV_X1    g248(.A(new_n667), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n665), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n664), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n668), .B1(new_n676), .B2(new_n667), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n673), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n683), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G229));
  NAND2_X1  g273(.A1(new_n615), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G4), .B2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G1348), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G19), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n557), .B2(new_n704), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(G1341), .Z(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT90), .B(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G26), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n495), .A2(G140), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT94), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n469), .A2(G116), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n631), .A2(G128), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n711), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2067), .ZN(new_n722));
  OR3_X1    g297(.A1(new_n708), .A2(KEYINPUT95), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(KEYINPUT95), .B1(new_n708), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n704), .A2(G20), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT23), .Z(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G299), .B2(G16), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1956), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT24), .B(G34), .ZN(new_n729));
  AOI22_X1  g304(.A1(G160), .A2(G29), .B1(new_n709), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G2084), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(G2084), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n638), .B2(new_n709), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n704), .A2(G5), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G171), .B2(new_n704), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n731), .B(new_n733), .C1(G1961), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n495), .A2(G139), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n738), .B(new_n739), .C1(new_n469), .C2(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G33), .B(new_n741), .S(G29), .Z(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G2072), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n704), .A2(G21), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G168), .B2(new_n704), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G1966), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT98), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(G1966), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT96), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n736), .A2(new_n743), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT31), .B(G11), .ZN(new_n751));
  INV_X1    g326(.A(G28), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n752), .B2(KEYINPUT30), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(KEYINPUT97), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(KEYINPUT97), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(KEYINPUT30), .B2(new_n752), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n751), .B1(new_n754), .B2(new_n756), .C1(new_n735), .C2(G1961), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G105), .B2(new_n470), .ZN(new_n762));
  INV_X1    g337(.A(G129), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n489), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n495), .B2(G141), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(new_n720), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n720), .B2(G32), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n757), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n709), .A2(G27), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT99), .Z(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G164), .B2(new_n709), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(KEYINPUT100), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(KEYINPUT100), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n767), .A2(new_n768), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n769), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n709), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(G35), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G162), .B2(new_n779), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT29), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2090), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n750), .A2(new_n778), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n723), .A2(new_n724), .A3(new_n728), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n704), .A2(G23), .ZN(new_n786));
  INV_X1    g361(.A(G288), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n704), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n788), .B(new_n789), .Z(new_n790));
  MUX2_X1   g365(.A(G6), .B(G305), .S(G16), .Z(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G22), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G166), .B2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n793), .B1(G1971), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n790), .B(new_n796), .C1(G1971), .C2(new_n795), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT34), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n779), .A2(G25), .ZN(new_n799));
  OAI221_X1 g374(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n469), .C2(G107), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT91), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n495), .A2(G131), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n631), .A2(G119), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n799), .B1(new_n809), .B2(new_n779), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT93), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n798), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n704), .A2(G24), .ZN(new_n815));
  INV_X1    g390(.A(G290), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n704), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G1986), .Z(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n811), .B2(new_n812), .ZN(new_n819));
  OR3_X1    g394(.A1(new_n814), .A2(KEYINPUT36), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT36), .B1(new_n814), .B2(new_n819), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n785), .B1(new_n820), .B2(new_n821), .ZN(G311));
  INV_X1    g397(.A(G311), .ZN(G150));
  NAND2_X1  g398(.A1(new_n516), .A2(G55), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(new_n523), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n511), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT37), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n614), .A2(new_n622), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n829), .A2(KEYINPUT102), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n829), .A2(KEYINPUT102), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n624), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n557), .A2(KEYINPUT102), .A3(new_n829), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n835), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n830), .B1(new_n842), .B2(KEYINPUT39), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n832), .B1(new_n843), .B2(new_n844), .ZN(G145));
  NAND2_X1  g420(.A1(new_n495), .A2(G142), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n631), .A2(G130), .ZN(new_n847));
  OAI221_X1 g422(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n808), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n502), .A2(new_n505), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n502), .B2(new_n505), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n498), .A2(new_n855), .A3(new_n500), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n498), .B2(new_n500), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n741), .B(new_n858), .Z(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n850), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n850), .A2(new_n860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n718), .B(new_n765), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n643), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n861), .A2(new_n865), .A3(new_n862), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G160), .B(G162), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n638), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n871), .B2(new_n869), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g449(.A(G288), .B(KEYINPUT107), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G305), .ZN(new_n876));
  XNOR2_X1  g451(.A(G303), .B(new_n816), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT42), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n840), .B(new_n627), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n615), .A2(G299), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n619), .A2(new_n614), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n881), .A2(KEYINPUT105), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(KEYINPUT41), .ZN(new_n887));
  XOR2_X1   g462(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n888));
  NOR2_X1   g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n881), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT105), .B1(new_n881), .B2(new_n885), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n880), .B1(new_n892), .B2(KEYINPUT108), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(KEYINPUT108), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n880), .A2(new_n892), .A3(KEYINPUT108), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G868), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n829), .A2(G868), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(G295));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n902), .A3(new_n900), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n625), .B1(new_n895), .B2(new_n896), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT109), .B1(new_n904), .B2(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(G331));
  OAI21_X1  g481(.A(G168), .B1(G301), .B2(KEYINPUT110), .ZN(new_n907));
  NAND2_X1  g482(.A1(G301), .A2(KEYINPUT110), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n907), .B(new_n908), .Z(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n840), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(new_n885), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n887), .A2(new_n889), .ZN(new_n913));
  INV_X1    g488(.A(new_n910), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n912), .B(new_n878), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n878), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n913), .A2(new_n914), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(new_n911), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT43), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n915), .A2(new_n916), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n884), .A2(KEYINPUT41), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n910), .B(new_n924), .C1(new_n885), .C2(new_n888), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n878), .B1(new_n912), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n921), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n923), .B1(new_n917), .B2(new_n920), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n922), .A2(KEYINPUT43), .A3(new_n926), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n928), .B1(new_n931), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT45), .B1(new_n858), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n471), .A2(G40), .A3(new_n483), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G2067), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n718), .B(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT111), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n939), .B2(new_n765), .ZN(new_n940));
  INV_X1    g515(.A(G1996), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n936), .A2(G1996), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n765), .ZN(new_n945));
  INV_X1    g520(.A(new_n936), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n809), .A2(new_n812), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n809), .A2(new_n812), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n936), .A2(G1986), .A3(G290), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT48), .Z(new_n952));
  NAND4_X1  g527(.A1(new_n943), .A2(new_n945), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n944), .B(KEYINPUT46), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n940), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n955), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n947), .B(KEYINPUT127), .Z(new_n961));
  NAND3_X1  g536(.A1(new_n943), .A2(new_n945), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n719), .A2(new_n937), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n936), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n501), .B2(new_n506), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  OR3_X1    g543(.A1(new_n967), .A2(KEYINPUT113), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT113), .B1(new_n967), .B2(new_n968), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n471), .A2(G40), .A3(new_n483), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(G2084), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n497), .A2(new_n482), .A3(KEYINPUT4), .ZN(new_n974));
  INV_X1    g549(.A(G138), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n465), .B2(new_n466), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n499), .B1(new_n976), .B2(new_n469), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT103), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n498), .A2(new_n500), .A3(new_n855), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n980), .B2(new_n854), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT112), .B1(new_n981), .B2(new_n968), .ZN(new_n982));
  AND4_X1   g557(.A1(KEYINPUT112), .A2(new_n858), .A3(new_n968), .A4(new_n933), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n971), .B(new_n973), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1966), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n507), .A2(new_n933), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n935), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n934), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT118), .B(new_n985), .C1(new_n934), .C2(new_n988), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n984), .A2(G168), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n993), .A2(G8), .ZN(new_n994));
  INV_X1    g569(.A(new_n984), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n991), .A2(new_n992), .ZN(new_n996));
  OAI21_X1  g571(.A(G286), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n966), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(G8), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(KEYINPUT51), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT62), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n991), .A2(new_n992), .ZN(new_n1002));
  AOI21_X1  g577(.A(G168), .B1(new_n1002), .B2(new_n984), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT51), .B1(new_n1003), .B2(new_n999), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n994), .A2(new_n966), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT62), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n971), .B(new_n935), .C1(new_n982), .C2(new_n983), .ZN(new_n1008));
  INV_X1    g583(.A(G1961), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n858), .A2(KEYINPUT45), .A3(new_n933), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n972), .B1(new_n986), .B2(new_n987), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n773), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1008), .A2(new_n1009), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n934), .A2(new_n988), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(G2078), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(G301), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n858), .A2(new_n935), .A3(new_n933), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(G1981), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n594), .A2(new_n595), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n516), .A2(G48), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n536), .A2(new_n509), .A3(G86), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1023), .B(new_n1024), .C1(new_n1025), .C2(new_n511), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G1981), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1022), .A2(new_n1027), .A3(KEYINPUT49), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT115), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1022), .A2(new_n1027), .A3(new_n1032), .A4(KEYINPUT49), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1020), .A2(new_n1029), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n586), .A2(G1976), .A3(new_n589), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT114), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1020), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(G8), .A3(new_n1019), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1035), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1040), .A2(new_n1035), .A3(new_n1042), .A4(KEYINPUT117), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1971), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1008), .B2(G2090), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT55), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(G8), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n968), .B1(new_n858), .B2(new_n933), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n935), .B1(new_n986), .B2(KEYINPUT50), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1056), .A2(new_n1057), .A3(G2090), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1055), .B1(new_n1058), .B2(new_n1048), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G8), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1058), .A2(new_n1048), .A3(new_n1055), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1052), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AND4_X1   g637(.A1(new_n1018), .A2(new_n1047), .A3(new_n1054), .A4(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1001), .A2(new_n1007), .A3(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1035), .A2(new_n1038), .A3(new_n787), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1022), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1020), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1054), .B2(new_n1043), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G168), .A2(G8), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n1002), .B2(new_n984), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1047), .A2(new_n1062), .A3(new_n1054), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1050), .A2(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1052), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1043), .A2(new_n1072), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1054), .A3(new_n1070), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1068), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n569), .A2(new_n570), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n573), .A2(G651), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1079), .A2(new_n583), .A3(KEYINPUT57), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n574), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n583), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n581), .A2(new_n580), .A3(new_n575), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n1087));
  INV_X1    g662(.A(new_n579), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT119), .B(new_n1086), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n574), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1085), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1956), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1010), .A2(new_n1011), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n615), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1019), .A2(G2067), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(new_n1008), .B2(new_n701), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1085), .A2(new_n1105), .A3(new_n1095), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1083), .A2(new_n1084), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(new_n1105), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1102), .A2(new_n1104), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1101), .B(KEYINPUT61), .C1(new_n1109), .C2(new_n1106), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1010), .A2(new_n1011), .A3(new_n941), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1010), .A2(new_n1011), .A3(KEYINPUT122), .A4(new_n941), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1019), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n557), .ZN(new_n1124));
  NAND2_X1  g699(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1123), .A2(KEYINPUT123), .A3(KEYINPUT59), .A4(new_n557), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1104), .A2(KEYINPUT60), .A3(new_n614), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1116), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n614), .B1(new_n1104), .B2(KEYINPUT60), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(KEYINPUT60), .B2(new_n1104), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1110), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1010), .A2(new_n935), .A3(new_n1016), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1136), .A2(new_n934), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1014), .A2(new_n1135), .A3(G301), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1139), .A2(G301), .A3(new_n1140), .A4(new_n1137), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT125), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1134), .B(new_n1138), .C1(new_n1142), .C2(new_n1018), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1014), .A2(G301), .A3(new_n1017), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1014), .A2(new_n1137), .ZN(new_n1146));
  OAI211_X1 g721(.A(KEYINPUT54), .B(new_n1145), .C1(new_n1146), .C2(G301), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1047), .A2(new_n1054), .A3(new_n1062), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1143), .A2(new_n1144), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1064), .B(new_n1078), .C1(new_n1133), .C2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(G290), .B(G1986), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n946), .A2(new_n1151), .ZN(new_n1152));
  AND4_X1   g727(.A1(new_n1152), .A2(new_n943), .A3(new_n945), .A4(new_n950), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1150), .A2(KEYINPUT126), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT126), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n965), .B1(new_n1154), .B2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g731(.A(new_n461), .ZN(new_n1158));
  NOR4_X1   g732(.A1(G229), .A2(new_n1158), .A3(G401), .A4(G227), .ZN(new_n1159));
  OAI211_X1 g733(.A(new_n873), .B(new_n1159), .C1(new_n929), .C2(new_n930), .ZN(G225));
  INV_X1    g734(.A(G225), .ZN(G308));
endmodule


