

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n624, n625, n626, n627, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n656,
         n657, n658, n659, n660, n661, n662, n663, n665, n666, n667, n668,
         n669, n670, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762;

  INV_X1 U379 ( .A(n684), .ZN(n357) );
  INV_X1 U380 ( .A(n684), .ZN(n360) );
  INV_X1 U381 ( .A(n684), .ZN(n363) );
  INV_X1 U382 ( .A(n684), .ZN(n367) );
  BUF_X1 U383 ( .A(G122), .Z(n370) );
  NAND2_X1 U384 ( .A1(n620), .A2(n619), .ZN(n366) );
  AND2_X2 U385 ( .A1(n358), .A2(n357), .ZN(n630) );
  XNOR2_X1 U386 ( .A(n627), .B(n359), .ZN(n358) );
  INV_X1 U387 ( .A(n626), .ZN(n359) );
  AND2_X2 U388 ( .A1(n361), .A2(n360), .ZN(n657) );
  XNOR2_X1 U389 ( .A(n654), .B(n362), .ZN(n361) );
  INV_X1 U390 ( .A(n653), .ZN(n362) );
  AND2_X2 U391 ( .A1(n364), .A2(n363), .ZN(n665) );
  XNOR2_X1 U392 ( .A(n663), .B(n365), .ZN(n364) );
  INV_X1 U393 ( .A(n662), .ZN(n365) );
  AND2_X4 U394 ( .A1(n366), .A2(n622), .ZN(n674) );
  AND2_X2 U395 ( .A1(n368), .A2(n367), .ZN(n673) );
  XNOR2_X1 U396 ( .A(n670), .B(n369), .ZN(n368) );
  INV_X1 U397 ( .A(n669), .ZN(n369) );
  NOR2_X1 U398 ( .A1(n761), .A2(n762), .ZN(n580) );
  OR2_X2 U399 ( .A1(n709), .A2(n613), .ZN(n622) );
  NAND2_X1 U400 ( .A1(n635), .A2(n757), .ZN(n621) );
  XNOR2_X2 U401 ( .A(n544), .B(n409), .ZN(n585) );
  XNOR2_X2 U402 ( .A(n571), .B(n570), .ZN(n742) );
  XNOR2_X2 U403 ( .A(n449), .B(n448), .ZN(n750) );
  XNOR2_X2 U404 ( .A(n437), .B(n436), .ZN(n449) );
  XNOR2_X2 U405 ( .A(n385), .B(n391), .ZN(n531) );
  INV_X1 U406 ( .A(n718), .ZN(n573) );
  OR2_X1 U407 ( .A1(n625), .A2(G902), .ZN(n474) );
  BUF_X1 U408 ( .A(n621), .Z(n709) );
  NOR2_X1 U409 ( .A1(n704), .A2(n599), .ZN(n601) );
  XNOR2_X1 U410 ( .A(G110), .B(KEYINPUT16), .ZN(n392) );
  OR2_X2 U411 ( .A1(n549), .A2(n498), .ZN(n712) );
  XNOR2_X2 U412 ( .A(n371), .B(KEYINPUT0), .ZN(n516) );
  NOR2_X2 U413 ( .A1(n585), .A2(n416), .ZN(n371) );
  BUF_X1 U414 ( .A(n641), .Z(n372) );
  XNOR2_X2 U415 ( .A(n388), .B(n387), .ZN(n544) );
  XNOR2_X1 U416 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U417 ( .A(n750), .B(G146), .ZN(n472) );
  NAND2_X1 U418 ( .A1(n377), .A2(n713), .ZN(n509) );
  NAND2_X1 U419 ( .A1(n531), .A2(n390), .ZN(n540) );
  INV_X1 U420 ( .A(KEYINPUT71), .ZN(n390) );
  XNOR2_X1 U421 ( .A(G131), .B(KEYINPUT4), .ZN(n448) );
  XNOR2_X1 U422 ( .A(n428), .B(n427), .ZN(n668) );
  XNOR2_X1 U423 ( .A(n426), .B(n374), .ZN(n427) );
  XNOR2_X1 U424 ( .A(G107), .B(G110), .ZN(n455) );
  XNOR2_X1 U425 ( .A(G101), .B(G104), .ZN(n456) );
  OR2_X1 U426 ( .A1(n661), .A2(G902), .ZN(n461) );
  INV_X1 U427 ( .A(G237), .ZN(n405) );
  NOR2_X1 U428 ( .A1(n536), .A2(KEYINPUT44), .ZN(n535) );
  XOR2_X1 U429 ( .A(KEYINPUT12), .B(G143), .Z(n425) );
  XNOR2_X1 U430 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n398) );
  NAND2_X1 U431 ( .A1(G234), .A2(G237), .ZN(n410) );
  XNOR2_X1 U432 ( .A(G475), .B(KEYINPUT13), .ZN(n429) );
  INV_X1 U433 ( .A(KEYINPUT81), .ZN(n387) );
  XNOR2_X1 U434 ( .A(G101), .B(G113), .ZN(n395) );
  XNOR2_X1 U435 ( .A(KEYINPUT3), .B(G119), .ZN(n394) );
  XNOR2_X1 U436 ( .A(G119), .B(G128), .ZN(n475) );
  XNOR2_X1 U437 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n566) );
  XNOR2_X1 U438 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U439 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U440 ( .A(n472), .B(n373), .ZN(n661) );
  XNOR2_X1 U441 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X1 U442 ( .A1(n450), .A2(G952), .ZN(n684) );
  INV_X1 U443 ( .A(KEYINPUT35), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n497), .B(KEYINPUT32), .ZN(n632) );
  NAND2_X1 U445 ( .A1(n515), .A2(n514), .ZN(n633) );
  INV_X1 U446 ( .A(KEYINPUT80), .ZN(n512) );
  XOR2_X1 U447 ( .A(n458), .B(n457), .Z(n373) );
  NAND2_X1 U448 ( .A1(G214), .A2(n463), .ZN(n374) );
  NOR2_X1 U449 ( .A1(n496), .A2(n551), .ZN(n375) );
  XOR2_X1 U450 ( .A(KEYINPUT74), .B(KEYINPUT22), .Z(n376) );
  NAND2_X1 U451 ( .A1(n408), .A2(G214), .ZN(n726) );
  NAND2_X1 U452 ( .A1(n377), .A2(n375), .ZN(n497) );
  XNOR2_X2 U453 ( .A(n447), .B(n376), .ZN(n377) );
  NAND2_X1 U454 ( .A1(n378), .A2(n543), .ZN(n380) );
  NAND2_X1 U455 ( .A1(n537), .A2(KEYINPUT64), .ZN(n378) );
  XNOR2_X2 U456 ( .A(n379), .B(KEYINPUT45), .ZN(n635) );
  NAND2_X2 U457 ( .A1(n381), .A2(n380), .ZN(n379) );
  NOR2_X2 U458 ( .A1(n382), .A2(n535), .ZN(n381) );
  NAND2_X1 U459 ( .A1(n384), .A2(n534), .ZN(n382) );
  INV_X1 U460 ( .A(n532), .ZN(n541) );
  NAND2_X1 U461 ( .A1(n532), .A2(n383), .ZN(n536) );
  INV_X1 U462 ( .A(n540), .ZN(n383) );
  AND2_X2 U463 ( .A1(n647), .A2(n632), .ZN(n532) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n565) );
  NAND2_X1 U465 ( .A1(n533), .A2(KEYINPUT71), .ZN(n384) );
  NAND2_X1 U466 ( .A1(n386), .A2(n583), .ZN(n385) );
  XNOR2_X1 U467 ( .A(n505), .B(n504), .ZN(n386) );
  NOR2_X2 U468 ( .A1(n565), .A2(n389), .ZN(n388) );
  INV_X1 U469 ( .A(n726), .ZN(n389) );
  XNOR2_X1 U470 ( .A(n531), .B(n370), .ZN(G24) );
  BUF_X1 U471 ( .A(n674), .Z(n679) );
  XNOR2_X1 U472 ( .A(n430), .B(n429), .ZN(n524) );
  INV_X4 U473 ( .A(G953), .ZN(n450) );
  XNOR2_X1 U474 ( .A(n513), .B(n512), .ZN(n515) );
  XNOR2_X2 U475 ( .A(G104), .B(G122), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n419), .B(n392), .ZN(n393) );
  XNOR2_X1 U477 ( .A(G107), .B(G116), .ZN(n438) );
  XNOR2_X1 U478 ( .A(n393), .B(n438), .ZN(n396) );
  XNOR2_X1 U479 ( .A(n395), .B(n394), .ZN(n467) );
  XNOR2_X1 U480 ( .A(n396), .B(n467), .ZN(n641) );
  NAND2_X1 U481 ( .A1(n450), .A2(G224), .ZN(n397) );
  XNOR2_X1 U482 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U483 ( .A(G146), .B(G125), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n399), .B(n422), .ZN(n402) );
  XNOR2_X2 U485 ( .A(G143), .B(G128), .ZN(n437) );
  XNOR2_X1 U486 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n400) );
  XNOR2_X1 U487 ( .A(n437), .B(n400), .ZN(n401) );
  XNOR2_X1 U488 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U489 ( .A(n641), .B(n403), .ZN(n650) );
  XNOR2_X1 U490 ( .A(G902), .B(KEYINPUT15), .ZN(n616) );
  INV_X1 U491 ( .A(n616), .ZN(n404) );
  NOR2_X1 U492 ( .A1(n650), .A2(n404), .ZN(n407) );
  INV_X1 U493 ( .A(G902), .ZN(n487) );
  NAND2_X1 U494 ( .A1(n487), .A2(n405), .ZN(n408) );
  AND2_X1 U495 ( .A1(n408), .A2(G210), .ZN(n406) );
  XNOR2_X1 U496 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n409) );
  XNOR2_X1 U497 ( .A(KEYINPUT14), .B(n410), .ZN(n411) );
  NAND2_X1 U498 ( .A1(G952), .A2(n411), .ZN(n740) );
  NOR2_X1 U499 ( .A1(G953), .A2(n740), .ZN(n547) );
  NAND2_X1 U500 ( .A1(G902), .A2(n411), .ZN(n545) );
  NOR2_X1 U501 ( .A1(G898), .A2(n450), .ZN(n412) );
  XNOR2_X1 U502 ( .A(KEYINPUT85), .B(n412), .ZN(n642) );
  NOR2_X1 U503 ( .A1(n545), .A2(n642), .ZN(n413) );
  OR2_X1 U504 ( .A1(n547), .A2(n413), .ZN(n415) );
  INV_X1 U505 ( .A(KEYINPUT86), .ZN(n414) );
  XNOR2_X1 U506 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U507 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n418) );
  XNOR2_X1 U508 ( .A(G140), .B(KEYINPUT95), .ZN(n417) );
  XNOR2_X1 U509 ( .A(n418), .B(n417), .ZN(n421) );
  XOR2_X1 U510 ( .A(KEYINPUT11), .B(n419), .Z(n420) );
  XNOR2_X1 U511 ( .A(n421), .B(n420), .ZN(n423) );
  XNOR2_X1 U512 ( .A(n422), .B(KEYINPUT10), .ZN(n485) );
  XNOR2_X1 U513 ( .A(n423), .B(n485), .ZN(n428) );
  XNOR2_X1 U514 ( .A(G113), .B(G131), .ZN(n424) );
  XNOR2_X1 U515 ( .A(n425), .B(n424), .ZN(n426) );
  NOR2_X2 U516 ( .A1(G953), .A2(G237), .ZN(n463) );
  NOR2_X1 U517 ( .A1(G902), .A2(n668), .ZN(n430) );
  INV_X1 U518 ( .A(n524), .ZN(n506) );
  XOR2_X1 U519 ( .A(KEYINPUT9), .B(KEYINPUT98), .Z(n432) );
  XNOR2_X1 U520 ( .A(n370), .B(KEYINPUT7), .ZN(n431) );
  XNOR2_X1 U521 ( .A(n432), .B(n431), .ZN(n435) );
  NAND2_X1 U522 ( .A1(G234), .A2(n450), .ZN(n433) );
  XOR2_X1 U523 ( .A(KEYINPUT8), .B(n433), .Z(n481) );
  NAND2_X1 U524 ( .A1(G217), .A2(n481), .ZN(n434) );
  XNOR2_X1 U525 ( .A(n435), .B(n434), .ZN(n441) );
  INV_X1 U526 ( .A(G134), .ZN(n436) );
  XNOR2_X1 U527 ( .A(n438), .B(KEYINPUT97), .ZN(n439) );
  XNOR2_X1 U528 ( .A(n449), .B(n439), .ZN(n440) );
  XNOR2_X1 U529 ( .A(n441), .B(n440), .ZN(n681) );
  NAND2_X1 U530 ( .A1(n681), .A2(n487), .ZN(n442) );
  XNOR2_X1 U531 ( .A(n442), .B(G478), .ZN(n526) );
  INV_X1 U532 ( .A(n526), .ZN(n443) );
  NAND2_X1 U533 ( .A1(n506), .A2(n443), .ZN(n729) );
  NAND2_X1 U534 ( .A1(n616), .A2(G234), .ZN(n444) );
  XNOR2_X1 U535 ( .A(n444), .B(KEYINPUT20), .ZN(n488) );
  AND2_X1 U536 ( .A1(n488), .A2(G221), .ZN(n445) );
  XNOR2_X1 U537 ( .A(n445), .B(KEYINPUT21), .ZN(n710) );
  INV_X1 U538 ( .A(n710), .ZN(n498) );
  NOR2_X1 U539 ( .A1(n729), .A2(n498), .ZN(n446) );
  NAND2_X1 U540 ( .A1(n516), .A2(n446), .ZN(n447) );
  NAND2_X1 U541 ( .A1(n450), .A2(G227), .ZN(n451) );
  XNOR2_X1 U542 ( .A(n451), .B(KEYINPUT87), .ZN(n454) );
  INV_X1 U543 ( .A(G140), .ZN(n452) );
  XNOR2_X1 U544 ( .A(n452), .B(G137), .ZN(n484) );
  INV_X1 U545 ( .A(n484), .ZN(n453) );
  XNOR2_X1 U546 ( .A(n454), .B(n453), .ZN(n458) );
  XNOR2_X1 U547 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U548 ( .A(KEYINPUT69), .ZN(n459) );
  XNOR2_X1 U549 ( .A(n459), .B(G469), .ZN(n460) );
  XNOR2_X2 U550 ( .A(n461), .B(n460), .ZN(n576) );
  INV_X1 U551 ( .A(KEYINPUT1), .ZN(n462) );
  XNOR2_X2 U552 ( .A(n576), .B(n462), .ZN(n713) );
  XNOR2_X1 U553 ( .A(n509), .B(KEYINPUT101), .ZN(n494) );
  XOR2_X1 U554 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n465) );
  NAND2_X1 U555 ( .A1(n463), .A2(G210), .ZN(n464) );
  XNOR2_X1 U556 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U557 ( .A(n466), .B(KEYINPUT92), .Z(n470) );
  XNOR2_X1 U558 ( .A(G137), .B(G116), .ZN(n468) );
  XNOR2_X1 U559 ( .A(n467), .B(n468), .ZN(n469) );
  XNOR2_X1 U560 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U561 ( .A(n472), .B(n471), .ZN(n625) );
  INV_X1 U562 ( .A(G472), .ZN(n473) );
  XNOR2_X2 U563 ( .A(n474), .B(n473), .ZN(n718) );
  XOR2_X1 U564 ( .A(KEYINPUT24), .B(G110), .Z(n476) );
  XNOR2_X1 U565 ( .A(n476), .B(n475), .ZN(n480) );
  XOR2_X1 U566 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n478) );
  XNOR2_X1 U567 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n477) );
  XNOR2_X1 U568 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U569 ( .A(n480), .B(n479), .Z(n483) );
  NAND2_X1 U570 ( .A1(G221), .A2(n481), .ZN(n482) );
  XNOR2_X1 U571 ( .A(n483), .B(n482), .ZN(n486) );
  XNOR2_X1 U572 ( .A(n485), .B(n484), .ZN(n752) );
  XNOR2_X1 U573 ( .A(n486), .B(n752), .ZN(n675) );
  NAND2_X1 U574 ( .A1(n675), .A2(n487), .ZN(n492) );
  XOR2_X1 U575 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n490) );
  NAND2_X1 U576 ( .A1(n488), .A2(G217), .ZN(n489) );
  XNOR2_X1 U577 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U578 ( .A(n492), .B(n491), .ZN(n549) );
  AND2_X1 U579 ( .A1(n718), .A2(n549), .ZN(n493) );
  NAND2_X1 U580 ( .A1(n494), .A2(n493), .ZN(n647) );
  OR2_X1 U581 ( .A1(n713), .A2(n514), .ZN(n495) );
  XNOR2_X1 U582 ( .A(n495), .B(KEYINPUT100), .ZN(n496) );
  XNOR2_X1 U583 ( .A(n718), .B(KEYINPUT6), .ZN(n551) );
  NOR2_X1 U584 ( .A1(n713), .A2(n712), .ZN(n499) );
  NAND2_X1 U585 ( .A1(n499), .A2(n551), .ZN(n502) );
  XNOR2_X1 U586 ( .A(KEYINPUT82), .B(KEYINPUT33), .ZN(n500) );
  XNOR2_X1 U587 ( .A(n500), .B(KEYINPUT70), .ZN(n501) );
  XNOR2_X1 U588 ( .A(n502), .B(n501), .ZN(n734) );
  NAND2_X1 U589 ( .A1(n734), .A2(n516), .ZN(n505) );
  XNOR2_X1 U590 ( .A(KEYINPUT76), .B(KEYINPUT34), .ZN(n503) );
  XNOR2_X1 U591 ( .A(n503), .B(KEYINPUT73), .ZN(n504) );
  NAND2_X1 U592 ( .A1(n524), .A2(n526), .ZN(n508) );
  INV_X1 U593 ( .A(KEYINPUT102), .ZN(n507) );
  XNOR2_X1 U594 ( .A(n508), .B(n507), .ZN(n583) );
  INV_X1 U595 ( .A(n509), .ZN(n511) );
  INV_X1 U596 ( .A(n551), .ZN(n510) );
  NAND2_X1 U597 ( .A1(n511), .A2(n510), .ZN(n513) );
  INV_X1 U598 ( .A(n549), .ZN(n514) );
  BUF_X1 U599 ( .A(n516), .Z(n517) );
  INV_X1 U600 ( .A(n713), .ZN(n602) );
  NOR2_X1 U601 ( .A1(n718), .A2(n712), .ZN(n518) );
  AND2_X1 U602 ( .A1(n602), .A2(n518), .ZN(n721) );
  NAND2_X1 U603 ( .A1(n517), .A2(n721), .ZN(n520) );
  INV_X1 U604 ( .A(KEYINPUT31), .ZN(n519) );
  XNOR2_X1 U605 ( .A(n520), .B(n519), .ZN(n700) );
  INV_X1 U606 ( .A(n712), .ZN(n521) );
  NAND2_X1 U607 ( .A1(n521), .A2(n576), .ZN(n522) );
  NOR2_X1 U608 ( .A1(n573), .A2(n522), .ZN(n523) );
  NAND2_X1 U609 ( .A1(n517), .A2(n523), .ZN(n688) );
  NAND2_X1 U610 ( .A1(n700), .A2(n688), .ZN(n529) );
  XOR2_X1 U611 ( .A(n524), .B(KEYINPUT96), .Z(n527) );
  NOR2_X1 U612 ( .A1(n527), .A2(n526), .ZN(n525) );
  XOR2_X1 U613 ( .A(n525), .B(KEYINPUT99), .Z(n558) );
  AND2_X1 U614 ( .A1(n527), .A2(n526), .ZN(n692) );
  NOR2_X1 U615 ( .A1(n558), .A2(n692), .ZN(n591) );
  XNOR2_X1 U616 ( .A(n591), .B(KEYINPUT77), .ZN(n528) );
  NAND2_X1 U617 ( .A1(n529), .A2(n528), .ZN(n530) );
  AND2_X1 U618 ( .A1(n633), .A2(n530), .ZN(n534) );
  NAND2_X1 U619 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U620 ( .A1(n536), .A2(KEYINPUT44), .ZN(n537) );
  INV_X1 U621 ( .A(KEYINPUT64), .ZN(n538) );
  NAND2_X1 U622 ( .A1(n538), .A2(KEYINPUT44), .ZN(n539) );
  NOR2_X1 U623 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U624 ( .A1(n542), .A2(n541), .ZN(n543) );
  BUF_X1 U625 ( .A(n544), .Z(n554) );
  OR2_X1 U626 ( .A1(n450), .A2(n545), .ZN(n546) );
  NOR2_X1 U627 ( .A1(G900), .A2(n546), .ZN(n548) );
  NOR2_X1 U628 ( .A1(n548), .A2(n547), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n549), .A2(n710), .ZN(n550) );
  NOR2_X1 U630 ( .A1(n561), .A2(n550), .ZN(n572) );
  AND2_X1 U631 ( .A1(n551), .A2(n572), .ZN(n552) );
  AND2_X1 U632 ( .A1(n558), .A2(n552), .ZN(n553) );
  XOR2_X1 U633 ( .A(KEYINPUT103), .B(n553), .Z(n604) );
  NAND2_X1 U634 ( .A1(n554), .A2(n604), .ZN(n556) );
  INV_X1 U635 ( .A(KEYINPUT36), .ZN(n555) );
  XNOR2_X1 U636 ( .A(n556), .B(n555), .ZN(n557) );
  AND2_X1 U637 ( .A1(n557), .A2(n602), .ZN(n704) );
  INV_X1 U638 ( .A(n558), .ZN(n686) );
  NAND2_X1 U639 ( .A1(n573), .A2(n726), .ZN(n559) );
  XNOR2_X1 U640 ( .A(KEYINPUT30), .B(n559), .ZN(n560) );
  INV_X1 U641 ( .A(n560), .ZN(n564) );
  NOR2_X1 U642 ( .A1(n712), .A2(n561), .ZN(n562) );
  AND2_X1 U643 ( .A1(n562), .A2(n576), .ZN(n563) );
  NAND2_X1 U644 ( .A1(n564), .A2(n563), .ZN(n581) );
  BUF_X1 U645 ( .A(n565), .Z(n606) );
  XOR2_X1 U646 ( .A(KEYINPUT38), .B(n606), .Z(n569) );
  NOR2_X1 U647 ( .A1(n581), .A2(n569), .ZN(n567) );
  XNOR2_X1 U648 ( .A(n567), .B(n566), .ZN(n608) );
  NOR2_X1 U649 ( .A1(n686), .A2(n608), .ZN(n568) );
  XNOR2_X1 U650 ( .A(n568), .B(KEYINPUT40), .ZN(n761) );
  INV_X1 U651 ( .A(n569), .ZN(n727) );
  NAND2_X1 U652 ( .A1(n727), .A2(n726), .ZN(n730) );
  NOR2_X1 U653 ( .A1(n730), .A2(n729), .ZN(n571) );
  XNOR2_X1 U654 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n570) );
  NAND2_X1 U655 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U656 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n574) );
  XNOR2_X1 U657 ( .A(n575), .B(n574), .ZN(n577) );
  NAND2_X1 U658 ( .A1(n577), .A2(n576), .ZN(n586) );
  NOR2_X1 U659 ( .A1(n742), .A2(n586), .ZN(n578) );
  XNOR2_X1 U660 ( .A(KEYINPUT42), .B(n578), .ZN(n762) );
  XOR2_X1 U661 ( .A(KEYINPUT46), .B(KEYINPUT79), .Z(n579) );
  XNOR2_X1 U662 ( .A(n580), .B(n579), .ZN(n598) );
  NOR2_X1 U663 ( .A1(n581), .A2(n606), .ZN(n582) );
  XNOR2_X1 U664 ( .A(n582), .B(KEYINPUT104), .ZN(n584) );
  NAND2_X1 U665 ( .A1(n584), .A2(n583), .ZN(n695) );
  NOR2_X1 U666 ( .A1(n586), .A2(n585), .ZN(n696) );
  INV_X1 U667 ( .A(n591), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n696), .A2(n590), .ZN(n587) );
  NAND2_X1 U669 ( .A1(KEYINPUT47), .A2(n587), .ZN(n588) );
  AND2_X1 U670 ( .A1(n695), .A2(n588), .ZN(n596) );
  NOR2_X1 U671 ( .A1(KEYINPUT77), .A2(KEYINPUT47), .ZN(n589) );
  NAND2_X1 U672 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n591), .A2(KEYINPUT77), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n594), .A2(n696), .ZN(n595) );
  AND2_X1 U676 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U678 ( .A(KEYINPUT48), .B(KEYINPUT68), .ZN(n600) );
  XNOR2_X1 U679 ( .A(n601), .B(n600), .ZN(n611) );
  NOR2_X1 U680 ( .A1(n602), .A2(n389), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n605), .B(KEYINPUT43), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n634) );
  INV_X1 U684 ( .A(n692), .ZN(n701) );
  NOR2_X1 U685 ( .A1(n608), .A2(n701), .ZN(n707) );
  INV_X1 U686 ( .A(n707), .ZN(n609) );
  AND2_X1 U687 ( .A1(n634), .A2(n609), .ZN(n610) );
  AND2_X2 U688 ( .A1(n611), .A2(n610), .ZN(n757) );
  INV_X1 U689 ( .A(n621), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n612), .A2(KEYINPUT78), .ZN(n614) );
  INV_X1 U691 ( .A(KEYINPUT2), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n615), .A2(n404), .ZN(n620) );
  NOR2_X1 U694 ( .A1(n621), .A2(n616), .ZN(n617) );
  NOR2_X1 U695 ( .A1(n617), .A2(KEYINPUT78), .ZN(n618) );
  INV_X1 U696 ( .A(n618), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n674), .A2(G472), .ZN(n627) );
  XOR2_X1 U698 ( .A(KEYINPUT107), .B(KEYINPUT62), .Z(n624) );
  INV_X1 U699 ( .A(KEYINPUT63), .ZN(n629) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(G57) );
  XOR2_X1 U701 ( .A(G119), .B(KEYINPUT127), .Z(n631) );
  XNOR2_X1 U702 ( .A(n632), .B(n631), .ZN(G21) );
  XNOR2_X1 U703 ( .A(n633), .B(G101), .ZN(G3) );
  XNOR2_X1 U704 ( .A(n634), .B(G140), .ZN(G42) );
  AND2_X1 U705 ( .A1(n635), .A2(n450), .ZN(n640) );
  NAND2_X1 U706 ( .A1(G224), .A2(G953), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n636), .B(KEYINPUT124), .ZN(n637) );
  XNOR2_X1 U708 ( .A(KEYINPUT61), .B(n637), .ZN(n638) );
  AND2_X1 U709 ( .A1(n638), .A2(G898), .ZN(n639) );
  NOR2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n646) );
  INV_X1 U711 ( .A(n642), .ZN(n643) );
  NOR2_X1 U712 ( .A1(n372), .A2(n643), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n644), .B(KEYINPUT125), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n646), .B(n645), .ZN(G69) );
  BUF_X1 U715 ( .A(n647), .Z(n648) );
  XNOR2_X1 U716 ( .A(G110), .B(KEYINPUT108), .ZN(n649) );
  XNOR2_X1 U717 ( .A(n648), .B(n649), .ZN(G12) );
  NAND2_X1 U718 ( .A1(n674), .A2(G210), .ZN(n654) );
  BUF_X1 U719 ( .A(n650), .Z(n652) );
  XOR2_X1 U720 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n651) );
  XOR2_X1 U721 ( .A(KEYINPUT117), .B(KEYINPUT56), .Z(n656) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(G51) );
  NAND2_X1 U723 ( .A1(n674), .A2(G469), .ZN(n663) );
  XOR2_X1 U724 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n659) );
  XNOR2_X1 U725 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n658) );
  XOR2_X1 U726 ( .A(n659), .B(n658), .Z(n660) );
  XNOR2_X1 U727 ( .A(n665), .B(KEYINPUT120), .ZN(G54) );
  NAND2_X1 U728 ( .A1(n674), .A2(G475), .ZN(n670) );
  XOR2_X1 U729 ( .A(KEYINPUT65), .B(KEYINPUT83), .Z(n666) );
  XNOR2_X1 U730 ( .A(n666), .B(KEYINPUT59), .ZN(n667) );
  XOR2_X1 U731 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n672) );
  XNOR2_X1 U732 ( .A(n673), .B(n672), .ZN(G60) );
  NAND2_X1 U733 ( .A1(n679), .A2(G217), .ZN(n677) );
  XNOR2_X1 U734 ( .A(n675), .B(KEYINPUT123), .ZN(n676) );
  XNOR2_X1 U735 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U736 ( .A1(n678), .A2(n684), .ZN(G66) );
  NAND2_X1 U737 ( .A1(n679), .A2(G478), .ZN(n683) );
  XNOR2_X1 U738 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n680) );
  XNOR2_X1 U739 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U740 ( .A(n683), .B(n682), .ZN(n685) );
  NOR2_X1 U741 ( .A1(n685), .A2(n684), .ZN(G63) );
  NOR2_X1 U742 ( .A1(n686), .A2(n688), .ZN(n687) );
  XOR2_X1 U743 ( .A(G104), .B(n687), .Z(G6) );
  NOR2_X1 U744 ( .A1(n701), .A2(n688), .ZN(n690) );
  XNOR2_X1 U745 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U747 ( .A(G107), .B(n691), .ZN(G9) );
  XOR2_X1 U748 ( .A(G128), .B(KEYINPUT29), .Z(n694) );
  NAND2_X1 U749 ( .A1(n692), .A2(n696), .ZN(n693) );
  XNOR2_X1 U750 ( .A(n694), .B(n693), .ZN(G30) );
  XNOR2_X1 U751 ( .A(G143), .B(n695), .ZN(G45) );
  XOR2_X1 U752 ( .A(G146), .B(KEYINPUT109), .Z(n698) );
  NAND2_X1 U753 ( .A1(n558), .A2(n696), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n698), .B(n697), .ZN(G48) );
  NOR2_X1 U755 ( .A1(n686), .A2(n700), .ZN(n699) );
  XOR2_X1 U756 ( .A(G113), .B(n699), .Z(G15) );
  NOR2_X1 U757 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U758 ( .A(KEYINPUT110), .B(n702), .Z(n703) );
  XNOR2_X1 U759 ( .A(G116), .B(n703), .ZN(G18) );
  XOR2_X1 U760 ( .A(KEYINPUT111), .B(KEYINPUT37), .Z(n706) );
  XNOR2_X1 U761 ( .A(n704), .B(G125), .ZN(n705) );
  XNOR2_X1 U762 ( .A(n706), .B(n705), .ZN(G27) );
  XOR2_X1 U763 ( .A(G134), .B(n707), .Z(n708) );
  XNOR2_X1 U764 ( .A(KEYINPUT112), .B(n708), .ZN(G36) );
  XNOR2_X1 U765 ( .A(n709), .B(KEYINPUT2), .ZN(n747) );
  NOR2_X1 U766 ( .A1(n514), .A2(n710), .ZN(n711) );
  XOR2_X1 U767 ( .A(KEYINPUT49), .B(n711), .Z(n717) );
  NAND2_X1 U768 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U769 ( .A(n714), .B(KEYINPUT113), .ZN(n715) );
  XNOR2_X1 U770 ( .A(KEYINPUT50), .B(n715), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n720), .B(KEYINPUT114), .ZN(n723) );
  INV_X1 U774 ( .A(n721), .ZN(n722) );
  NAND2_X1 U775 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U776 ( .A(KEYINPUT51), .B(n724), .ZN(n725) );
  NOR2_X1 U777 ( .A1(n742), .A2(n725), .ZN(n737) );
  NOR2_X1 U778 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U779 ( .A1(n729), .A2(n728), .ZN(n732) );
  NOR2_X1 U780 ( .A1(n591), .A2(n730), .ZN(n731) );
  NOR2_X1 U781 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U782 ( .A(KEYINPUT115), .B(n733), .Z(n735) );
  INV_X1 U783 ( .A(n734), .ZN(n741) );
  NOR2_X1 U784 ( .A1(n735), .A2(n741), .ZN(n736) );
  NOR2_X1 U785 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U786 ( .A(n738), .B(KEYINPUT52), .ZN(n739) );
  NOR2_X1 U787 ( .A1(n740), .A2(n739), .ZN(n745) );
  NOR2_X1 U788 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U789 ( .A(n743), .B(KEYINPUT116), .ZN(n744) );
  OR2_X1 U790 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U791 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U792 ( .A1(n748), .A2(G953), .ZN(n749) );
  XNOR2_X1 U793 ( .A(n749), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U794 ( .A(n750), .B(KEYINPUT87), .ZN(n751) );
  XOR2_X1 U795 ( .A(n752), .B(n751), .Z(n756) );
  XOR2_X1 U796 ( .A(KEYINPUT126), .B(n756), .Z(n753) );
  XNOR2_X1 U797 ( .A(G227), .B(n753), .ZN(n754) );
  NAND2_X1 U798 ( .A1(G900), .A2(n754), .ZN(n755) );
  NAND2_X1 U799 ( .A1(n755), .A2(G953), .ZN(n760) );
  XNOR2_X1 U800 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U801 ( .A1(n758), .A2(n450), .ZN(n759) );
  NAND2_X1 U802 ( .A1(n760), .A2(n759), .ZN(G72) );
  XOR2_X1 U803 ( .A(G131), .B(n761), .Z(G33) );
  XOR2_X1 U804 ( .A(G137), .B(n762), .Z(G39) );
endmodule

