//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1198, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AND2_X1   g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  XOR2_X1   g0017(.A(KEYINPUT65), .B(G244), .Z(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n205), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n211), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n214), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G50), .B(G68), .Z(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G274), .ZN(new_n243));
  NAND2_X1  g0043(.A1(G33), .A2(G41), .ZN(new_n244));
  AOI21_X1  g0044(.A(new_n243), .B1(new_n215), .B2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n215), .A2(new_n244), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n252), .B(new_n246), .C1(G41), .C2(G45), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G226), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n249), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G222), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n260), .B1(new_n205), .B2(new_n258), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n257), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n269), .A2(G179), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT8), .B(G58), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n272), .A2(new_n274), .B1(G150), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G20), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n204), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(new_n211), .B2(new_n273), .ZN(new_n280));
  NAND4_X1  g0080(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n265), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n246), .A2(G13), .A3(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n277), .A2(G1), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(G50), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n285), .A2(new_n202), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n283), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n269), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n270), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n283), .A2(KEYINPUT9), .A3(new_n289), .A4(new_n290), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n257), .A2(new_n267), .A3(G190), .A4(new_n268), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n269), .A2(G200), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n299), .A2(new_n300), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n302), .A2(new_n297), .A3(new_n301), .A4(new_n298), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n295), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G68), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n274), .A2(G77), .B1(G20), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n275), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n202), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT71), .B1(new_n310), .B2(new_n282), .ZN(new_n313));
  OR3_X1    g0113(.A1(new_n312), .A2(KEYINPUT11), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT11), .B1(new_n312), .B2(new_n313), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT72), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n284), .B2(G68), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT12), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n287), .A2(new_n307), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n286), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n314), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n258), .A2(G226), .A3(new_n259), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n266), .ZN(new_n327));
  OAI21_X1  g0127(.A(G274), .B1(new_n264), .B2(new_n265), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n247), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(G238), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n327), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(G169), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(G179), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n337), .B1(new_n336), .B2(G169), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n322), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n336), .A2(G200), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n333), .A2(G190), .A3(new_n335), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n321), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n280), .A2(new_n265), .A3(new_n281), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n284), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n347), .A2(new_n205), .A3(new_n287), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT15), .B(G87), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n274), .B1(G20), .B2(G77), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n272), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n346), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n284), .A2(G77), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n348), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n249), .B1(new_n254), .B2(new_n218), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n360));
  INV_X1    g0160(.A(G238), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n360), .B1(new_n208), .B2(new_n258), .C1(new_n261), .C2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n359), .B1(new_n362), .B2(new_n266), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n357), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n363), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n365), .A2(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n362), .A2(new_n266), .ZN(new_n370));
  INV_X1    g0170(.A(new_n359), .ZN(new_n371));
  AOI21_X1  g0171(.A(G169), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n357), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n373), .B2(KEYINPUT70), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT70), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n357), .B2(new_n372), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n368), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n306), .A2(new_n342), .A3(new_n345), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  INV_X1    g0179(.A(G58), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n307), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n381), .B2(new_n201), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n275), .A2(G159), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n258), .B2(G20), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT3), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(G33), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT7), .B(new_n277), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n307), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n385), .B1(new_n392), .B2(KEYINPUT73), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT73), .ZN(new_n394));
  AOI211_X1 g0194(.A(new_n394), .B(new_n307), .C1(new_n387), .C2(new_n391), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n379), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n392), .A2(new_n384), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n346), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n272), .A2(new_n288), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n347), .A2(new_n400), .B1(new_n284), .B2(new_n272), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G232), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n249), .B1(new_n254), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n258), .A2(G226), .A3(G1698), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n258), .A2(G223), .A3(new_n259), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n405), .B1(new_n266), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(new_n292), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n266), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n329), .B1(new_n330), .B2(G232), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n412), .A2(new_n413), .A3(G179), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n403), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n401), .B1(new_n396), .B2(new_n398), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n411), .A2(new_n414), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT18), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n412), .A2(new_n413), .A3(new_n366), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n410), .B2(G200), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n258), .A2(new_n386), .A3(G20), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n388), .A2(G33), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n428), .B2(new_n277), .ZN(new_n429));
  OAI21_X1  g0229(.A(G68), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n384), .B1(new_n430), .B2(new_n394), .ZN(new_n431));
  INV_X1    g0231(.A(new_n395), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT16), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n385), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n282), .B1(new_n434), .B2(new_n379), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n424), .B(new_n402), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n424), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(KEYINPUT74), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT74), .B1(new_n438), .B2(new_n439), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n422), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT75), .B1(new_n378), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n342), .A2(new_n377), .A3(new_n345), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT75), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT74), .ZN(new_n447));
  AND4_X1   g0247(.A1(KEYINPUT17), .A2(new_n399), .A3(new_n402), .A4(new_n424), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT17), .B1(new_n418), .B2(new_n424), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n421), .B1(new_n450), .B2(new_n440), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n445), .A2(new_n446), .A3(new_n451), .A4(new_n306), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n246), .A2(G33), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n346), .A2(G116), .A3(new_n284), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n285), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(G20), .B1(G33), .B2(G283), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n273), .A2(G97), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n458), .A2(new_n459), .B1(G20), .B2(new_n456), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n282), .A2(KEYINPUT20), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT20), .B1(new_n282), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n455), .B(new_n457), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n426), .A2(new_n427), .A3(G257), .A4(new_n259), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n426), .A2(new_n427), .A3(G264), .A4(G1698), .ZN(new_n465));
  INV_X1    g0265(.A(G303), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n258), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n266), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT76), .B1(new_n474), .B2(new_n328), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT5), .B(G41), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT76), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n245), .A2(new_n476), .A3(new_n477), .A4(new_n470), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n266), .B1(new_n470), .B2(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G270), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n468), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n463), .A2(new_n482), .A3(G169), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n463), .A2(new_n482), .A3(KEYINPUT80), .A4(G169), .ZN(new_n486));
  XOR2_X1   g0286(.A(KEYINPUT81), .B(KEYINPUT21), .Z(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n482), .A2(KEYINPUT21), .A3(G169), .ZN(new_n489));
  INV_X1    g0289(.A(G179), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n463), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n482), .A2(G200), .ZN(new_n493));
  INV_X1    g0293(.A(new_n463), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n494), .C1(new_n366), .C2(new_n482), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n488), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n426), .A2(new_n427), .A3(G257), .A4(G1698), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT85), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n258), .A2(KEYINPUT85), .A3(G257), .A4(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n426), .A2(new_n427), .A3(G250), .A4(new_n259), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G294), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n266), .B1(G264), .B2(new_n480), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n490), .A3(new_n479), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n480), .A2(G264), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n505), .B1(new_n500), .B2(new_n501), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n479), .B(new_n510), .C1(new_n511), .C2(new_n251), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n292), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT23), .B1(new_n277), .B2(G107), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT23), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n208), .A3(G20), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n277), .A2(G33), .A3(G116), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT83), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n426), .A2(new_n427), .A3(new_n277), .A4(G87), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT82), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n258), .A2(new_n277), .A3(G87), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n522), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT24), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n522), .A2(new_n531), .A3(new_n526), .A4(new_n528), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n346), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  XOR2_X1   g0333(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n534));
  NOR2_X1   g0334(.A1(new_n284), .A2(G107), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n286), .A2(new_n454), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(new_n208), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n509), .B(new_n513), .C1(new_n533), .C2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n426), .A2(new_n427), .A3(G238), .A4(new_n259), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n426), .A2(new_n427), .A3(G244), .A4(G1698), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n273), .C2(new_n456), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n266), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n246), .A2(G45), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT78), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n544), .B(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n251), .A2(G250), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n546), .A2(new_n547), .B1(new_n245), .B2(new_n470), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT79), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n543), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n543), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n292), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n543), .A2(new_n548), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT79), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n543), .A2(new_n548), .A3(new_n549), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n490), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n258), .A2(new_n277), .A3(G68), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n277), .B1(new_n325), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(G87), .B2(new_n209), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n273), .A2(new_n207), .A3(G20), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n557), .B(new_n560), .C1(KEYINPUT19), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n282), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n349), .A2(new_n285), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n564), .C1(new_n349), .C2(new_n537), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n552), .A2(new_n556), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n550), .B2(new_n551), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n554), .A2(G190), .A3(new_n555), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  INV_X1    g0369(.A(G87), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n537), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n567), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n539), .A2(new_n566), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT86), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n508), .A2(new_n575), .A3(new_n366), .A4(new_n479), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT86), .B1(new_n512), .B2(G190), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n512), .A2(new_n358), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n533), .A2(new_n538), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT6), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n582), .A2(new_n207), .A3(G107), .ZN(new_n583));
  XNOR2_X1  g0383(.A(G97), .B(G107), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n585), .A2(new_n277), .B1(new_n205), .B2(new_n309), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n208), .B1(new_n387), .B2(new_n391), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n282), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n286), .A2(G97), .A3(new_n454), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n284), .A2(G97), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G283), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n426), .A2(new_n427), .A3(G250), .A4(G1698), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n426), .A2(new_n427), .A3(G244), .A4(new_n259), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n266), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n475), .A2(new_n478), .B1(new_n480), .B2(G257), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n292), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n490), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n592), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT77), .B1(new_n601), .B2(G200), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT77), .ZN(new_n606));
  AOI211_X1 g0406(.A(new_n606), .B(new_n358), .C1(new_n599), .C2(new_n600), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n599), .A2(new_n600), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n592), .B1(G190), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n604), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n497), .A2(new_n574), .A3(new_n581), .A4(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n453), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n614), .B(KEYINPUT87), .ZN(G372));
  NAND3_X1  g0415(.A1(new_n566), .A2(new_n573), .A3(new_n604), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT26), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n553), .A2(new_n292), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n553), .A2(KEYINPUT88), .A3(new_n292), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n556), .A2(new_n620), .A3(new_n565), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n553), .A2(G200), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n568), .A2(new_n572), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n622), .A2(new_n604), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n617), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n488), .A2(new_n539), .A3(new_n492), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n622), .A2(new_n624), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n611), .A2(new_n628), .A3(new_n629), .A4(new_n581), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n453), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n374), .A2(new_n376), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n345), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n342), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n442), .B2(new_n441), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n422), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n303), .A2(new_n305), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n295), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n632), .A2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(G13), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n642), .A2(G1), .A3(G20), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT89), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n463), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n497), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n488), .A2(new_n492), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n650), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n539), .A2(new_n649), .ZN(new_n655));
  INV_X1    g0455(.A(new_n649), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n581), .B1(new_n580), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n657), .B2(new_n539), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n652), .A2(new_n649), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n539), .B2(new_n649), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n660), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n212), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G1), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n217), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT29), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n622), .A2(new_n604), .A3(new_n624), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT26), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n566), .A2(new_n573), .A3(new_n604), .A4(new_n625), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n622), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT91), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT92), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n630), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n604), .ZN(new_n681));
  INV_X1    g0481(.A(new_n592), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n609), .A2(G190), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n682), .B(new_n683), .C1(new_n605), .C2(new_n607), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n581), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n685), .A2(KEYINPUT92), .A3(new_n628), .A4(new_n629), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n674), .A2(KEYINPUT91), .A3(new_n622), .A4(new_n675), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n678), .A2(new_n680), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n672), .B1(new_n688), .B2(new_n656), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n468), .A2(new_n479), .A3(new_n481), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n609), .A2(new_n508), .A3(G179), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n554), .A2(new_n555), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n512), .A2(new_n601), .ZN(new_n696));
  AOI21_X1  g0496(.A(G179), .B1(new_n543), .B2(new_n548), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT90), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n697), .A2(new_n698), .A3(new_n482), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n697), .B2(new_n482), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n550), .A2(new_n551), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n510), .B1(new_n511), .B2(new_n251), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n601), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n702), .A2(new_n704), .A3(KEYINPUT30), .A4(new_n491), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n695), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n649), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n581), .A2(new_n681), .A3(new_n684), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n539), .A2(new_n566), .A3(new_n573), .ZN(new_n714));
  NOR4_X1   g0514(.A1(new_n713), .A2(new_n496), .A3(new_n714), .A4(new_n649), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n690), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g0517(.A(KEYINPUT29), .B(new_n649), .C1(new_n627), .C2(new_n630), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n689), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n671), .B1(new_n719), .B2(G1), .ZN(G364));
  NOR2_X1   g0520(.A1(new_n642), .A2(G20), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n246), .B1(new_n721), .B2(G45), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n666), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n653), .A2(G330), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n724), .B1(new_n725), .B2(new_n654), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT94), .Z(new_n730));
  OR2_X1    g0530(.A1(new_n653), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n277), .A2(new_n366), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n490), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G190), .ZN(new_n737));
  XNOR2_X1  g0537(.A(KEYINPUT33), .B(G317), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n735), .A2(G322), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT98), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n490), .A2(G200), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT97), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(new_n277), .A3(G190), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n743), .A2(new_n277), .A3(new_n366), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G283), .A2(new_n744), .B1(new_n745), .B2(G303), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n277), .A2(G190), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n733), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G311), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n428), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G179), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n750), .B1(G329), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n277), .B1(new_n751), .B2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n736), .A2(new_n366), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n756), .A2(G294), .B1(G326), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n740), .A2(new_n746), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n744), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n208), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n755), .A2(new_n207), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n761), .A2(new_n428), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n753), .A2(G159), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT32), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(G68), .B2(new_n737), .ZN(new_n766));
  INV_X1    g0566(.A(new_n745), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n570), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n763), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n748), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G58), .A2(new_n735), .B1(new_n771), .B2(G77), .ZN(new_n772));
  INV_X1    g0572(.A(new_n757), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n202), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT96), .Z(new_n775));
  OAI21_X1  g0575(.A(new_n759), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n265), .B1(G20), .B2(new_n292), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT95), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(KEYINPUT95), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n730), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n780), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n217), .A2(G45), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n665), .A2(new_n258), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n783), .B(new_n784), .C1(new_n238), .C2(new_n469), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n258), .A2(new_n212), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(KEYINPUT93), .B2(G355), .ZN(new_n787));
  OR2_X1    g0587(.A1(G355), .A2(KEYINPUT93), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n787), .A2(new_n788), .B1(new_n456), .B2(new_n665), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n776), .A2(new_n780), .B1(new_n782), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n731), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n726), .B1(new_n724), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT99), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  AOI21_X1  g0595(.A(new_n649), .B1(new_n627), .B2(new_n630), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n656), .A2(new_n357), .ZN(new_n797));
  MUX2_X1   g0597(.A(new_n377), .B(new_n633), .S(new_n797), .Z(new_n798));
  XNOR2_X1  g0598(.A(new_n796), .B(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n717), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n724), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n778), .A2(new_n728), .A3(new_n779), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n724), .B1(new_n804), .B2(G77), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n428), .B1(new_n752), .B2(new_n749), .C1(new_n806), .C2(new_n734), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n762), .B(new_n807), .C1(G303), .C2(new_n757), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G87), .A2(new_n744), .B1(new_n745), .B2(G107), .ZN(new_n809));
  INV_X1    g0609(.A(new_n737), .ZN(new_n810));
  INV_X1    g0610(.A(G283), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n811), .B1(new_n748), .B2(new_n456), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT100), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G143), .A2(new_n735), .B1(new_n771), .B2(G159), .ZN(new_n815));
  INV_X1    g0615(.A(G150), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n810), .B2(new_n816), .C1(new_n817), .C2(new_n773), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT34), .Z(new_n819));
  NAND2_X1  g0619(.A1(new_n744), .A2(G68), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n745), .A2(G50), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n756), .A2(G58), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n428), .B1(new_n753), .B2(G132), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n814), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n805), .B1(new_n825), .B2(new_n780), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n798), .B2(new_n728), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT101), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n803), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G384));
  OAI21_X1  g0630(.A(G77), .B1(new_n380), .B2(new_n307), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n831), .A2(new_n217), .B1(G50), .B2(new_n307), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n832), .A2(G1), .A3(new_n642), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT102), .ZN(new_n834));
  INV_X1    g0634(.A(new_n585), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n456), .B(new_n216), .C1(new_n835), .C2(KEYINPUT35), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(KEYINPUT35), .B2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT36), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  INV_X1    g0640(.A(new_n341), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(new_n339), .A3(new_n338), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n322), .A3(new_n656), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n398), .B1(KEYINPUT16), .B2(new_n397), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n402), .ZN(new_n845));
  INV_X1    g0645(.A(new_n647), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n443), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n403), .A2(new_n415), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n403), .A2(new_n846), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n436), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n419), .A2(new_n647), .B1(new_n844), .B2(new_n402), .ZN(new_n854));
  INV_X1    g0654(.A(new_n436), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT38), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(KEYINPUT38), .B(new_n857), .C1(new_n451), .C2(new_n847), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT39), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n436), .B1(new_n418), .B2(new_n419), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n418), .A2(new_n647), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n853), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n438), .A2(new_n439), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n864), .B1(new_n421), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT39), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n859), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n861), .A2(new_n862), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n857), .B1(new_n451), .B2(new_n847), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n870), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n872), .B1(new_n876), .B2(new_n859), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n859), .A2(new_n871), .A3(new_n872), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT103), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n843), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n634), .A2(new_n649), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n796), .B2(new_n798), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n322), .B(new_n649), .C1(new_n842), .C2(new_n635), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n342), .B(new_n345), .C1(new_n321), .C2(new_n656), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n876), .A2(new_n859), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(new_n889), .B1(new_n421), .B2(new_n647), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n453), .B1(new_n689), .B2(new_n718), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n640), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n891), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n859), .A2(new_n871), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n886), .A2(new_n798), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n709), .B(new_n710), .C1(new_n612), .C2(new_n649), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT40), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n798), .A3(new_n886), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n876), .B2(new_n859), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n900), .B2(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n453), .A2(new_n897), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(G330), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n894), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n246), .B2(new_n721), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n894), .A2(new_n905), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n840), .B1(new_n907), .B2(new_n908), .ZN(G367));
  OAI21_X1  g0709(.A(new_n611), .B1(new_n682), .B2(new_n656), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT105), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n681), .A2(new_n656), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n663), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT44), .Z(new_n915));
  NOR2_X1   g0715(.A1(new_n913), .A2(new_n663), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT45), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n660), .A2(KEYINPUT107), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n662), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n658), .A2(new_n661), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(new_n654), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n719), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n915), .A2(new_n919), .A3(new_n917), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n929), .A2(new_n719), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n666), .B(KEYINPUT41), .Z(new_n931));
  OAI21_X1  g0731(.A(new_n722), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n922), .B1(new_n911), .B2(new_n912), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  INV_X1    g0734(.A(new_n539), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n604), .B1(new_n911), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n934), .B1(new_n649), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(KEYINPUT106), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n649), .B1(new_n569), .B2(new_n571), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n629), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n622), .B2(new_n942), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT104), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n949), .B1(new_n941), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n660), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n913), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n932), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n234), .A2(new_n784), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n782), .B1(new_n212), .B2(new_n349), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n744), .A2(G77), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n258), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT109), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n748), .A2(new_n202), .B1(new_n752), .B2(new_n817), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G159), .B2(new_n737), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n962), .B(new_n964), .C1(new_n380), .C2(new_n767), .ZN(new_n965));
  INV_X1    g0765(.A(G143), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n773), .A2(new_n966), .B1(new_n734), .B2(new_n816), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n755), .A2(new_n307), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT108), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n961), .B2(new_n960), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n745), .A2(G116), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT46), .Z(new_n973));
  OAI22_X1  g0773(.A1(new_n810), .A2(new_n806), .B1(new_n773), .B2(new_n749), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G107), .B2(new_n756), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n744), .A2(G97), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n258), .B1(new_n735), .B2(G303), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G283), .A2(new_n771), .B1(new_n753), .B2(G317), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n965), .A2(new_n971), .B1(new_n973), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT47), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n780), .B1(new_n980), .B2(new_n981), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n724), .B1(new_n957), .B2(new_n958), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT110), .Z(new_n985));
  OR2_X1    g0785(.A1(new_n944), .A2(new_n730), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n956), .A2(new_n987), .ZN(G387));
  OAI21_X1  g0788(.A(new_n258), .B1(new_n748), .B2(new_n307), .ZN(new_n989));
  INV_X1    g0789(.A(G159), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n990), .A2(new_n773), .B1(new_n810), .B2(new_n271), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n989), .B(new_n991), .C1(G150), .C2(new_n753), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n734), .A2(new_n202), .B1(new_n755), .B2(new_n349), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n745), .A2(G77), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n992), .A2(new_n976), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n767), .A2(new_n806), .B1(new_n811), .B2(new_n755), .ZN(new_n997));
  INV_X1    g0797(.A(G317), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n734), .A2(new_n998), .B1(new_n748), .B2(new_n466), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT113), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(KEYINPUT113), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n737), .A2(G311), .B1(new_n757), .B2(G322), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n997), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(KEYINPUT49), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n258), .B1(new_n753), .B2(G326), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n456), .C2(new_n760), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT49), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n996), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n780), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n231), .A2(new_n469), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n272), .A2(new_n202), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT50), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n668), .B(new_n469), .C1(new_n307), .C2(new_n205), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n784), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1013), .B1(KEYINPUT111), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT111), .B2(new_n1017), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(G107), .B2(new_n212), .C1(new_n668), .C2(new_n786), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n782), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1012), .A2(new_n1021), .A3(new_n724), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n659), .B2(new_n781), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n925), .B2(new_n723), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n926), .A2(new_n666), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n925), .A2(new_n719), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(G393));
  XNOR2_X1  g0827(.A(new_n918), .B(new_n953), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n929), .B(new_n666), .C1(new_n1028), .C2(new_n927), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n913), .A2(new_n781), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n782), .B1(new_n207), .B2(new_n212), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n241), .A2(new_n665), .A3(new_n258), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n724), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n755), .A2(new_n205), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n258), .B1(new_n752), .B2(new_n966), .C1(new_n271), .C2(new_n748), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G50), .C2(new_n737), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n773), .A2(new_n816), .B1(new_n734), .B2(new_n990), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT51), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G68), .A2(new_n745), .B1(new_n744), .B2(G87), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n761), .B1(G283), .B2(new_n745), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n428), .B1(new_n748), .B2(new_n806), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G322), .B2(new_n753), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n756), .A2(G116), .B1(G303), .B2(new_n737), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n773), .A2(new_n998), .B1(new_n734), .B2(new_n749), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT52), .Z(new_n1047));
  OAI21_X1  g0847(.A(new_n1040), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1033), .B1(new_n1048), .B2(new_n780), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1028), .A2(new_n723), .B1(new_n1030), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT114), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n1029), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n1029), .B2(new_n1050), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(G390));
  NAND3_X1  g0855(.A1(new_n874), .A2(new_n879), .A3(new_n727), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n724), .B1(new_n804), .B2(new_n272), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n773), .A2(new_n811), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1034), .B(new_n1058), .C1(G107), .C2(new_n737), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n748), .A2(new_n207), .B1(new_n752), .B2(new_n806), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n258), .B(new_n1060), .C1(G116), .C2(new_n735), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n769), .A2(new_n820), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n428), .B1(new_n753), .B2(G125), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n760), .B2(new_n202), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT116), .Z(new_n1065));
  INV_X1    g0865(.A(G128), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n773), .A2(new_n1066), .B1(new_n755), .B2(new_n990), .ZN(new_n1067));
  INV_X1    g0867(.A(G132), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n810), .A2(new_n817), .B1(new_n734), .B2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT54), .B(G143), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT115), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1067), .B(new_n1069), .C1(new_n771), .C2(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n745), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT53), .B1(new_n745), .B2(G150), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1062), .B1(new_n1065), .B2(new_n1075), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT117), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1077), .A2(new_n780), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(KEYINPUT117), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1057), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1056), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n843), .B1(new_n883), .B2(new_n887), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n874), .A2(new_n879), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n688), .A2(new_n656), .A3(new_n798), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n882), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n843), .B(new_n895), .C1(new_n1086), .C2(new_n887), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n897), .A2(new_n886), .A3(G330), .A4(new_n798), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1083), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1081), .B1(new_n1093), .B2(new_n722), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n453), .A2(new_n717), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n892), .A2(new_n640), .A3(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(G330), .B(new_n798), .C1(new_n711), .C2(new_n715), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n887), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1098), .A2(new_n1084), .A3(new_n1085), .A4(new_n1089), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1098), .A2(new_n1089), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n883), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1091), .A2(new_n1092), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n667), .B1(new_n1093), .B2(new_n1102), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1094), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G378));
  INV_X1    g0907(.A(KEYINPUT119), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n898), .B(G330), .C1(new_n900), .C2(KEYINPUT40), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n291), .A2(new_n846), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n306), .B(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n890), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1114), .A2(new_n1115), .B1(new_n880), .B2(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n881), .A2(new_n1118), .A3(new_n890), .A4(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1104), .A2(new_n1096), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1108), .B1(new_n1121), .B2(KEYINPUT57), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1117), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1083), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1089), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n1102), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n892), .A2(new_n640), .A3(new_n1095), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1123), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT57), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(KEYINPUT119), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1104), .A2(new_n1096), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT118), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1117), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1120), .A2(new_n1117), .A3(new_n1132), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1131), .A2(new_n1133), .A3(KEYINPUT57), .A4(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1122), .A2(new_n1130), .A3(new_n666), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1113), .A2(new_n727), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n724), .B1(new_n804), .B2(G50), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1139));
  INV_X1    g0939(.A(G41), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n428), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n773), .A2(new_n456), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n968), .B(new_n1142), .C1(G97), .C2(new_n737), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n744), .A2(G58), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n734), .A2(new_n208), .B1(new_n748), .B2(new_n349), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1140), .B(new_n428), .C1(new_n752), .C2(new_n811), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1143), .A2(new_n995), .A3(new_n1144), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT58), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1141), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n745), .A2(new_n1071), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n734), .A2(new_n1066), .B1(new_n748), .B2(new_n817), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G132), .B2(new_n737), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n756), .A2(G150), .B1(G125), .B2(new_n757), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n744), .A2(G159), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G33), .B(G41), .C1(new_n753), .C2(G124), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1150), .B1(new_n1149), .B2(new_n1148), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1138), .B1(new_n1161), .B2(new_n780), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1123), .A2(new_n723), .B1(new_n1137), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1136), .A2(new_n1163), .ZN(G375));
  NOR2_X1   g0964(.A1(new_n1103), .A2(new_n931), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT120), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n883), .B1(new_n1098), .B2(new_n1089), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1086), .B2(new_n1100), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1169), .B2(new_n722), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1101), .A2(KEYINPUT120), .A3(new_n723), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n724), .B1(new_n804), .B2(G68), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n773), .A2(new_n1068), .B1(new_n755), .B2(new_n202), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n734), .A2(new_n817), .B1(new_n748), .B2(new_n816), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n258), .B1(new_n752), .B2(new_n1066), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n745), .A2(G159), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1071), .A2(new_n737), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1176), .A2(new_n1144), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n745), .A2(G97), .B1(G303), .B2(new_n753), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT121), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n428), .B1(new_n734), .B2(new_n811), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G107), .B2(new_n771), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n757), .A2(G294), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n756), .A2(new_n350), .B1(G116), .B2(new_n737), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n959), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1179), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1172), .B1(new_n1187), .B2(new_n780), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n886), .B2(new_n728), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1170), .A2(new_n1171), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1166), .A2(new_n1191), .ZN(G381));
  OR3_X1    g0992(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(G387), .A2(G381), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(G375), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1194), .A2(new_n1195), .A3(new_n1054), .A4(new_n1106), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT122), .ZN(G407));
  NAND2_X1  g0997(.A1(new_n1106), .A2(new_n648), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G407), .B(G213), .C1(G375), .C2(new_n1198), .ZN(G409));
  INV_X1    g0999(.A(KEYINPUT60), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n667), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1169), .A2(new_n1127), .A3(KEYINPUT60), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT123), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT123), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1201), .A2(new_n1202), .A3(new_n1206), .A4(new_n1203), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G384), .B1(new_n1208), .B2(new_n1191), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n829), .B(new_n1190), .C1(new_n1205), .C2(new_n1207), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n648), .A2(G213), .ZN(new_n1212));
  INV_X1    g1012(.A(G2897), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(KEYINPUT124), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(KEYINPUT124), .B2(new_n1213), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n666), .B1(new_n1169), .B2(new_n1127), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT60), .B1(new_n1169), .B2(new_n1127), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1206), .B1(new_n1219), .B2(new_n1203), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1207), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1191), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n829), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1208), .A2(G384), .A3(new_n1191), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT125), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(KEYINPUT125), .B(new_n1226), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1216), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1136), .A2(G378), .A3(new_n1163), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1133), .A2(new_n723), .A3(new_n1134), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1137), .A2(new_n1162), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1128), .A2(new_n931), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1106), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1212), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT61), .B1(new_n1231), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT63), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1239), .B2(new_n1225), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1054), .A2(G387), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n956), .B(new_n987), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G393), .B(new_n794), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1212), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(KEYINPUT63), .A3(new_n1211), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1240), .A2(new_n1242), .A3(new_n1248), .A4(new_n1251), .ZN(new_n1252));
  XOR2_X1   g1052(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1253));
  AND3_X1   g1053(.A1(new_n1250), .A2(new_n1211), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT61), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1250), .B2(new_n1230), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1250), .B2(new_n1211), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1254), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1252), .B1(new_n1259), .B2(new_n1248), .ZN(G405));
  NAND2_X1  g1060(.A1(G375), .A2(new_n1106), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1232), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(KEYINPUT127), .A3(new_n1211), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1211), .A2(KEYINPUT127), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1261), .A2(new_n1232), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1248), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(G402));
endmodule


