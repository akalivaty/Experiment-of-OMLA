//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  INV_X1    g000(.A(KEYINPUT107), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT91), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n203), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  OAI221_X1 g007(.A(new_n207), .B1(KEYINPUT92), .B2(new_n208), .C1(new_n205), .C2(new_n204), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n208), .A2(KEYINPUT92), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT96), .ZN(new_n213));
  XOR2_X1   g012(.A(G57gat), .B(G64gat), .Z(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(KEYINPUT96), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G71gat), .B(G78gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT21), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(G183gat), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n222));
  NOR2_X1   g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n221), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n223), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n221), .B(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n225), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G127gat), .B(G155gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(G211gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(G231gat), .A2(G233gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n235), .B(new_n236), .Z(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n227), .A2(new_n230), .A3(new_n237), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G218gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT14), .ZN(new_n244));
  INV_X1    g043(.A(G29gat), .ZN(new_n245));
  INV_X1    g044(.A(G36gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(KEYINPUT87), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT87), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n250), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT88), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT89), .B(G36gat), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n252), .A2(new_n253), .B1(G29gat), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(new_n253), .B2(new_n252), .ZN(new_n256));
  INV_X1    g055(.A(G50gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT15), .B1(new_n257), .B2(G43gat), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(G43gat), .B2(new_n257), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n248), .B2(new_n247), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(G29gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n257), .A2(G43gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT90), .B(G43gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(new_n257), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n261), .B(new_n262), .C1(KEYINPUT15), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT17), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT101), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(G85gat), .A3(G92gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT100), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT100), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(G85gat), .A3(G92gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT7), .ZN(new_n275));
  NAND2_X1  g074(.A1(G99gat), .A2(G106gat), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n270), .A2(new_n275), .B1(KEYINPUT8), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT102), .B(G85gat), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT103), .B(G92gat), .Z(new_n279));
  OAI211_X1 g078(.A(new_n274), .B(new_n277), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(G99gat), .B(G106gat), .Z(new_n281));
  OR2_X1    g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n281), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT104), .A3(new_n283), .ZN(new_n284));
  OR3_X1    g083(.A1(new_n280), .A2(KEYINPUT104), .A3(new_n281), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  AND3_X1   g088(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n286), .B2(new_n267), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n289), .B1(new_n288), .B2(new_n291), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n243), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n288), .A2(new_n291), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G190gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(G218gat), .A3(new_n292), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(KEYINPUT105), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G134gat), .B(G162gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT105), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n293), .A2(new_n243), .A3(new_n294), .ZN(new_n306));
  AOI21_X1  g105(.A(G218gat), .B1(new_n297), .B2(new_n292), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n299), .A3(new_n303), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n242), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G230gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n218), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n284), .A2(new_n315), .A3(new_n285), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT10), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n282), .A2(new_n218), .A3(new_n283), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n286), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n314), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n314), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G176gat), .B(G204gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT106), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(G120gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G148gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n325), .B(new_n329), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n202), .B1(new_n311), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n242), .A2(new_n310), .A3(KEYINPUT107), .A4(new_n330), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n267), .ZN(new_n335));
  OR3_X1    g134(.A1(new_n211), .A2(new_n335), .A3(KEYINPUT93), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT93), .B1(new_n335), .B2(new_n211), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G229gat), .A2(G233gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n268), .A2(new_n211), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n338), .A2(KEYINPUT18), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n211), .ZN(new_n342));
  INV_X1    g141(.A(new_n337), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n335), .A2(new_n211), .A3(KEYINPUT93), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n339), .B(KEYINPUT13), .Z(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n336), .A2(new_n337), .B1(new_n268), .B2(new_n211), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT18), .B1(new_n349), .B2(new_n339), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT11), .B(G169gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(G197gat), .ZN(new_n353));
  XOR2_X1   g152(.A(G113gat), .B(G141gat), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT12), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n348), .B(new_n351), .C1(KEYINPUT94), .C2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n347), .A3(KEYINPUT94), .ZN(new_n358));
  INV_X1    g157(.A(new_n356), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n347), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n358), .B(new_n359), .C1(new_n360), .C2(new_n350), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n357), .A2(KEYINPUT95), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT95), .B1(new_n357), .B2(new_n361), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT31), .B(G50gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT3), .ZN(new_n367));
  XOR2_X1   g166(.A(G211gat), .B(G218gat), .Z(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT77), .ZN(new_n369));
  XNOR2_X1  g168(.A(G197gat), .B(G204gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT22), .ZN(new_n371));
  INV_X1    g170(.A(G211gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n243), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n369), .B(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n367), .B1(new_n375), .B2(KEYINPUT29), .ZN(new_n376));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT2), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT81), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G141gat), .B(G148gat), .Z(new_n381));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n382), .A3(KEYINPUT2), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n379), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n377), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n381), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n376), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n375), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n384), .A2(new_n389), .B1(new_n381), .B2(new_n392), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n367), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(G228gat), .B(G233gat), .C1(new_n395), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n374), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n404), .A2(new_n368), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n399), .B1(new_n404), .B2(new_n368), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT3), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n403), .B1(new_n407), .B2(new_n397), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n366), .B1(new_n402), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n412), .B(G22gat), .Z(new_n413));
  NAND3_X1  g212(.A1(new_n402), .A2(new_n366), .A3(new_n409), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n411), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT39), .ZN(new_n419));
  XOR2_X1   g218(.A(G113gat), .B(G120gat), .Z(new_n420));
  INV_X1    g219(.A(KEYINPUT1), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G127gat), .B(G134gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n426));
  NAND2_X1  g225(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n420), .A2(new_n423), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n428), .A2(KEYINPUT73), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(KEYINPUT73), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n394), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n428), .B(KEYINPUT73), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n397), .B1(new_n433), .B2(new_n425), .ZN(new_n434));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n394), .A2(KEYINPUT3), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n431), .A2(new_n440), .A3(new_n398), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n425), .A3(new_n397), .ZN(new_n442));
  INV_X1    g241(.A(new_n438), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  AOI211_X1 g244(.A(new_n419), .B(new_n437), .C1(new_n445), .C2(new_n436), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n419), .A3(new_n436), .ZN(new_n447));
  XOR2_X1   g246(.A(G1gat), .B(G29gat), .Z(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT85), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n447), .A2(new_n455), .A3(new_n452), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n446), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(KEYINPUT40), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n436), .B1(new_n432), .B2(new_n434), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n432), .B1(new_n441), .B2(KEYINPUT4), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT4), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n442), .B2(new_n435), .ZN(new_n462));
  OAI211_X1 g261(.A(KEYINPUT5), .B(new_n459), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n436), .A2(KEYINPUT5), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n439), .A2(new_n441), .A3(new_n444), .A4(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n452), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n457), .B2(KEYINPUT40), .ZN(new_n467));
  NAND2_X1  g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g269(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT27), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT27), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n474));
  AND4_X1   g273(.A1(new_n470), .A2(new_n472), .A3(new_n474), .A4(new_n289), .ZN(new_n475));
  AOI21_X1  g274(.A(G190gat), .B1(new_n471), .B2(KEYINPUT27), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n470), .B1(new_n476), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n469), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT70), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT70), .B(new_n469), .C1(new_n475), .C2(new_n477), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT27), .B(G183gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT71), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n483), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT28), .B(new_n289), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G183gat), .A2(G190gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(G169gat), .A2(G176gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n489), .B(KEYINPUT65), .Z(new_n490));
  INV_X1    g289(.A(G169gat), .ZN(new_n491));
  INV_X1    g290(.A(G176gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT26), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n493), .A2(KEYINPUT26), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n487), .A2(new_n488), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n498));
  MUX2_X1   g297(.A(KEYINPUT24), .B(new_n498), .S(new_n488), .Z(new_n499));
  INV_X1    g298(.A(KEYINPUT64), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n493), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(G169gat), .A2(G176gat), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT64), .B1(new_n503), .B2(KEYINPUT23), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(KEYINPUT23), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n499), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT66), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT25), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n499), .A2(new_n490), .A3(new_n505), .A4(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n507), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(new_n508), .A3(KEYINPUT25), .A4(new_n490), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n497), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n468), .B1(new_n515), .B2(KEYINPUT29), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n514), .ZN(new_n517));
  INV_X1    g316(.A(new_n468), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n396), .ZN(new_n521));
  XOR2_X1   g320(.A(G8gat), .B(G36gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G64gat), .ZN(new_n523));
  INV_X1    g322(.A(G92gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n399), .B1(new_n497), .B2(new_n514), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT79), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n526), .A2(new_n527), .A3(new_n518), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n517), .A2(new_n400), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n468), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT79), .B1(new_n517), .B2(new_n518), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n521), .B(new_n525), .C1(new_n532), .C2(new_n396), .ZN(new_n533));
  INV_X1    g332(.A(new_n525), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n519), .B(new_n527), .C1(new_n518), .C2(new_n526), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(KEYINPUT79), .A3(new_n468), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n396), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n375), .B1(new_n516), .B2(new_n519), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(new_n539), .A3(KEYINPUT30), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n541), .B(new_n534), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n458), .A2(new_n467), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT6), .ZN(new_n544));
  AOI211_X1 g343(.A(new_n544), .B(new_n452), .C1(new_n463), .C2(new_n465), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n441), .A2(KEYINPUT4), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n462), .B1(new_n546), .B2(new_n442), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n459), .A2(KEYINPUT5), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n452), .B(new_n465), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(new_n466), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n545), .B1(new_n551), .B2(new_n544), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n521), .B(new_n553), .C1(new_n532), .C2(new_n396), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT37), .B1(new_n537), .B2(new_n538), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n534), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT38), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n539), .B(new_n552), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n520), .A2(new_n375), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n559), .B(KEYINPUT37), .C1(new_n532), .C2(new_n375), .ZN(new_n560));
  AOI211_X1 g359(.A(KEYINPUT38), .B(new_n534), .C1(new_n560), .C2(new_n554), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n418), .B(new_n543), .C1(new_n558), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G227gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(new_n313), .ZN(new_n564));
  INV_X1    g363(.A(new_n431), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n497), .A2(new_n565), .A3(new_n514), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n565), .B1(new_n497), .B2(new_n514), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT34), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n566), .A2(new_n567), .ZN(new_n570));
  INV_X1    g369(.A(new_n564), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR4_X1   g371(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT34), .A4(new_n564), .ZN(new_n573));
  OAI211_X1 g372(.A(KEYINPUT32), .B(new_n568), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n497), .A2(new_n565), .A3(new_n514), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT34), .B1(new_n577), .B2(new_n564), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n568), .A2(KEYINPUT32), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n570), .A2(new_n569), .A3(new_n571), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT33), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n568), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT74), .B(G71gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G99gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G15gat), .B(G43gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n574), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n574), .B2(new_n581), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT75), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT76), .ZN(new_n592));
  INV_X1    g391(.A(new_n590), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n581), .A3(new_n588), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(KEYINPUT36), .B(new_n591), .C1(new_n595), .C2(KEYINPUT75), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n540), .A2(new_n542), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n551), .A2(KEYINPUT84), .A3(new_n544), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n463), .A2(new_n465), .ZN(new_n599));
  INV_X1    g398(.A(new_n452), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n544), .A3(new_n549), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT84), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n545), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n598), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n417), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT75), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n589), .A2(new_n590), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n592), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n562), .A2(new_n596), .A3(new_n608), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n593), .A2(new_n418), .A3(new_n594), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT35), .B1(new_n607), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT86), .ZN(new_n616));
  INV_X1    g415(.A(new_n552), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n597), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT35), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n589), .A2(new_n590), .A3(new_n417), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n552), .B1(new_n540), .B2(new_n542), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n621), .B1(new_n622), .B2(new_n616), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n615), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n364), .B1(new_n613), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n334), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(new_n606), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT108), .B(G1gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1324gat));
  INV_X1    g428(.A(new_n626), .ZN(new_n630));
  INV_X1    g429(.A(new_n597), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT16), .B(G8gat), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT109), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n634), .A2(KEYINPUT42), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(G8gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(KEYINPUT42), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(G1325gat));
  INV_X1    g437(.A(new_n596), .ZN(new_n639));
  INV_X1    g438(.A(new_n612), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n630), .A2(G15gat), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(G15gat), .B1(new_n630), .B2(new_n611), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(G1326gat));
  NOR2_X1   g444(.A1(new_n626), .A2(new_n418), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT43), .B(G22gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1327gat));
  AOI21_X1  g447(.A(new_n310), .B1(new_n613), .B2(new_n624), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n241), .A2(new_n330), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n364), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(G29gat), .A3(new_n606), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n624), .A2(KEYINPUT111), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT111), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n615), .B(new_n657), .C1(new_n620), .C2(new_n623), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n613), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n310), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n357), .A2(new_n361), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n665), .ZN(new_n666));
  AOI211_X1 g465(.A(new_n662), .B(new_n310), .C1(new_n613), .C2(new_n624), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n663), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT112), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n667), .B1(new_n661), .B2(new_n662), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT112), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n672), .A3(new_n666), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n606), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n655), .B1(new_n674), .B2(new_n245), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT113), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT113), .B(new_n655), .C1(new_n674), .C2(new_n245), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1328gat));
  AND3_X1   g478(.A1(new_n671), .A2(new_n672), .A3(new_n666), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n672), .B1(new_n671), .B2(new_n666), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n631), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT115), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n670), .A2(new_n673), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(KEYINPUT115), .A3(new_n631), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n254), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT114), .ZN(new_n689));
  NOR4_X1   g488(.A1(new_n652), .A2(new_n597), .A3(new_n254), .A4(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n652), .A2(new_n597), .A3(new_n254), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(KEYINPUT114), .B2(new_n688), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n690), .B1(new_n692), .B2(new_n689), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n687), .A2(new_n693), .ZN(G1329gat));
  OAI21_X1  g493(.A(new_n264), .B1(new_n669), .B2(new_n641), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n649), .A2(new_n651), .ZN(new_n696));
  INV_X1    g495(.A(new_n611), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n264), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(KEYINPUT47), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n699), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n642), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n264), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n703), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g503(.A(G50gat), .B1(new_n669), .B2(new_n418), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n652), .A2(KEYINPUT116), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n652), .A2(KEYINPUT116), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n706), .A2(new_n257), .A3(new_n417), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(KEYINPUT48), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n708), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n685), .A2(new_n417), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(G50gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n712), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g512(.A1(new_n659), .A2(new_n665), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n311), .A2(new_n330), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n606), .B(KEYINPUT117), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n597), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT49), .B(G64gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(G1333gat));
  NOR3_X1   g523(.A1(new_n716), .A2(G71gat), .A3(new_n697), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n714), .A2(new_n642), .A3(new_n715), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(G71gat), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g527(.A1(new_n716), .A2(new_n418), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g529(.A1(new_n242), .A2(new_n664), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n671), .A2(new_n331), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n278), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n732), .A2(new_n606), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n659), .A2(new_n660), .A3(new_n731), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT118), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n736), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n606), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n735), .A2(KEYINPUT118), .A3(new_n736), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n331), .A4(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n734), .B1(new_n743), .B2(new_n733), .ZN(G1336gat));
  INV_X1    g543(.A(new_n279), .ZN(new_n745));
  INV_X1    g544(.A(new_n732), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n631), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n597), .A2(G92gat), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g548(.A(new_n330), .B(new_n749), .C1(new_n737), .C2(new_n739), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT52), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n740), .A2(new_n331), .A3(new_n742), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n749), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n751), .B1(new_n747), .B2(new_n754), .ZN(G1337gat));
  OAI21_X1  g554(.A(G99gat), .B1(new_n732), .B2(new_n641), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n753), .A2(G99gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(new_n697), .ZN(G1338gat));
  INV_X1    g557(.A(G106gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n746), .B2(new_n417), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n418), .A2(G106gat), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g561(.A(new_n330), .B(new_n762), .C1(new_n737), .C2(new_n739), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT53), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n753), .B2(new_n762), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n760), .B2(new_n766), .ZN(G1339gat));
  OR2_X1    g566(.A1(new_n325), .A2(new_n329), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n319), .A2(new_n314), .A3(new_n320), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n322), .A2(KEYINPUT120), .A3(new_n769), .A4(KEYINPUT54), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n322), .A2(KEYINPUT54), .A3(new_n769), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n321), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n770), .B(new_n329), .C1(new_n771), .C2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n664), .A2(new_n768), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n348), .A2(new_n351), .A3(new_n356), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n349), .A2(new_n339), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n345), .A2(new_n346), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n355), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n331), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n779), .A2(new_n786), .B1(new_n304), .B2(new_n309), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n778), .A2(new_n768), .A3(new_n777), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n310), .A2(new_n788), .A3(new_n784), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT121), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n778), .A2(new_n768), .A3(new_n777), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(new_n304), .A3(new_n309), .A4(new_n785), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n784), .A2(new_n330), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n792), .B2(new_n664), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n791), .B(new_n793), .C1(new_n795), .C2(new_n660), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(new_n796), .A3(new_n241), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n242), .A2(new_n310), .A3(new_n665), .A4(new_n330), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT119), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n614), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n717), .A2(new_n631), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(G113gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(new_n664), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n631), .A2(new_n606), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n800), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT122), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n800), .A2(KEYINPUT122), .A3(new_n806), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n810), .A2(new_n364), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n805), .B1(new_n813), .B2(new_n804), .ZN(G1340gat));
  INV_X1    g613(.A(G120gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n803), .A2(new_n815), .A3(new_n331), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n810), .A2(new_n330), .A3(new_n812), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n815), .ZN(G1341gat));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n809), .A2(G127gat), .A3(new_n242), .A4(new_n811), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n802), .A2(new_n241), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(G127gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n819), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n820), .B(KEYINPUT123), .C1(G127gat), .C2(new_n822), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1342gat));
  NOR3_X1   g625(.A1(new_n802), .A2(G134gat), .A3(new_n310), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT56), .ZN(new_n828));
  INV_X1    g627(.A(G134gat), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n810), .A2(new_n310), .A3(new_n812), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n641), .A2(new_n806), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n792), .B1(new_n362), .B2(new_n363), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n660), .B1(new_n833), .B2(new_n786), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n241), .B1(new_n834), .B2(new_n789), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n799), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n417), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n832), .B1(new_n837), .B2(KEYINPUT57), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n418), .B1(new_n797), .B2(new_n799), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G141gat), .B1(new_n842), .B2(new_n364), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n418), .B(new_n642), .C1(new_n797), .C2(new_n799), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n801), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n364), .A2(G141gat), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT58), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n838), .A2(new_n664), .A3(new_n841), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n851), .A2(G141gat), .B1(new_n846), .B2(new_n847), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(G1344gat));
  OR3_X1    g652(.A1(new_n845), .A2(G148gat), .A3(new_n330), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n797), .A2(new_n799), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n417), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n332), .A2(new_n364), .A3(new_n333), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n835), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n857), .A2(KEYINPUT57), .B1(new_n417), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n832), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT124), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(KEYINPUT124), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n860), .A2(new_n331), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n855), .B1(new_n864), .B2(G148gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n838), .A2(new_n331), .A3(new_n841), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n866), .A2(new_n855), .A3(G148gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n854), .B1(new_n865), .B2(new_n867), .ZN(G1345gat));
  INV_X1    g667(.A(G155gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n845), .B2(new_n241), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n838), .A2(G155gat), .A3(new_n242), .A4(new_n841), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT125), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1346gat));
  INV_X1    g675(.A(G162gat), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n842), .A2(new_n877), .A3(new_n310), .ZN(new_n878));
  AOI21_X1  g677(.A(G162gat), .B1(new_n846), .B2(new_n660), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(G1347gat));
  AOI211_X1 g679(.A(new_n597), .B(new_n614), .C1(new_n797), .C2(new_n799), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(new_n606), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n491), .A3(new_n664), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n717), .A2(new_n631), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n800), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G169gat), .B1(new_n886), .B2(new_n364), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(G1348gat));
  NOR3_X1   g687(.A1(new_n886), .A2(new_n492), .A3(new_n330), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n882), .A2(new_n331), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n492), .ZN(G1349gat));
  NOR2_X1   g690(.A1(new_n484), .A2(new_n485), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n241), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n800), .A2(new_n606), .A3(new_n631), .A4(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n881), .A2(KEYINPUT126), .A3(new_n606), .A4(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G183gat), .B1(new_n886), .B2(new_n241), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT60), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n882), .A2(new_n289), .A3(new_n660), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n800), .A2(new_n660), .A3(new_n885), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n906), .A2(new_n907), .A3(G190gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(G190gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1351gat));
  NAND2_X1  g709(.A1(new_n859), .A2(new_n417), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n642), .A2(new_n884), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n911), .B(new_n912), .C1(new_n840), .C2(new_n839), .ZN(new_n913));
  OAI21_X1  g712(.A(G197gat), .B1(new_n913), .B2(new_n364), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n741), .A2(new_n597), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n844), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n916), .A2(G197gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n917), .B2(new_n665), .ZN(G1352gat));
  NOR3_X1   g717(.A1(new_n916), .A2(G204gat), .A3(new_n330), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n860), .A2(new_n331), .A3(new_n912), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G204gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n920), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(G1353gat));
  NAND4_X1  g724(.A1(new_n844), .A2(new_n372), .A3(new_n242), .A4(new_n915), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n860), .A2(new_n242), .A3(new_n912), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n928));
  OAI211_X1 g727(.A(KEYINPUT63), .B(G211gat), .C1(new_n913), .C2(new_n241), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n928), .B2(new_n930), .ZN(G1354gat));
  OAI21_X1  g730(.A(G218gat), .B1(new_n913), .B2(new_n310), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n844), .A2(new_n243), .A3(new_n915), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n310), .B2(new_n933), .ZN(G1355gat));
endmodule


