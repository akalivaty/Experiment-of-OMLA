

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594;

  NOR2_X1 U326 ( .A1(n554), .A2(n553), .ZN(n563) );
  XNOR2_X1 U327 ( .A(n344), .B(n343), .ZN(n356) );
  XNOR2_X1 U328 ( .A(n353), .B(n352), .ZN(n528) );
  XNOR2_X1 U329 ( .A(n335), .B(n334), .ZN(n550) );
  XNOR2_X1 U330 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U331 ( .A(n479), .B(KEYINPUT120), .ZN(n480) );
  INV_X1 U332 ( .A(KEYINPUT99), .ZN(n345) );
  XNOR2_X1 U333 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U334 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U335 ( .A(n348), .B(n347), .ZN(n351) );
  XOR2_X1 U336 ( .A(n571), .B(KEYINPUT36), .Z(n591) );
  XNOR2_X1 U337 ( .A(n486), .B(KEYINPUT121), .ZN(n572) );
  INV_X1 U338 ( .A(G106GAT), .ZN(n457) );
  XNOR2_X1 U339 ( .A(n314), .B(n313), .ZN(n532) );
  XNOR2_X1 U340 ( .A(n488), .B(KEYINPUT122), .ZN(n489) );
  XNOR2_X1 U341 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U342 ( .A(n490), .B(n489), .ZN(G1350GAT) );
  XNOR2_X1 U343 ( .A(KEYINPUT86), .B(KEYINPUT19), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n294), .B(KEYINPUT17), .ZN(n295) );
  XOR2_X1 U345 ( .A(n295), .B(KEYINPUT85), .Z(n297) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n339) );
  XOR2_X1 U348 ( .A(G134GAT), .B(G190GAT), .Z(n299) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G99GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U351 ( .A(KEYINPUT84), .B(KEYINPUT87), .Z(n301) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(G71GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U354 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U355 ( .A(G183GAT), .B(G176GAT), .Z(n305) );
  NAND2_X1 U356 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U358 ( .A(KEYINPUT20), .B(n306), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n339), .B(n309), .ZN(n314) );
  XOR2_X1 U361 ( .A(KEYINPUT0), .B(G127GAT), .Z(n311) );
  XNOR2_X1 U362 ( .A(KEYINPUT83), .B(G120GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U364 ( .A(G113GAT), .B(n312), .Z(n333) );
  INV_X1 U365 ( .A(n333), .ZN(n313) );
  XOR2_X1 U366 ( .A(G85GAT), .B(G155GAT), .Z(n316) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(G162GAT), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U369 ( .A(KEYINPUT95), .B(KEYINPUT1), .Z(n318) );
  XNOR2_X1 U370 ( .A(G148GAT), .B(KEYINPUT6), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U372 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U373 ( .A(G134GAT), .B(KEYINPUT79), .Z(n415) );
  XOR2_X1 U374 ( .A(KEYINPUT4), .B(KEYINPUT97), .Z(n322) );
  NAND2_X1 U375 ( .A1(G225GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n415), .B(n323), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U379 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n327) );
  XNOR2_X1 U380 ( .A(G1GAT), .B(G57GAT), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U382 ( .A(n329), .B(n328), .Z(n335) );
  XOR2_X1 U383 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n331) );
  XNOR2_X1 U384 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U386 ( .A(G141GAT), .B(n332), .Z(n371) );
  XNOR2_X1 U387 ( .A(n333), .B(n371), .ZN(n334) );
  XOR2_X1 U388 ( .A(G64GAT), .B(KEYINPUT75), .Z(n337) );
  XNOR2_X1 U389 ( .A(G204GAT), .B(G92GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(G176GAT), .B(n338), .Z(n446) );
  XNOR2_X1 U392 ( .A(n339), .B(n446), .ZN(n353) );
  XOR2_X1 U393 ( .A(G36GAT), .B(G190GAT), .Z(n401) );
  XNOR2_X1 U394 ( .A(KEYINPUT91), .B(KEYINPUT89), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n340), .B(KEYINPUT21), .ZN(n344) );
  XNOR2_X1 U396 ( .A(G197GAT), .B(G218GAT), .ZN(n342) );
  INV_X1 U397 ( .A(KEYINPUT90), .ZN(n341) );
  XOR2_X1 U398 ( .A(n401), .B(n356), .Z(n348) );
  NAND2_X1 U399 ( .A1(G226GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U400 ( .A(G8GAT), .B(G183GAT), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n349), .B(G211GAT), .ZN(n386) );
  XNOR2_X1 U402 ( .A(n386), .B(KEYINPUT98), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n352) );
  INV_X1 U404 ( .A(KEYINPUT100), .ZN(n354) );
  XNOR2_X1 U405 ( .A(n528), .B(n354), .ZN(n355) );
  XNOR2_X1 U406 ( .A(KEYINPUT27), .B(n355), .ZN(n375) );
  XOR2_X1 U407 ( .A(KEYINPUT22), .B(G211GAT), .Z(n358) );
  XNOR2_X1 U408 ( .A(KEYINPUT24), .B(n356), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U410 ( .A(n359), .B(KEYINPUT88), .Z(n369) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(KEYINPUT78), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n360), .B(G162GAT), .ZN(n406) );
  XOR2_X1 U413 ( .A(n406), .B(KEYINPUT23), .Z(n362) );
  NAND2_X1 U414 ( .A1(G228GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n367) );
  XNOR2_X1 U416 ( .A(G106GAT), .B(G78GAT), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n363), .B(G148GAT), .ZN(n451) );
  XOR2_X1 U418 ( .A(G22GAT), .B(G155GAT), .Z(n385) );
  XOR2_X1 U419 ( .A(n451), .B(n385), .Z(n365) );
  XNOR2_X1 U420 ( .A(G204GAT), .B(KEYINPUT94), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n483) );
  XOR2_X1 U425 ( .A(KEYINPUT28), .B(n483), .Z(n522) );
  NOR2_X1 U426 ( .A1(n375), .A2(n522), .ZN(n372) );
  NAND2_X1 U427 ( .A1(n550), .A2(n372), .ZN(n534) );
  NOR2_X1 U428 ( .A1(n532), .A2(n534), .ZN(n382) );
  NOR2_X1 U429 ( .A1(n532), .A2(n483), .ZN(n374) );
  XNOR2_X1 U430 ( .A(KEYINPUT101), .B(KEYINPUT26), .ZN(n373) );
  XOR2_X1 U431 ( .A(n374), .B(n373), .Z(n577) );
  INV_X1 U432 ( .A(n577), .ZN(n376) );
  NOR2_X1 U433 ( .A1(n376), .A2(n375), .ZN(n552) );
  NAND2_X1 U434 ( .A1(n528), .A2(n532), .ZN(n377) );
  NAND2_X1 U435 ( .A1(n483), .A2(n377), .ZN(n378) );
  XNOR2_X1 U436 ( .A(KEYINPUT25), .B(n378), .ZN(n379) );
  NOR2_X1 U437 ( .A1(n552), .A2(n379), .ZN(n380) );
  NOR2_X1 U438 ( .A1(n550), .A2(n380), .ZN(n381) );
  NOR2_X1 U439 ( .A1(n382), .A2(n381), .ZN(n495) );
  XOR2_X1 U440 ( .A(KEYINPUT15), .B(G64GAT), .Z(n384) );
  XNOR2_X1 U441 ( .A(G127GAT), .B(G78GAT), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n399) );
  XOR2_X1 U443 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U446 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n390) );
  XNOR2_X1 U447 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U449 ( .A(n392), .B(n391), .Z(n397) );
  XNOR2_X1 U450 ( .A(G15GAT), .B(G1GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n393), .B(KEYINPUT69), .ZN(n429) );
  XOR2_X1 U452 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n395) );
  XNOR2_X1 U453 ( .A(G71GAT), .B(G57GAT), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n450) );
  XNOR2_X1 U455 ( .A(n429), .B(n450), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U457 ( .A(n399), .B(n398), .Z(n492) );
  INV_X1 U458 ( .A(n492), .ZN(n588) );
  NOR2_X1 U459 ( .A1(n495), .A2(n588), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n400), .B(KEYINPUT103), .ZN(n419) );
  XOR2_X1 U461 ( .A(G99GAT), .B(G85GAT), .Z(n442) );
  XOR2_X1 U462 ( .A(n442), .B(n401), .Z(n403) );
  NAND2_X1 U463 ( .A1(G232GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n411) );
  XOR2_X1 U465 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n409) );
  XOR2_X1 U466 ( .A(KEYINPUT9), .B(G92GAT), .Z(n405) );
  XNOR2_X1 U467 ( .A(G106GAT), .B(G218GAT), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U471 ( .A(n411), .B(n410), .Z(n418) );
  XOR2_X1 U472 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n413) );
  XNOR2_X1 U473 ( .A(G43GAT), .B(G29GAT), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U475 ( .A(KEYINPUT7), .B(n414), .ZN(n437) );
  INV_X1 U476 ( .A(n437), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X2 U478 ( .A(n418), .B(n417), .ZN(n571) );
  NOR2_X1 U479 ( .A1(n419), .A2(n591), .ZN(n420) );
  XNOR2_X1 U480 ( .A(KEYINPUT37), .B(n420), .ZN(n506) );
  XOR2_X1 U481 ( .A(KEYINPUT66), .B(G8GAT), .Z(n422) );
  XNOR2_X1 U482 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n436) );
  XOR2_X1 U484 ( .A(G141GAT), .B(G197GAT), .Z(n424) );
  XNOR2_X1 U485 ( .A(G169GAT), .B(G22GAT), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U487 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n426) );
  XNOR2_X1 U488 ( .A(G113GAT), .B(KEYINPUT65), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n434) );
  XOR2_X1 U491 ( .A(G36GAT), .B(n429), .Z(n431) );
  NAND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U494 ( .A(G50GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U497 ( .A(n438), .B(n437), .Z(n465) );
  XOR2_X1 U498 ( .A(KEYINPUT73), .B(KEYINPUT76), .Z(n440) );
  XNOR2_X1 U499 ( .A(KEYINPUT32), .B(KEYINPUT74), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U501 ( .A(n441), .B(KEYINPUT77), .Z(n444) );
  XNOR2_X1 U502 ( .A(G120GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n455) );
  XOR2_X1 U505 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n448) );
  NAND2_X1 U506 ( .A1(G230GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U508 ( .A(n449), .B(KEYINPUT31), .Z(n453) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n455), .B(n454), .ZN(n582) );
  INV_X1 U512 ( .A(n582), .ZN(n491) );
  XNOR2_X1 U513 ( .A(KEYINPUT41), .B(n491), .ZN(n567) );
  NAND2_X1 U514 ( .A1(n465), .A2(n567), .ZN(n517) );
  NOR2_X1 U515 ( .A1(n506), .A2(n517), .ZN(n456) );
  XOR2_X1 U516 ( .A(KEYINPUT105), .B(n456), .Z(n530) );
  AND2_X1 U517 ( .A1(n530), .A2(n522), .ZN(n460) );
  XNOR2_X1 U518 ( .A(KEYINPUT106), .B(KEYINPUT44), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n460), .B(n459), .ZN(G1339GAT) );
  INV_X1 U520 ( .A(KEYINPUT45), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n492), .A2(n591), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n463), .A2(n582), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n464), .B(KEYINPUT109), .ZN(n466) );
  INV_X1 U525 ( .A(n465), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n466), .A2(n469), .ZN(n468) );
  INV_X1 U527 ( .A(KEYINPUT110), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n468), .B(n467), .ZN(n476) );
  NAND2_X1 U529 ( .A1(n567), .A2(n469), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT108), .B(KEYINPUT46), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U532 ( .A(KEYINPUT107), .B(n588), .ZN(n544) );
  NAND2_X1 U533 ( .A1(n472), .A2(n544), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n473), .A2(n571), .ZN(n474) );
  XNOR2_X1 U535 ( .A(KEYINPUT47), .B(n474), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n551) );
  AND2_X1 U539 ( .A1(n528), .A2(n551), .ZN(n481) );
  INV_X1 U540 ( .A(KEYINPUT54), .ZN(n479) );
  NOR2_X1 U541 ( .A1(n550), .A2(n482), .ZN(n576) );
  NAND2_X1 U542 ( .A1(n576), .A2(n483), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(KEYINPUT55), .ZN(n485) );
  NAND2_X1 U544 ( .A1(n485), .A2(n532), .ZN(n486) );
  INV_X1 U545 ( .A(n572), .ZN(n487) );
  NOR2_X1 U546 ( .A1(n487), .A2(n544), .ZN(n490) );
  INV_X1 U547 ( .A(G183GAT), .ZN(n488) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n499) );
  NAND2_X1 U549 ( .A1(n469), .A2(n491), .ZN(n507) );
  XNOR2_X1 U550 ( .A(KEYINPUT82), .B(KEYINPUT16), .ZN(n494) );
  NOR2_X1 U551 ( .A1(n571), .A2(n492), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(n497) );
  INV_X1 U553 ( .A(n495), .ZN(n496) );
  NAND2_X1 U554 ( .A1(n497), .A2(n496), .ZN(n516) );
  NOR2_X1 U555 ( .A1(n507), .A2(n516), .ZN(n503) );
  NAND2_X1 U556 ( .A1(n550), .A2(n503), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(G1324GAT) );
  NAND2_X1 U558 ( .A1(n503), .A2(n528), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U561 ( .A1(n503), .A2(n532), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  NAND2_X1 U563 ( .A1(n522), .A2(n503), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n504), .B(KEYINPUT102), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G22GAT), .B(n505), .ZN(G1327GAT) );
  XOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT39), .Z(n510) );
  NOR2_X1 U567 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n508), .B(KEYINPUT38), .ZN(n514) );
  NAND2_X1 U569 ( .A1(n550), .A2(n514), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  NAND2_X1 U571 ( .A1(n514), .A2(n528), .ZN(n511) );
  XNOR2_X1 U572 ( .A(n511), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U573 ( .A1(n514), .A2(n532), .ZN(n512) );
  XNOR2_X1 U574 ( .A(n512), .B(KEYINPUT40), .ZN(n513) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(n513), .ZN(G1330GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n522), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n515), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n519) );
  NOR2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n550), .A2(n523), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n519), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U582 ( .A1(n523), .A2(n528), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n532), .A2(n523), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(n526), .ZN(G1335GAT) );
  NAND2_X1 U590 ( .A1(n530), .A2(n550), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n530), .A2(n528), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n532), .A2(n530), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n536) );
  NAND2_X1 U597 ( .A1(n532), .A2(n551), .ZN(n533) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n547) );
  NAND2_X1 U599 ( .A1(n547), .A2(n469), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U603 ( .A1(n547), .A2(n567), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U605 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n542) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n546) );
  INV_X1 U609 ( .A(n547), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(n546), .B(n545), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U613 ( .A1(n547), .A2(n571), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n556) );
  INV_X1 U616 ( .A(n550), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n563), .A2(n469), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n556), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n558) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(n559), .Z(n561) );
  NAND2_X1 U624 ( .A1(n563), .A2(n567), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n588), .A2(n563), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U628 ( .A(G162GAT), .B(KEYINPUT119), .Z(n565) );
  NAND2_X1 U629 ( .A1(n571), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n469), .A2(n572), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n569) );
  NAND2_X1 U634 ( .A1(n572), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(n570), .ZN(G1349GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G190GAT), .B(n575), .ZN(G1351GAT) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n581) );
  XOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT124), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n590) );
  INV_X1 U644 ( .A(n590), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n587), .A2(n469), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n584) );
  NAND2_X1 U649 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n586) );
  XOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT125), .Z(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

