

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726;

  NOR2_X2 U365 ( .A1(n685), .A2(n552), .ZN(n540) );
  XNOR2_X2 U366 ( .A(n541), .B(KEYINPUT104), .ZN(n722) );
  NOR2_X2 U367 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U368 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X2 U369 ( .A1(n671), .A2(n669), .ZN(n531) );
  INV_X1 U370 ( .A(n536), .ZN(n654) );
  XNOR2_X2 U371 ( .A(G119), .B(G116), .ZN(n357) );
  AND2_X1 U372 ( .A1(n576), .A2(n575), .ZN(n577) );
  AND2_X1 U373 ( .A1(n599), .A2(n596), .ZN(n484) );
  XNOR2_X1 U374 ( .A(n496), .B(n495), .ZN(n644) );
  XNOR2_X1 U375 ( .A(n344), .B(KEYINPUT38), .ZN(n530) );
  XNOR2_X1 U376 ( .A(n354), .B(n400), .ZN(n538) );
  NAND2_X1 U377 ( .A1(n370), .A2(n580), .ZN(n373) );
  BUF_X1 U378 ( .A(n598), .Z(n343) );
  XNOR2_X1 U379 ( .A(n373), .B(n372), .ZN(n344) );
  BUF_X1 U380 ( .A(n427), .Z(n345) );
  XNOR2_X1 U381 ( .A(n582), .B(KEYINPUT65), .ZN(n346) );
  XNOR2_X1 U382 ( .A(n582), .B(KEYINPUT65), .ZN(n347) );
  XNOR2_X1 U383 ( .A(n472), .B(n471), .ZN(n598) );
  XNOR2_X1 U384 ( .A(n582), .B(KEYINPUT65), .ZN(n617) );
  NAND2_X2 U385 ( .A1(n649), .A2(n581), .ZN(n582) );
  XNOR2_X2 U386 ( .A(n376), .B(KEYINPUT83), .ZN(n546) );
  OR2_X1 U387 ( .A1(n483), .A2(n545), .ZN(n508) );
  OR2_X1 U388 ( .A1(n612), .A2(G902), .ZN(n354) );
  XNOR2_X1 U389 ( .A(n456), .B(n396), .ZN(n428) );
  XNOR2_X1 U390 ( .A(n658), .B(n479), .ZN(n549) );
  XNOR2_X1 U391 ( .A(n476), .B(n353), .ZN(n483) );
  XOR2_X1 U392 ( .A(KEYINPUT99), .B(n502), .Z(n670) );
  NOR2_X1 U393 ( .A1(G237), .A2(G953), .ZN(n422) );
  XNOR2_X1 U394 ( .A(n395), .B(n394), .ZN(n456) );
  XNOR2_X1 U395 ( .A(n538), .B(KEYINPUT1), .ZN(n478) );
  XNOR2_X1 U396 ( .A(KEYINPUT15), .B(G902), .ZN(n580) );
  INV_X1 U397 ( .A(n714), .ZN(n576) );
  NOR2_X1 U398 ( .A1(n572), .A2(KEYINPUT77), .ZN(n573) );
  OR2_X2 U399 ( .A1(n483), .A2(n355), .ZN(n489) );
  NAND2_X1 U400 ( .A1(n549), .A2(n352), .ZN(n355) );
  XNOR2_X1 U401 ( .A(n414), .B(n413), .ZN(n583) );
  XNOR2_X1 U402 ( .A(n713), .B(n398), .ZN(n612) );
  XNOR2_X1 U403 ( .A(n621), .B(n620), .ZN(n622) );
  NAND2_X1 U404 ( .A1(n585), .A2(G953), .ZN(n624) );
  NAND2_X1 U405 ( .A1(n470), .A2(n469), .ZN(n472) );
  AND2_X1 U406 ( .A1(n598), .A2(n596), .ZN(n348) );
  NOR2_X1 U407 ( .A1(n501), .A2(n500), .ZN(n349) );
  XOR2_X1 U408 ( .A(KEYINPUT16), .B(G122), .Z(n350) );
  XNOR2_X1 U409 ( .A(n546), .B(n377), .ZN(n551) );
  XOR2_X1 U410 ( .A(n489), .B(n488), .Z(n351) );
  AND2_X1 U411 ( .A1(n477), .A2(n651), .ZN(n352) );
  XOR2_X1 U412 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n353) );
  XNOR2_X2 U413 ( .A(G143), .B(G128), .ZN(n395) );
  XNOR2_X1 U414 ( .A(n360), .B(G104), .ZN(n387) );
  XNOR2_X1 U415 ( .A(n387), .B(n350), .ZN(n361) );
  XNOR2_X2 U416 ( .A(n519), .B(n518), .ZN(n702) );
  INV_X1 U417 ( .A(KEYINPUT34), .ZN(n436) );
  XNOR2_X1 U418 ( .A(n437), .B(n436), .ZN(n470) );
  BUF_X1 U419 ( .A(n478), .Z(n658) );
  INV_X1 U420 ( .A(KEYINPUT120), .ZN(n587) );
  XNOR2_X2 U421 ( .A(G113), .B(KEYINPUT70), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n359) );
  XNOR2_X1 U423 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n427) );
  XNOR2_X2 U425 ( .A(G110), .B(G107), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n427), .B(n361), .ZN(n693) );
  XNOR2_X1 U427 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n363) );
  INV_X4 U428 ( .A(G953), .ZN(n703) );
  NAND2_X1 U429 ( .A1(n703), .A2(G224), .ZN(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n366) );
  XNOR2_X2 U431 ( .A(KEYINPUT66), .B(G101), .ZN(n392) );
  XNOR2_X1 U432 ( .A(KEYINPUT86), .B(KEYINPUT4), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n392), .B(n364), .ZN(n365) );
  XNOR2_X1 U434 ( .A(n366), .B(n365), .ZN(n368) );
  XNOR2_X1 U435 ( .A(G146), .B(G125), .ZN(n409) );
  XNOR2_X1 U436 ( .A(n395), .B(n409), .ZN(n367) );
  XNOR2_X1 U437 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n693), .B(n369), .ZN(n618) );
  INV_X1 U439 ( .A(n618), .ZN(n370) );
  INV_X1 U440 ( .A(G902), .ZN(n466) );
  INV_X1 U441 ( .A(G237), .ZN(n371) );
  NAND2_X1 U442 ( .A1(n466), .A2(n371), .ZN(n374) );
  NAND2_X1 U443 ( .A1(n374), .A2(G210), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n373), .B(n372), .ZN(n524) );
  NAND2_X1 U445 ( .A1(n374), .A2(G214), .ZN(n667) );
  INV_X1 U446 ( .A(n667), .ZN(n375) );
  OR2_X2 U447 ( .A1(n524), .A2(n375), .ZN(n376) );
  XNOR2_X1 U448 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n377) );
  NAND2_X1 U449 ( .A1(G237), .A2(G234), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n378), .B(KEYINPUT14), .ZN(n650) );
  NOR2_X1 U451 ( .A1(G902), .A2(n703), .ZN(n380) );
  NOR2_X1 U452 ( .A1(G953), .A2(G952), .ZN(n379) );
  NOR2_X1 U453 ( .A1(n380), .A2(n379), .ZN(n381) );
  NAND2_X1 U454 ( .A1(n650), .A2(n381), .ZN(n520) );
  AND2_X1 U455 ( .A1(G953), .A2(G898), .ZN(n382) );
  OR2_X1 U456 ( .A1(n520), .A2(n382), .ZN(n383) );
  OR2_X2 U457 ( .A1(n551), .A2(n383), .ZN(n386) );
  INV_X1 U458 ( .A(KEYINPUT84), .ZN(n384) );
  XNOR2_X1 U459 ( .A(n384), .B(KEYINPUT0), .ZN(n385) );
  XNOR2_X2 U460 ( .A(n386), .B(n385), .ZN(n492) );
  BUF_X1 U461 ( .A(n387), .Z(n391) );
  XNOR2_X1 U462 ( .A(KEYINPUT87), .B(G140), .ZN(n389) );
  NAND2_X1 U463 ( .A1(n703), .A2(G227), .ZN(n388) );
  XNOR2_X1 U464 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U465 ( .A(n391), .B(n390), .ZN(n393) );
  XNOR2_X1 U466 ( .A(n392), .B(G146), .ZN(n426) );
  XNOR2_X1 U467 ( .A(n393), .B(n426), .ZN(n398) );
  INV_X1 U468 ( .A(G134), .ZN(n394) );
  XNOR2_X1 U469 ( .A(KEYINPUT4), .B(G131), .ZN(n396) );
  INV_X1 U470 ( .A(KEYINPUT68), .ZN(n397) );
  XNOR2_X1 U471 ( .A(n397), .B(G137), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n428), .B(n401), .ZN(n713) );
  INV_X1 U473 ( .A(KEYINPUT69), .ZN(n399) );
  XNOR2_X1 U474 ( .A(n399), .B(G469), .ZN(n400) );
  XNOR2_X1 U475 ( .A(G119), .B(G110), .ZN(n402) );
  XNOR2_X1 U476 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U477 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n404) );
  XNOR2_X1 U478 ( .A(G128), .B(KEYINPUT79), .ZN(n403) );
  XNOR2_X1 U479 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U480 ( .A(n406), .B(n405), .Z(n414) );
  INV_X1 U481 ( .A(KEYINPUT10), .ZN(n407) );
  XNOR2_X1 U482 ( .A(n407), .B(G140), .ZN(n408) );
  XNOR2_X1 U483 ( .A(n409), .B(n408), .ZN(n711) );
  XOR2_X1 U484 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n411) );
  NAND2_X1 U485 ( .A1(G234), .A2(n703), .ZN(n410) );
  XNOR2_X1 U486 ( .A(n411), .B(n410), .ZN(n459) );
  NAND2_X1 U487 ( .A1(n459), .A2(G221), .ZN(n412) );
  XNOR2_X1 U488 ( .A(n711), .B(n412), .ZN(n413) );
  NAND2_X1 U489 ( .A1(n583), .A2(n466), .ZN(n418) );
  NAND2_X1 U490 ( .A1(G234), .A2(n580), .ZN(n415) );
  XNOR2_X1 U491 ( .A(KEYINPUT20), .B(n415), .ZN(n419) );
  AND2_X1 U492 ( .A1(n419), .A2(G217), .ZN(n416) );
  XNOR2_X1 U493 ( .A(KEYINPUT25), .B(n416), .ZN(n417) );
  XNOR2_X1 U494 ( .A(n418), .B(n417), .ZN(n533) );
  AND2_X1 U495 ( .A1(n419), .A2(G221), .ZN(n421) );
  INV_X1 U496 ( .A(KEYINPUT21), .ZN(n420) );
  XNOR2_X1 U497 ( .A(n421), .B(n420), .ZN(n652) );
  INV_X1 U498 ( .A(n652), .ZN(n534) );
  AND2_X1 U499 ( .A1(n533), .A2(n534), .ZN(n657) );
  AND2_X1 U500 ( .A1(n478), .A2(n657), .ZN(n494) );
  XNOR2_X1 U501 ( .A(KEYINPUT76), .B(n422), .ZN(n443) );
  NAND2_X1 U502 ( .A1(n443), .A2(G210), .ZN(n424) );
  XNOR2_X1 U503 ( .A(G137), .B(KEYINPUT5), .ZN(n423) );
  XNOR2_X1 U504 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U505 ( .A(n426), .B(n425), .ZN(n430) );
  XNOR2_X1 U506 ( .A(n345), .B(n428), .ZN(n429) );
  XNOR2_X1 U507 ( .A(n430), .B(n429), .ZN(n601) );
  NOR2_X1 U508 ( .A1(n601), .A2(G902), .ZN(n433) );
  XNOR2_X1 U509 ( .A(KEYINPUT89), .B(G472), .ZN(n431) );
  XOR2_X1 U510 ( .A(n431), .B(KEYINPUT74), .Z(n432) );
  XNOR2_X1 U511 ( .A(n433), .B(n432), .ZN(n536) );
  XNOR2_X1 U512 ( .A(n536), .B(KEYINPUT6), .ZN(n545) );
  NAND2_X1 U513 ( .A1(n494), .A2(n545), .ZN(n435) );
  XNOR2_X1 U514 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n434) );
  XNOR2_X1 U515 ( .A(n435), .B(n434), .ZN(n676) );
  NAND2_X1 U516 ( .A1(n492), .A2(n676), .ZN(n437) );
  XOR2_X1 U517 ( .A(KEYINPUT91), .B(KEYINPUT11), .Z(n442) );
  XOR2_X1 U518 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n439) );
  XNOR2_X1 U519 ( .A(G131), .B(KEYINPUT12), .ZN(n438) );
  XNOR2_X1 U520 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U521 ( .A(n711), .B(n440), .ZN(n441) );
  XNOR2_X1 U522 ( .A(n442), .B(n441), .ZN(n449) );
  AND2_X1 U523 ( .A1(n443), .A2(G214), .ZN(n447) );
  XNOR2_X1 U524 ( .A(G113), .B(G122), .ZN(n445) );
  XOR2_X1 U525 ( .A(G143), .B(G104), .Z(n444) );
  XNOR2_X1 U526 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U527 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U528 ( .A(n449), .B(n448), .ZN(n589) );
  NAND2_X1 U529 ( .A1(n589), .A2(n466), .ZN(n451) );
  XOR2_X1 U530 ( .A(KEYINPUT13), .B(G475), .Z(n450) );
  XNOR2_X1 U531 ( .A(n451), .B(n450), .ZN(n501) );
  INV_X1 U532 ( .A(n501), .ZN(n468) );
  XOR2_X1 U533 ( .A(KEYINPUT96), .B(KEYINPUT93), .Z(n453) );
  XNOR2_X1 U534 ( .A(KEYINPUT7), .B(KEYINPUT94), .ZN(n452) );
  XNOR2_X1 U535 ( .A(n453), .B(n452), .ZN(n455) );
  XOR2_X1 U536 ( .A(KEYINPUT9), .B(G107), .Z(n454) );
  XNOR2_X1 U537 ( .A(n455), .B(n454), .ZN(n458) );
  INV_X1 U538 ( .A(n456), .ZN(n457) );
  XNOR2_X1 U539 ( .A(n458), .B(n457), .ZN(n465) );
  NAND2_X1 U540 ( .A1(G217), .A2(n459), .ZN(n463) );
  XNOR2_X1 U541 ( .A(G116), .B(G122), .ZN(n460) );
  XNOR2_X1 U542 ( .A(KEYINPUT95), .B(n460), .ZN(n461) );
  XNOR2_X1 U543 ( .A(n461), .B(KEYINPUT97), .ZN(n462) );
  XNOR2_X1 U544 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U545 ( .A(n465), .B(n464), .ZN(n607) );
  NAND2_X1 U546 ( .A1(n607), .A2(n466), .ZN(n467) );
  XNOR2_X1 U547 ( .A(n467), .B(G478), .ZN(n474) );
  INV_X1 U548 ( .A(n474), .ZN(n500) );
  OR2_X1 U549 ( .A1(n468), .A2(n500), .ZN(n555) );
  INV_X1 U550 ( .A(n555), .ZN(n469) );
  INV_X1 U551 ( .A(KEYINPUT35), .ZN(n471) );
  INV_X1 U552 ( .A(KEYINPUT44), .ZN(n490) );
  NAND2_X1 U553 ( .A1(n598), .A2(n490), .ZN(n473) );
  XNOR2_X1 U554 ( .A(n473), .B(KEYINPUT67), .ZN(n485) );
  OR2_X1 U555 ( .A1(n501), .A2(n474), .ZN(n669) );
  NOR2_X1 U556 ( .A1(n669), .A2(n652), .ZN(n475) );
  NAND2_X1 U557 ( .A1(n492), .A2(n475), .ZN(n476) );
  INV_X1 U558 ( .A(n545), .ZN(n477) );
  INV_X1 U559 ( .A(KEYINPUT85), .ZN(n479) );
  XNOR2_X1 U560 ( .A(n533), .B(KEYINPUT101), .ZN(n651) );
  XNOR2_X2 U561 ( .A(n489), .B(KEYINPUT32), .ZN(n599) );
  INV_X1 U562 ( .A(n533), .ZN(n480) );
  NAND2_X1 U563 ( .A1(n480), .A2(n536), .ZN(n481) );
  OR2_X1 U564 ( .A1(n658), .A2(n481), .ZN(n482) );
  OR2_X1 U565 ( .A1(n483), .A2(n482), .ZN(n596) );
  NAND2_X1 U566 ( .A1(n485), .A2(n484), .ZN(n487) );
  INV_X1 U567 ( .A(KEYINPUT73), .ZN(n486) );
  XNOR2_X1 U568 ( .A(n487), .B(n486), .ZN(n515) );
  INV_X1 U569 ( .A(KEYINPUT32), .ZN(n488) );
  NAND2_X1 U570 ( .A1(n351), .A2(n348), .ZN(n491) );
  NAND2_X1 U571 ( .A1(n491), .A2(KEYINPUT44), .ZN(n506) );
  BUF_X1 U572 ( .A(n492), .Z(n493) );
  AND2_X1 U573 ( .A1(n494), .A2(n654), .ZN(n662) );
  NAND2_X1 U574 ( .A1(n493), .A2(n662), .ZN(n496) );
  INV_X1 U575 ( .A(KEYINPUT31), .ZN(n495) );
  NAND2_X1 U576 ( .A1(n538), .A2(n657), .ZN(n498) );
  INV_X1 U577 ( .A(KEYINPUT88), .ZN(n497) );
  XNOR2_X1 U578 ( .A(n498), .B(n497), .ZN(n558) );
  AND2_X1 U579 ( .A1(n558), .A2(n536), .ZN(n499) );
  NAND2_X1 U580 ( .A1(n493), .A2(n499), .ZN(n631) );
  NAND2_X1 U581 ( .A1(n644), .A2(n631), .ZN(n503) );
  XOR2_X1 U582 ( .A(KEYINPUT98), .B(n349), .Z(n565) );
  NAND2_X1 U583 ( .A1(n501), .A2(n500), .ZN(n642) );
  NAND2_X1 U584 ( .A1(n565), .A2(n642), .ZN(n502) );
  NAND2_X1 U585 ( .A1(n503), .A2(n670), .ZN(n504) );
  XNOR2_X1 U586 ( .A(n504), .B(KEYINPUT100), .ZN(n505) );
  NAND2_X1 U587 ( .A1(n506), .A2(n505), .ZN(n513) );
  INV_X1 U588 ( .A(KEYINPUT82), .ZN(n507) );
  XNOR2_X1 U589 ( .A(n508), .B(n507), .ZN(n510) );
  NOR2_X1 U590 ( .A1(n658), .A2(n651), .ZN(n509) );
  NAND2_X1 U591 ( .A1(n510), .A2(n509), .ZN(n512) );
  INV_X1 U592 ( .A(KEYINPUT102), .ZN(n511) );
  XNOR2_X1 U593 ( .A(n512), .B(n511), .ZN(n597) );
  NOR2_X1 U594 ( .A1(n513), .A2(n597), .ZN(n514) );
  NAND2_X1 U595 ( .A1(n515), .A2(n514), .ZN(n519) );
  XNOR2_X1 U596 ( .A(KEYINPUT81), .B(KEYINPUT45), .ZN(n517) );
  INV_X1 U597 ( .A(KEYINPUT64), .ZN(n516) );
  XNOR2_X1 U598 ( .A(n517), .B(n516), .ZN(n518) );
  INV_X1 U599 ( .A(n520), .ZN(n521) );
  NAND2_X1 U600 ( .A1(G953), .A2(G900), .ZN(n718) );
  NAND2_X1 U601 ( .A1(n521), .A2(n718), .ZN(n532) );
  NAND2_X1 U602 ( .A1(n654), .A2(n667), .ZN(n522) );
  XNOR2_X1 U603 ( .A(n522), .B(KEYINPUT30), .ZN(n523) );
  NOR2_X1 U604 ( .A1(n532), .A2(n523), .ZN(n557) );
  NAND2_X1 U605 ( .A1(n557), .A2(n530), .ZN(n526) );
  INV_X1 U606 ( .A(n558), .ZN(n525) );
  XNOR2_X1 U607 ( .A(n527), .B(KEYINPUT39), .ZN(n564) );
  NOR2_X1 U608 ( .A1(n564), .A2(n642), .ZN(n529) );
  XNOR2_X1 U609 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n528) );
  XNOR2_X1 U610 ( .A(n529), .B(n528), .ZN(n726) );
  NAND2_X1 U611 ( .A1(n530), .A2(n667), .ZN(n671) );
  XNOR2_X1 U612 ( .A(KEYINPUT41), .B(n531), .ZN(n685) );
  NOR2_X1 U613 ( .A1(n533), .A2(n532), .ZN(n535) );
  NAND2_X1 U614 ( .A1(n535), .A2(n534), .ZN(n543) );
  NOR2_X1 U615 ( .A1(n543), .A2(n536), .ZN(n537) );
  XNOR2_X1 U616 ( .A(n537), .B(KEYINPUT28), .ZN(n539) );
  NAND2_X1 U617 ( .A1(n539), .A2(n538), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT42), .B(n540), .Z(n541) );
  NAND2_X1 U619 ( .A1(n726), .A2(n722), .ZN(n542) );
  XNOR2_X1 U620 ( .A(n542), .B(KEYINPUT46), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n642), .A2(n543), .ZN(n544) );
  AND2_X1 U622 ( .A1(n545), .A2(n544), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n566), .A2(n546), .ZN(n547) );
  XOR2_X1 U624 ( .A(KEYINPUT36), .B(n547), .Z(n548) );
  NAND2_X1 U625 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U626 ( .A(n550), .B(KEYINPUT105), .ZN(n723) );
  NOR2_X1 U627 ( .A1(n552), .A2(n551), .ZN(n640) );
  NAND2_X1 U628 ( .A1(n670), .A2(n640), .ZN(n553) );
  XNOR2_X1 U629 ( .A(KEYINPUT47), .B(n553), .ZN(n554) );
  NOR2_X1 U630 ( .A1(n723), .A2(n554), .ZN(n560) );
  NOR2_X1 U631 ( .A1(n555), .A2(n344), .ZN(n556) );
  AND2_X1 U632 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U633 ( .A1(n559), .A2(n558), .ZN(n638) );
  NAND2_X1 U634 ( .A1(n560), .A2(n638), .ZN(n561) );
  XNOR2_X1 U635 ( .A(n563), .B(KEYINPUT48), .ZN(n571) );
  NOR2_X1 U636 ( .A1(n565), .A2(n564), .ZN(n648) );
  NAND2_X1 U637 ( .A1(n566), .A2(n667), .ZN(n567) );
  OR2_X1 U638 ( .A1(n658), .A2(n567), .ZN(n568) );
  XNOR2_X1 U639 ( .A(n568), .B(KEYINPUT43), .ZN(n569) );
  AND2_X1 U640 ( .A1(n569), .A2(n344), .ZN(n595) );
  NOR2_X1 U641 ( .A1(n648), .A2(n595), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n714) );
  NAND2_X1 U643 ( .A1(n702), .A2(n576), .ZN(n574) );
  INV_X1 U644 ( .A(KEYINPUT2), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n579) );
  XNOR2_X1 U646 ( .A(KEYINPUT77), .B(KEYINPUT2), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n577), .A2(n702), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n649) );
  INV_X1 U649 ( .A(n580), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n617), .A2(G217), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n584), .B(n583), .ZN(n586) );
  INV_X1 U652 ( .A(G952), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n624), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(G66) );
  NAND2_X1 U655 ( .A1(n617), .A2(G475), .ZN(n591) );
  XOR2_X1 U656 ( .A(n589), .B(KEYINPUT59), .Z(n590) );
  XNOR2_X1 U657 ( .A(n591), .B(n590), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n592), .A2(n624), .ZN(n594) );
  INV_X1 U659 ( .A(KEYINPUT60), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n594), .B(n593), .ZN(G60) );
  XOR2_X1 U661 ( .A(G140), .B(n595), .Z(G42) );
  XNOR2_X1 U662 ( .A(n596), .B(G110), .ZN(G12) );
  XOR2_X1 U663 ( .A(G101), .B(n597), .Z(G3) );
  XNOR2_X1 U664 ( .A(n343), .B(G122), .ZN(G24) );
  XNOR2_X1 U665 ( .A(n599), .B(G119), .ZN(G21) );
  NAND2_X1 U666 ( .A1(n347), .A2(G472), .ZN(n603) );
  XOR2_X1 U667 ( .A(KEYINPUT106), .B(KEYINPUT62), .Z(n600) );
  XNOR2_X1 U668 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U669 ( .A(n603), .B(n602), .ZN(n604) );
  NAND2_X1 U670 ( .A1(n604), .A2(n624), .ZN(n605) );
  XNOR2_X1 U671 ( .A(n605), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U672 ( .A1(n347), .A2(G478), .ZN(n606) );
  XOR2_X1 U673 ( .A(n607), .B(n606), .Z(n608) );
  INV_X1 U674 ( .A(n624), .ZN(n615) );
  NOR2_X1 U675 ( .A1(n608), .A2(n615), .ZN(G63) );
  BUF_X1 U676 ( .A(n346), .Z(n609) );
  NAND2_X1 U677 ( .A1(n609), .A2(G469), .ZN(n614) );
  XNOR2_X1 U678 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n610) );
  XNOR2_X1 U679 ( .A(n610), .B(KEYINPUT58), .ZN(n611) );
  XNOR2_X1 U680 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U681 ( .A(n614), .B(n613), .ZN(n616) );
  NOR2_X1 U682 ( .A1(n616), .A2(n615), .ZN(G54) );
  NAND2_X1 U683 ( .A1(n346), .A2(G210), .ZN(n623) );
  BUF_X1 U684 ( .A(n618), .Z(n621) );
  XNOR2_X1 U685 ( .A(KEYINPUT117), .B(KEYINPUT54), .ZN(n619) );
  XOR2_X1 U686 ( .A(n619), .B(KEYINPUT55), .Z(n620) );
  XNOR2_X1 U687 ( .A(n623), .B(n622), .ZN(n625) );
  NAND2_X1 U688 ( .A1(n625), .A2(n624), .ZN(n627) );
  XOR2_X1 U689 ( .A(KEYINPUT118), .B(KEYINPUT56), .Z(n626) );
  XNOR2_X1 U690 ( .A(n627), .B(n626), .ZN(G51) );
  NOR2_X1 U691 ( .A1(n642), .A2(n631), .ZN(n629) );
  XNOR2_X1 U692 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n628) );
  XNOR2_X1 U693 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U694 ( .A(G104), .B(n630), .ZN(G6) );
  INV_X1 U695 ( .A(n349), .ZN(n645) );
  NOR2_X1 U696 ( .A1(n645), .A2(n631), .ZN(n633) );
  XNOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n632) );
  XNOR2_X1 U698 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U699 ( .A(G107), .B(n634), .ZN(G9) );
  XOR2_X1 U700 ( .A(KEYINPUT109), .B(KEYINPUT29), .Z(n636) );
  NAND2_X1 U701 ( .A1(n640), .A2(n349), .ZN(n635) );
  XNOR2_X1 U702 ( .A(n636), .B(n635), .ZN(n637) );
  XOR2_X1 U703 ( .A(G128), .B(n637), .Z(G30) );
  XNOR2_X1 U704 ( .A(G143), .B(n638), .ZN(G45) );
  INV_X1 U705 ( .A(n642), .ZN(n639) );
  NAND2_X1 U706 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U707 ( .A(G146), .B(n641), .ZN(G48) );
  NOR2_X1 U708 ( .A1(n642), .A2(n644), .ZN(n643) );
  XOR2_X1 U709 ( .A(G113), .B(n643), .Z(G15) );
  NOR2_X1 U710 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U711 ( .A(KEYINPUT110), .B(n646), .Z(n647) );
  XNOR2_X1 U712 ( .A(G116), .B(n647), .ZN(G18) );
  XOR2_X1 U713 ( .A(G134), .B(n648), .Z(G36) );
  BUF_X1 U714 ( .A(n649), .Z(n691) );
  NAND2_X1 U715 ( .A1(G952), .A2(n650), .ZN(n683) );
  XOR2_X1 U716 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n665) );
  NAND2_X1 U717 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U718 ( .A(KEYINPUT49), .B(n653), .ZN(n655) );
  NOR2_X1 U719 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U720 ( .A(KEYINPUT112), .B(n656), .Z(n661) );
  NOR2_X1 U721 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U722 ( .A(n659), .B(KEYINPUT50), .ZN(n660) );
  NOR2_X1 U723 ( .A1(n661), .A2(n660), .ZN(n663) );
  OR2_X1 U724 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U725 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U726 ( .A1(n666), .A2(n685), .ZN(n679) );
  NOR2_X1 U727 ( .A1(n530), .A2(n667), .ZN(n668) );
  NOR2_X1 U728 ( .A1(n669), .A2(n668), .ZN(n675) );
  INV_X1 U729 ( .A(n670), .ZN(n672) );
  NOR2_X1 U730 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U731 ( .A(n673), .B(KEYINPUT114), .ZN(n674) );
  NOR2_X1 U732 ( .A1(n675), .A2(n674), .ZN(n677) );
  INV_X1 U733 ( .A(n676), .ZN(n684) );
  NOR2_X1 U734 ( .A1(n677), .A2(n684), .ZN(n678) );
  NOR2_X1 U735 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U736 ( .A(KEYINPUT52), .B(n680), .Z(n681) );
  XNOR2_X1 U737 ( .A(KEYINPUT115), .B(n681), .ZN(n682) );
  NOR2_X1 U738 ( .A1(n683), .A2(n682), .ZN(n687) );
  NOR2_X1 U739 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U740 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U741 ( .A(n688), .B(KEYINPUT116), .ZN(n689) );
  NAND2_X1 U742 ( .A1(n689), .A2(n703), .ZN(n690) );
  NOR2_X1 U743 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U744 ( .A(n692), .B(KEYINPUT53), .ZN(G75) );
  BUF_X1 U745 ( .A(n693), .Z(n694) );
  XNOR2_X1 U746 ( .A(G101), .B(KEYINPUT124), .ZN(n695) );
  XNOR2_X1 U747 ( .A(n694), .B(n695), .ZN(n697) );
  NOR2_X1 U748 ( .A1(G898), .A2(n703), .ZN(n696) );
  NOR2_X1 U749 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U750 ( .A(n698), .B(KEYINPUT123), .Z(n710) );
  NAND2_X1 U751 ( .A1(G953), .A2(G224), .ZN(n699) );
  XNOR2_X1 U752 ( .A(KEYINPUT61), .B(n699), .ZN(n700) );
  NAND2_X1 U753 ( .A1(n700), .A2(G898), .ZN(n701) );
  XNOR2_X1 U754 ( .A(KEYINPUT121), .B(n701), .ZN(n707) );
  BUF_X1 U755 ( .A(n702), .Z(n704) );
  NAND2_X1 U756 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U757 ( .A(KEYINPUT122), .B(n705), .Z(n706) );
  NOR2_X1 U758 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n708), .B(KEYINPUT125), .ZN(n709) );
  XNOR2_X1 U760 ( .A(n710), .B(n709), .ZN(G69) );
  XNOR2_X1 U761 ( .A(n711), .B(KEYINPUT126), .ZN(n712) );
  XNOR2_X1 U762 ( .A(n713), .B(n712), .ZN(n716) );
  XNOR2_X1 U763 ( .A(n716), .B(n714), .ZN(n715) );
  NOR2_X1 U764 ( .A1(G953), .A2(n715), .ZN(n720) );
  XOR2_X1 U765 ( .A(G227), .B(n716), .Z(n717) );
  NOR2_X1 U766 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U767 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U768 ( .A(KEYINPUT127), .B(n721), .Z(G72) );
  XNOR2_X1 U769 ( .A(G137), .B(n722), .ZN(G39) );
  XOR2_X1 U770 ( .A(KEYINPUT37), .B(KEYINPUT111), .Z(n725) );
  XNOR2_X1 U771 ( .A(G125), .B(n723), .ZN(n724) );
  XNOR2_X1 U772 ( .A(n725), .B(n724), .ZN(G27) );
  XNOR2_X1 U773 ( .A(G131), .B(n726), .ZN(G33) );
endmodule

