

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725;

  NOR2_X1 U379 ( .A1(n673), .A2(n688), .ZN(n379) );
  XNOR2_X1 U380 ( .A(n572), .B(n385), .ZN(n553) );
  NOR2_X1 U381 ( .A1(n516), .A2(n517), .ZN(n359) );
  NOR2_X1 U382 ( .A1(n678), .A2(n688), .ZN(n380) );
  OR2_X2 U383 ( .A1(n527), .A2(n526), .ZN(n382) );
  XNOR2_X2 U384 ( .A(n391), .B(KEYINPUT35), .ZN(n715) );
  NOR2_X1 U385 ( .A1(n656), .A2(n519), .ZN(n393) );
  XNOR2_X2 U386 ( .A(n540), .B(n541), .ZN(n577) );
  XNOR2_X2 U387 ( .A(n450), .B(n414), .ZN(n592) );
  NOR2_X2 U388 ( .A1(n686), .A2(G902), .ZN(n500) );
  NOR2_X1 U389 ( .A1(n553), .A2(n458), .ZN(n459) );
  NOR2_X1 U390 ( .A1(n669), .A2(n668), .ZN(n375) );
  AND2_X2 U391 ( .A1(n602), .A2(n631), .ZN(n684) );
  NOR2_X1 U392 ( .A1(n692), .A2(KEYINPUT2), .ZN(n629) );
  BUF_X1 U393 ( .A(n628), .Z(n692) );
  NOR2_X1 U394 ( .A1(n511), .A2(n510), .ZN(n528) );
  NAND2_X1 U395 ( .A1(n378), .A2(n359), .ZN(n410) );
  XNOR2_X1 U396 ( .A(n485), .B(KEYINPUT22), .ZN(n504) );
  XNOR2_X1 U397 ( .A(n459), .B(KEYINPUT0), .ZN(n523) );
  AND2_X1 U398 ( .A1(n538), .A2(n537), .ZN(n563) );
  OR2_X1 U399 ( .A1(n486), .A2(G902), .ZN(n487) );
  XNOR2_X1 U400 ( .A(n499), .B(n361), .ZN(n399) );
  XNOR2_X1 U401 ( .A(n467), .B(n404), .ZN(n496) );
  XNOR2_X1 U402 ( .A(n473), .B(n386), .ZN(n704) );
  XNOR2_X1 U403 ( .A(n431), .B(G122), .ZN(n465) );
  XNOR2_X1 U404 ( .A(n439), .B(G134), .ZN(n473) );
  XNOR2_X1 U405 ( .A(n372), .B(G107), .ZN(n430) );
  XNOR2_X1 U406 ( .A(G143), .B(G128), .ZN(n439) );
  XNOR2_X1 U407 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n422) );
  XOR2_X1 U408 ( .A(G137), .B(G140), .Z(n495) );
  XNOR2_X1 U409 ( .A(n432), .B(n465), .ZN(n435) );
  XNOR2_X1 U410 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U411 ( .A(KEYINPUT71), .B(KEYINPUT16), .Z(n429) );
  XNOR2_X1 U412 ( .A(n704), .B(n413), .ZN(n427) );
  XNOR2_X1 U413 ( .A(n445), .B(G146), .ZN(n413) );
  NAND2_X1 U414 ( .A1(n383), .A2(n381), .ZN(n529) );
  XNOR2_X1 U415 ( .A(n382), .B(KEYINPUT83), .ZN(n381) );
  NOR2_X1 U416 ( .A1(n528), .A2(n360), .ZN(n383) );
  INV_X1 U417 ( .A(n714), .ZN(n407) );
  XOR2_X1 U418 ( .A(KEYINPUT5), .B(G113), .Z(n425) );
  XNOR2_X1 U419 ( .A(n388), .B(n387), .ZN(n386) );
  INV_X1 U420 ( .A(KEYINPUT4), .ZN(n387) );
  XNOR2_X1 U421 ( .A(G131), .B(KEYINPUT68), .ZN(n388) );
  INV_X1 U422 ( .A(G110), .ZN(n372) );
  AND2_X1 U423 ( .A1(n576), .A2(n719), .ZN(n401) );
  XNOR2_X1 U424 ( .A(n584), .B(n368), .ZN(n409) );
  NOR2_X1 U425 ( .A1(n547), .A2(n546), .ZN(n569) );
  INV_X1 U426 ( .A(G469), .ZN(n412) );
  XOR2_X1 U427 ( .A(G122), .B(KEYINPUT9), .Z(n476) );
  XNOR2_X1 U428 ( .A(n470), .B(n403), .ZN(n675) );
  XNOR2_X1 U429 ( .A(n405), .B(n496), .ZN(n403) );
  XNOR2_X1 U430 ( .A(n465), .B(n469), .ZN(n405) );
  NAND2_X1 U431 ( .A1(n628), .A2(n601), .ZN(n631) );
  XNOR2_X1 U432 ( .A(n600), .B(KEYINPUT79), .ZN(n601) );
  XNOR2_X1 U433 ( .A(n481), .B(n480), .ZN(n517) );
  XNOR2_X1 U434 ( .A(n515), .B(n402), .ZN(n516) );
  INV_X1 U435 ( .A(KEYINPUT94), .ZN(n402) );
  OR2_X2 U436 ( .A1(n608), .A2(G902), .ZN(n389) );
  NAND2_X1 U437 ( .A1(n373), .A2(n636), .ZN(n512) );
  INV_X1 U438 ( .A(n504), .ZN(n373) );
  NOR2_X1 U439 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U440 ( .A(n398), .B(KEYINPUT15), .ZN(n596) );
  XNOR2_X1 U441 ( .A(KEYINPUT85), .B(G902), .ZN(n398) );
  XNOR2_X1 U442 ( .A(G113), .B(G104), .ZN(n431) );
  XNOR2_X1 U443 ( .A(G140), .B(KEYINPUT12), .ZN(n460) );
  XOR2_X1 U444 ( .A(KEYINPUT93), .B(KEYINPUT11), .Z(n461) );
  XNOR2_X1 U445 ( .A(G143), .B(G131), .ZN(n463) );
  INV_X1 U446 ( .A(KEYINPUT10), .ZN(n404) );
  XNOR2_X1 U447 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n441) );
  XOR2_X1 U448 ( .A(KEYINPUT17), .B(KEYINPUT75), .Z(n442) );
  OR2_X1 U449 ( .A1(G237), .A2(G902), .ZN(n451) );
  XNOR2_X1 U450 ( .A(n471), .B(n472), .ZN(n515) );
  XNOR2_X1 U451 ( .A(n390), .B(n427), .ZN(n608) );
  XNOR2_X1 U452 ( .A(n419), .B(n427), .ZN(n486) );
  XNOR2_X1 U453 ( .A(KEYINPUT97), .B(KEYINPUT33), .ZN(n507) );
  INV_X1 U454 ( .A(KEYINPUT19), .ZN(n385) );
  INV_X1 U455 ( .A(n518), .ZN(n411) );
  INV_X1 U456 ( .A(n592), .ZN(n560) );
  INV_X1 U457 ( .A(n547), .ZN(n535) );
  INV_X1 U458 ( .A(n688), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n479), .B(n376), .ZN(n680) );
  XNOR2_X1 U460 ( .A(n473), .B(n478), .ZN(n376) );
  XNOR2_X1 U461 ( .A(G116), .B(G107), .ZN(n478) );
  XNOR2_X1 U462 ( .A(n675), .B(n370), .ZN(n676) );
  XNOR2_X1 U463 ( .A(n670), .B(n369), .ZN(n671) );
  NOR2_X1 U464 ( .A1(G952), .A2(n474), .ZN(n688) );
  AND2_X1 U465 ( .A1(n631), .A2(n363), .ZN(n374) );
  NOR2_X1 U466 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U467 ( .A(n577), .ZN(n378) );
  NOR2_X1 U468 ( .A1(n512), .A2(n571), .ZN(n384) );
  AND2_X1 U469 ( .A1(n511), .A2(KEYINPUT44), .ZN(n360) );
  XNOR2_X1 U470 ( .A(KEYINPUT90), .B(KEYINPUT25), .ZN(n361) );
  NOR2_X1 U471 ( .A1(n625), .A2(n359), .ZN(n362) );
  OR2_X1 U472 ( .A1(n630), .A2(KEYINPUT2), .ZN(n363) );
  XOR2_X1 U473 ( .A(n561), .B(KEYINPUT76), .Z(n364) );
  XOR2_X1 U474 ( .A(n629), .B(KEYINPUT78), .Z(n365) );
  AND2_X1 U475 ( .A1(n468), .A2(G210), .ZN(n366) );
  XOR2_X1 U476 ( .A(n608), .B(n607), .Z(n367) );
  XOR2_X1 U477 ( .A(n583), .B(KEYINPUT81), .Z(n368) );
  INV_X2 U478 ( .A(G953), .ZN(n474) );
  XNOR2_X1 U479 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n369) );
  XNOR2_X1 U480 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n370) );
  XOR2_X1 U481 ( .A(n609), .B(KEYINPUT84), .Z(n371) );
  XNOR2_X1 U482 ( .A(n384), .B(KEYINPUT82), .ZN(n513) );
  NAND2_X1 U483 ( .A1(n513), .A2(n634), .ZN(n611) );
  NAND2_X1 U484 ( .A1(n670), .A2(n594), .ZN(n450) );
  XNOR2_X1 U485 ( .A(n689), .B(n448), .ZN(n670) );
  NAND2_X1 U486 ( .A1(n617), .A2(n718), .ZN(n511) );
  NAND2_X1 U487 ( .A1(n506), .A2(n545), .ZN(n617) );
  NAND2_X1 U488 ( .A1(n365), .A2(n374), .ZN(n632) );
  NOR2_X1 U489 ( .A1(n715), .A2(KEYINPUT44), .ZN(n509) );
  XNOR2_X1 U490 ( .A(n375), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U491 ( .A(n426), .B(n366), .ZN(n390) );
  NOR2_X2 U492 ( .A1(n594), .A2(n705), .ZN(n595) );
  XNOR2_X1 U493 ( .A(n377), .B(n476), .ZN(n477) );
  NAND2_X1 U494 ( .A1(n488), .A2(G217), .ZN(n377) );
  AND2_X1 U495 ( .A1(n722), .A2(n407), .ZN(n406) );
  XNOR2_X1 U496 ( .A(n379), .B(n674), .ZN(G51) );
  XNOR2_X1 U497 ( .A(n380), .B(n679), .ZN(G60) );
  NAND2_X1 U498 ( .A1(n592), .A2(n649), .ZN(n572) );
  XNOR2_X2 U499 ( .A(n389), .B(G472), .ZN(n548) );
  NAND2_X1 U500 ( .A1(n392), .A2(n364), .ZN(n391) );
  XNOR2_X1 U501 ( .A(n393), .B(KEYINPUT34), .ZN(n392) );
  XNOR2_X1 U502 ( .A(n394), .B(n371), .ZN(G57) );
  NAND2_X1 U503 ( .A1(n396), .A2(n395), .ZN(n394) );
  XNOR2_X1 U504 ( .A(n397), .B(n367), .ZN(n396) );
  NAND2_X1 U505 ( .A1(n684), .A2(G472), .ZN(n397) );
  INV_X1 U506 ( .A(n634), .ZN(n545) );
  XNOR2_X2 U507 ( .A(n500), .B(n399), .ZN(n634) );
  XNOR2_X1 U508 ( .A(n400), .B(n585), .ZN(n408) );
  NAND2_X1 U509 ( .A1(n401), .A2(n409), .ZN(n400) );
  AND2_X2 U510 ( .A1(n408), .A2(n406), .ZN(n630) );
  XNOR2_X2 U511 ( .A(n423), .B(n422), .ZN(n434) );
  NAND2_X1 U512 ( .A1(n723), .A2(n724), .ZN(n584) );
  XNOR2_X2 U513 ( .A(n410), .B(KEYINPUT40), .ZN(n723) );
  NAND2_X1 U514 ( .A1(n551), .A2(n411), .ZN(n552) );
  XNOR2_X2 U515 ( .A(n487), .B(n412), .ZN(n518) );
  XNOR2_X2 U516 ( .A(n548), .B(n428), .ZN(n571) );
  XNOR2_X1 U517 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U518 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U519 ( .A(n518), .B(KEYINPUT1), .ZN(n636) );
  XOR2_X1 U520 ( .A(n449), .B(KEYINPUT86), .Z(n414) );
  INV_X1 U521 ( .A(KEYINPUT46), .ZN(n583) );
  INV_X1 U522 ( .A(KEYINPUT48), .ZN(n585) );
  XNOR2_X1 U523 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U524 ( .A(n508), .B(n507), .ZN(n656) );
  INV_X1 U525 ( .A(n636), .ZN(n589) );
  XNOR2_X1 U526 ( .A(n494), .B(n493), .ZN(n497) );
  XNOR2_X1 U527 ( .A(KEYINPUT58), .B(KEYINPUT117), .ZN(n421) );
  XOR2_X1 U528 ( .A(KEYINPUT66), .B(G101), .Z(n445) );
  NAND2_X1 U529 ( .A1(n474), .A2(G227), .ZN(n415) );
  XNOR2_X1 U530 ( .A(n415), .B(n495), .ZN(n416) );
  XOR2_X1 U531 ( .A(n416), .B(G104), .Z(n418) );
  XNOR2_X1 U532 ( .A(n430), .B(KEYINPUT74), .ZN(n417) );
  XNOR2_X1 U533 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U534 ( .A(n486), .B(KEYINPUT57), .ZN(n420) );
  XNOR2_X1 U535 ( .A(n421), .B(n420), .ZN(n604) );
  XOR2_X2 U536 ( .A(G116), .B(G119), .Z(n423) );
  XNOR2_X1 U537 ( .A(n434), .B(G137), .ZN(n424) );
  XNOR2_X1 U538 ( .A(n425), .B(n424), .ZN(n426) );
  NOR2_X1 U539 ( .A1(G953), .A2(G237), .ZN(n468) );
  INV_X1 U540 ( .A(KEYINPUT6), .ZN(n428) );
  INV_X1 U541 ( .A(n596), .ZN(n594) );
  INV_X1 U542 ( .A(n435), .ZN(n433) );
  NAND2_X1 U543 ( .A1(n434), .A2(n433), .ZN(n438) );
  INV_X1 U544 ( .A(n434), .ZN(n436) );
  NAND2_X1 U545 ( .A1(n436), .A2(n435), .ZN(n437) );
  NAND2_X1 U546 ( .A1(n438), .A2(n437), .ZN(n689) );
  NAND2_X1 U547 ( .A1(G224), .A2(n474), .ZN(n440) );
  XNOR2_X1 U548 ( .A(n440), .B(n439), .ZN(n444) );
  XNOR2_X1 U549 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U550 ( .A(n444), .B(n443), .ZN(n447) );
  XNOR2_X1 U551 ( .A(G146), .B(G125), .ZN(n466) );
  XNOR2_X1 U552 ( .A(n445), .B(n466), .ZN(n446) );
  NAND2_X1 U553 ( .A1(n451), .A2(G210), .ZN(n449) );
  NAND2_X1 U554 ( .A1(G214), .A2(n451), .ZN(n649) );
  XOR2_X1 U555 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n453) );
  NAND2_X1 U556 ( .A1(G234), .A2(G237), .ZN(n452) );
  XNOR2_X1 U557 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U558 ( .A1(G952), .A2(n454), .ZN(n662) );
  NOR2_X1 U559 ( .A1(G953), .A2(n662), .ZN(n534) );
  NAND2_X1 U560 ( .A1(G902), .A2(n454), .ZN(n455) );
  XOR2_X1 U561 ( .A(KEYINPUT88), .B(n455), .Z(n456) );
  NAND2_X1 U562 ( .A1(G953), .A2(n456), .ZN(n532) );
  NOR2_X1 U563 ( .A1(G898), .A2(n532), .ZN(n457) );
  NOR2_X1 U564 ( .A1(n534), .A2(n457), .ZN(n458) );
  XNOR2_X1 U565 ( .A(KEYINPUT13), .B(G475), .ZN(n472) );
  XNOR2_X1 U566 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U567 ( .A(n462), .B(KEYINPUT92), .Z(n464) );
  XNOR2_X1 U568 ( .A(n464), .B(n463), .ZN(n470) );
  INV_X1 U569 ( .A(n466), .ZN(n467) );
  NAND2_X1 U570 ( .A1(G214), .A2(n468), .ZN(n469) );
  NOR2_X1 U571 ( .A1(G902), .A2(n675), .ZN(n471) );
  NAND2_X1 U572 ( .A1(G234), .A2(n474), .ZN(n475) );
  XOR2_X1 U573 ( .A(KEYINPUT8), .B(n475), .Z(n488) );
  XOR2_X1 U574 ( .A(n477), .B(KEYINPUT7), .Z(n479) );
  NOR2_X1 U575 ( .A1(G902), .A2(n680), .ZN(n481) );
  XNOR2_X1 U576 ( .A(KEYINPUT95), .B(G478), .ZN(n480) );
  NOR2_X1 U577 ( .A1(n515), .A2(n517), .ZN(n578) );
  NAND2_X1 U578 ( .A1(n594), .A2(G234), .ZN(n482) );
  XNOR2_X1 U579 ( .A(n482), .B(KEYINPUT20), .ZN(n498) );
  NAND2_X1 U580 ( .A1(n498), .A2(G221), .ZN(n483) );
  XOR2_X1 U581 ( .A(KEYINPUT21), .B(n483), .Z(n633) );
  AND2_X1 U582 ( .A1(n578), .A2(n633), .ZN(n484) );
  NAND2_X1 U583 ( .A1(n523), .A2(n484), .ZN(n485) );
  NOR2_X1 U584 ( .A1(n571), .A2(n504), .ZN(n502) );
  NAND2_X1 U585 ( .A1(G221), .A2(n488), .ZN(n494) );
  XOR2_X1 U586 ( .A(KEYINPUT89), .B(G110), .Z(n490) );
  XNOR2_X1 U587 ( .A(G128), .B(G119), .ZN(n489) );
  XNOR2_X1 U588 ( .A(n490), .B(n489), .ZN(n492) );
  XOR2_X1 U589 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n491) );
  XNOR2_X1 U590 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U591 ( .A(n496), .B(n495), .ZN(n701) );
  XNOR2_X1 U592 ( .A(n497), .B(n701), .ZN(n686) );
  NAND2_X1 U593 ( .A1(n498), .A2(G217), .ZN(n499) );
  NOR2_X1 U594 ( .A1(n636), .A2(n634), .ZN(n501) );
  NAND2_X1 U595 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U596 ( .A(KEYINPUT32), .B(n503), .ZN(n718) );
  XNOR2_X1 U597 ( .A(KEYINPUT96), .B(n512), .ZN(n505) );
  NOR2_X1 U598 ( .A1(n548), .A2(n505), .ZN(n506) );
  NAND2_X1 U599 ( .A1(n633), .A2(n634), .ZN(n637) );
  NOR2_X1 U600 ( .A1(n636), .A2(n637), .ZN(n522) );
  NAND2_X1 U601 ( .A1(n522), .A2(n571), .ZN(n508) );
  INV_X1 U602 ( .A(n523), .ZN(n519) );
  NAND2_X1 U603 ( .A1(n515), .A2(n517), .ZN(n561) );
  XNOR2_X1 U604 ( .A(n509), .B(KEYINPUT67), .ZN(n510) );
  NAND2_X1 U605 ( .A1(n715), .A2(KEYINPUT44), .ZN(n514) );
  NAND2_X1 U606 ( .A1(n611), .A2(n514), .ZN(n527) );
  NAND2_X1 U607 ( .A1(n517), .A2(n516), .ZN(n542) );
  INV_X1 U608 ( .A(n542), .ZN(n625) );
  NOR2_X2 U609 ( .A1(n518), .A2(n637), .ZN(n531) );
  NOR2_X1 U610 ( .A1(n548), .A2(n519), .ZN(n520) );
  NAND2_X1 U611 ( .A1(n531), .A2(n520), .ZN(n521) );
  XNOR2_X1 U612 ( .A(KEYINPUT91), .B(n521), .ZN(n613) );
  AND2_X1 U613 ( .A1(n548), .A2(n522), .ZN(n644) );
  NAND2_X1 U614 ( .A1(n523), .A2(n644), .ZN(n524) );
  XNOR2_X1 U615 ( .A(n524), .B(KEYINPUT31), .ZN(n626) );
  NOR2_X1 U616 ( .A1(n613), .A2(n626), .ZN(n525) );
  NOR2_X1 U617 ( .A1(n362), .A2(n525), .ZN(n526) );
  XNOR2_X2 U618 ( .A(n529), .B(KEYINPUT45), .ZN(n628) );
  XOR2_X1 U619 ( .A(KEYINPUT70), .B(KEYINPUT39), .Z(n541) );
  NAND2_X1 U620 ( .A1(n548), .A2(n649), .ZN(n530) );
  XOR2_X1 U621 ( .A(n530), .B(KEYINPUT30), .Z(n538) );
  XOR2_X1 U622 ( .A(KEYINPUT99), .B(n531), .Z(n536) );
  NOR2_X1 U623 ( .A1(G900), .A2(n532), .ZN(n533) );
  NOR2_X1 U624 ( .A1(n534), .A2(n533), .ZN(n547) );
  AND2_X1 U625 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U626 ( .A(KEYINPUT38), .B(KEYINPUT73), .ZN(n539) );
  XOR2_X1 U627 ( .A(n539), .B(n560), .Z(n648) );
  NAND2_X1 U628 ( .A1(n563), .A2(n648), .ZN(n540) );
  NOR2_X1 U629 ( .A1(n577), .A2(n542), .ZN(n543) );
  XOR2_X1 U630 ( .A(KEYINPUT105), .B(n543), .Z(n714) );
  INV_X1 U631 ( .A(KEYINPUT77), .ZN(n544) );
  NAND2_X1 U632 ( .A1(n544), .A2(n362), .ZN(n554) );
  NAND2_X1 U633 ( .A1(n545), .A2(n633), .ZN(n546) );
  NAND2_X1 U634 ( .A1(n569), .A2(n548), .ZN(n550) );
  XNOR2_X1 U635 ( .A(KEYINPUT101), .B(KEYINPUT28), .ZN(n549) );
  XNOR2_X1 U636 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U637 ( .A(KEYINPUT102), .B(n552), .ZN(n580) );
  NOR2_X2 U638 ( .A1(n580), .A2(n553), .ZN(n622) );
  NAND2_X1 U639 ( .A1(n554), .A2(n622), .ZN(n555) );
  NAND2_X1 U640 ( .A1(n555), .A2(KEYINPUT47), .ZN(n558) );
  NOR2_X1 U641 ( .A1(n362), .A2(KEYINPUT47), .ZN(n556) );
  NAND2_X1 U642 ( .A1(n556), .A2(n622), .ZN(n557) );
  NAND2_X1 U643 ( .A1(n558), .A2(n557), .ZN(n567) );
  NAND2_X1 U644 ( .A1(KEYINPUT47), .A2(n362), .ZN(n559) );
  NAND2_X1 U645 ( .A1(n559), .A2(KEYINPUT77), .ZN(n565) );
  NOR2_X1 U646 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U647 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U648 ( .A(KEYINPUT100), .B(n564), .ZN(n716) );
  NAND2_X1 U649 ( .A1(n565), .A2(n716), .ZN(n566) );
  XNOR2_X1 U650 ( .A(KEYINPUT72), .B(n568), .ZN(n576) );
  AND2_X1 U651 ( .A1(n359), .A2(n569), .ZN(n570) );
  NAND2_X1 U652 ( .A1(n571), .A2(n570), .ZN(n586) );
  NOR2_X1 U653 ( .A1(n572), .A2(n586), .ZN(n573) );
  XNOR2_X1 U654 ( .A(KEYINPUT36), .B(n573), .ZN(n574) );
  NAND2_X1 U655 ( .A1(n574), .A2(n589), .ZN(n575) );
  XNOR2_X1 U656 ( .A(n575), .B(KEYINPUT104), .ZN(n719) );
  INV_X1 U657 ( .A(n578), .ZN(n652) );
  NAND2_X1 U658 ( .A1(n649), .A2(n648), .ZN(n653) );
  NOR2_X1 U659 ( .A1(n652), .A2(n653), .ZN(n579) );
  XNOR2_X1 U660 ( .A(KEYINPUT41), .B(n579), .ZN(n664) );
  NOR2_X1 U661 ( .A1(n580), .A2(n664), .ZN(n582) );
  XNOR2_X1 U662 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n581) );
  XNOR2_X1 U663 ( .A(n582), .B(n581), .ZN(n724) );
  INV_X1 U664 ( .A(n586), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n587), .A2(n649), .ZN(n588) );
  NOR2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U667 ( .A(n590), .B(KEYINPUT43), .ZN(n591) );
  XOR2_X1 U668 ( .A(KEYINPUT98), .B(n593), .Z(n722) );
  INV_X1 U669 ( .A(n630), .ZN(n705) );
  NAND2_X1 U670 ( .A1(n628), .A2(n595), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n596), .A2(KEYINPUT2), .ZN(n597) );
  XNOR2_X1 U672 ( .A(KEYINPUT64), .B(n597), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n630), .A2(KEYINPUT2), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n684), .A2(G469), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(n605) );
  NOR2_X2 U677 ( .A1(n605), .A2(n688), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n606), .B(KEYINPUT118), .ZN(G54) );
  XNOR2_X1 U679 ( .A(KEYINPUT106), .B(KEYINPUT62), .ZN(n607) );
  INV_X1 U680 ( .A(KEYINPUT63), .ZN(n609) );
  XOR2_X1 U681 ( .A(G101), .B(KEYINPUT107), .Z(n610) );
  XNOR2_X1 U682 ( .A(n611), .B(n610), .ZN(G3) );
  NAND2_X1 U683 ( .A1(n613), .A2(n359), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n612), .B(G104), .ZN(G6) );
  XOR2_X1 U685 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n615) );
  NAND2_X1 U686 ( .A1(n613), .A2(n625), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U688 ( .A(G107), .B(n616), .ZN(G9) );
  XNOR2_X1 U689 ( .A(G110), .B(n617), .ZN(G12) );
  XOR2_X1 U690 ( .A(KEYINPUT29), .B(KEYINPUT109), .Z(n619) );
  NAND2_X1 U691 ( .A1(n622), .A2(n625), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n619), .B(n618), .ZN(n621) );
  XOR2_X1 U693 ( .A(G128), .B(KEYINPUT108), .Z(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(G30) );
  NAND2_X1 U695 ( .A1(n622), .A2(n359), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n623), .B(G146), .ZN(G48) );
  NAND2_X1 U697 ( .A1(n626), .A2(n359), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n624), .B(G113), .ZN(G15) );
  NAND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n627), .B(G116), .ZN(G18) );
  NAND2_X1 U701 ( .A1(n632), .A2(n474), .ZN(n669) );
  NOR2_X1 U702 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U703 ( .A(KEYINPUT49), .B(n635), .ZN(n641) );
  NAND2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U705 ( .A(n638), .B(KEYINPUT112), .ZN(n639) );
  XNOR2_X1 U706 ( .A(KEYINPUT50), .B(n639), .ZN(n640) );
  NAND2_X1 U707 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U708 ( .A1(n548), .A2(n642), .ZN(n643) );
  NOR2_X1 U709 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U710 ( .A(n645), .B(KEYINPUT113), .ZN(n646) );
  XNOR2_X1 U711 ( .A(KEYINPUT51), .B(n646), .ZN(n647) );
  NOR2_X1 U712 ( .A1(n664), .A2(n647), .ZN(n659) );
  NOR2_X1 U713 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U714 ( .A(n650), .B(KEYINPUT114), .ZN(n651) );
  NOR2_X1 U715 ( .A1(n652), .A2(n651), .ZN(n655) );
  NOR2_X1 U716 ( .A1(n362), .A2(n653), .ZN(n654) );
  NOR2_X1 U717 ( .A1(n655), .A2(n654), .ZN(n657) );
  NOR2_X1 U718 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U719 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U720 ( .A(n660), .B(KEYINPUT52), .ZN(n661) );
  NOR2_X1 U721 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U722 ( .A(KEYINPUT115), .B(n663), .Z(n666) );
  NOR2_X1 U723 ( .A1(n656), .A2(n664), .ZN(n665) );
  NOR2_X1 U724 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U725 ( .A(KEYINPUT116), .B(n667), .Z(n668) );
  NAND2_X1 U726 ( .A1(n684), .A2(G210), .ZN(n672) );
  XNOR2_X1 U727 ( .A(KEYINPUT80), .B(KEYINPUT56), .ZN(n674) );
  NAND2_X1 U728 ( .A1(n684), .A2(G475), .ZN(n677) );
  XOR2_X1 U729 ( .A(KEYINPUT65), .B(KEYINPUT60), .Z(n679) );
  XNOR2_X1 U730 ( .A(n680), .B(KEYINPUT120), .ZN(n682) );
  NAND2_X1 U731 ( .A1(G478), .A2(n684), .ZN(n681) );
  XNOR2_X1 U732 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U733 ( .A1(n688), .A2(n683), .ZN(G63) );
  NAND2_X1 U734 ( .A1(G217), .A2(n684), .ZN(n685) );
  XNOR2_X1 U735 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U736 ( .A1(n688), .A2(n687), .ZN(G66) );
  XNOR2_X1 U737 ( .A(n689), .B(G101), .ZN(n691) );
  NOR2_X1 U738 ( .A1(n474), .A2(G898), .ZN(n690) );
  NOR2_X1 U739 ( .A1(n691), .A2(n690), .ZN(n700) );
  NAND2_X1 U740 ( .A1(n692), .A2(n474), .ZN(n693) );
  XNOR2_X1 U741 ( .A(n693), .B(KEYINPUT122), .ZN(n698) );
  XOR2_X1 U742 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n695) );
  NAND2_X1 U743 ( .A1(G224), .A2(G953), .ZN(n694) );
  XNOR2_X1 U744 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U745 ( .A1(n696), .A2(G898), .ZN(n697) );
  NAND2_X1 U746 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U747 ( .A(n700), .B(n699), .ZN(G69) );
  XNOR2_X1 U748 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n702) );
  XNOR2_X1 U749 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U750 ( .A(n704), .B(n703), .ZN(n708) );
  XOR2_X1 U751 ( .A(n708), .B(n705), .Z(n706) );
  NOR2_X1 U752 ( .A1(G953), .A2(n706), .ZN(n707) );
  XNOR2_X1 U753 ( .A(KEYINPUT125), .B(n707), .ZN(n713) );
  XNOR2_X1 U754 ( .A(n708), .B(G227), .ZN(n709) );
  XNOR2_X1 U755 ( .A(n709), .B(KEYINPUT126), .ZN(n710) );
  NAND2_X1 U756 ( .A1(n710), .A2(G900), .ZN(n711) );
  NAND2_X1 U757 ( .A1(n711), .A2(G953), .ZN(n712) );
  NAND2_X1 U758 ( .A1(n713), .A2(n712), .ZN(G72) );
  XOR2_X1 U759 ( .A(G134), .B(n714), .Z(G36) );
  XOR2_X1 U760 ( .A(n715), .B(G122), .Z(G24) );
  XNOR2_X1 U761 ( .A(G143), .B(n716), .ZN(n717) );
  XNOR2_X1 U762 ( .A(n717), .B(KEYINPUT110), .ZN(G45) );
  XNOR2_X1 U763 ( .A(G119), .B(n718), .ZN(G21) );
  XNOR2_X1 U764 ( .A(n719), .B(KEYINPUT37), .ZN(n720) );
  XNOR2_X1 U765 ( .A(n720), .B(KEYINPUT111), .ZN(n721) );
  XNOR2_X1 U766 ( .A(G125), .B(n721), .ZN(G27) );
  XNOR2_X1 U767 ( .A(G140), .B(n722), .ZN(G42) );
  XNOR2_X1 U768 ( .A(G131), .B(n723), .ZN(G33) );
  XOR2_X1 U769 ( .A(G137), .B(n724), .Z(n725) );
  XNOR2_X1 U770 ( .A(KEYINPUT127), .B(n725), .ZN(G39) );
endmodule

