//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT67), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n465), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  AOI211_X1 g051(.A(new_n476), .B(new_n462), .C1(new_n472), .C2(new_n473), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n467), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n462), .ZN(new_n481));
  INV_X1    g056(.A(G137), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR3_X1   g058(.A1(new_n475), .A2(new_n477), .A3(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n463), .A2(new_n464), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n462), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  MUX2_X1   g064(.A(G100), .B(G112), .S(G2105), .Z(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2104), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(G162));
  NAND3_X1  g067(.A1(new_n480), .A2(KEYINPUT4), .A3(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n480), .B2(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT4), .B1(new_n498), .B2(new_n462), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n465), .A2(new_n471), .A3(G138), .A4(new_n462), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G88), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n508), .A2(new_n511), .ZN(G166));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT7), .ZN(new_n514));
  XOR2_X1   g089(.A(KEYINPUT69), .B(G51), .Z(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n506), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n503), .A2(G89), .ZN(new_n520));
  NAND2_X1  g095(.A1(G63), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G168));
  INV_X1    g098(.A(G90), .ZN(new_n524));
  INV_X1    g099(.A(G52), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n504), .A2(new_n524), .B1(new_n506), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n510), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(G171));
  AOI22_X1  g104(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(new_n510), .ZN(new_n531));
  AND2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n519), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(G81), .A2(new_n535), .B1(new_n537), .B2(G43), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n531), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n504), .A2(new_n541), .B1(new_n506), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n530), .A2(new_n510), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT70), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n537), .A2(new_n554), .A3(G53), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n506), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n535), .A2(G91), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n510), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(G299));
  NAND2_X1  g137(.A1(G171), .A2(KEYINPUT71), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n564), .B1(new_n526), .B2(new_n528), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  OR2_X1    g143(.A1(new_n508), .A2(new_n511), .ZN(G303));
  NAND2_X1  g144(.A1(new_n535), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n537), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND3_X1  g148(.A1(new_n502), .A2(new_n503), .A3(G86), .ZN(new_n574));
  AND2_X1   g149(.A1(G48), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n575), .B1(new_n532), .B2(new_n533), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT73), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n503), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n574), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n510), .ZN(new_n583));
  OAI21_X1  g158(.A(G61), .B1(new_n517), .B2(new_n518), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n586), .A2(KEYINPUT72), .A3(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n580), .A2(new_n583), .A3(new_n587), .ZN(G305));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n504), .A2(new_n589), .B1(new_n506), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n510), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  AND3_X1   g170(.A1(new_n502), .A2(new_n503), .A3(G92), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n519), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(new_n537), .B2(G54), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n566), .B2(new_n604), .ZN(G284));
  OAI21_X1  g181(.A(new_n605), .B1(new_n566), .B2(new_n604), .ZN(G321));
  MUX2_X1   g182(.A(G286), .B(G299), .S(new_n604), .Z(G297));
  MUX2_X1   g183(.A(G286), .B(G299), .S(new_n604), .Z(G280));
  INV_X1    g184(.A(G860), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n603), .B1(G559), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT75), .ZN(G148));
  OAI21_X1  g187(.A(G868), .B1(new_n603), .B2(G559), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n547), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(KEYINPUT76), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT76), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g192(.A1(new_n465), .A2(new_n471), .A3(new_n478), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT13), .Z(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT78), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(G2100), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT77), .ZN(new_n624));
  MUX2_X1   g199(.A(G99), .B(G111), .S(G2105), .Z(new_n625));
  AOI22_X1  g200(.A1(new_n488), .A2(G123), .B1(G2104), .B2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G135), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n481), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT79), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n622), .A2(new_n624), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT80), .Z(G156));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT15), .B(G2435), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2427), .ZN(new_n637));
  INV_X1    g212(.A(G2430), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n640), .A2(new_n646), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  INV_X1    g229(.A(new_n650), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(new_n652), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n650), .A2(new_n652), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n651), .B1(new_n660), .B2(KEYINPUT17), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n654), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n630), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(G227));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n667), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT81), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n673), .A2(new_n674), .A3(new_n670), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n673), .B1(new_n674), .B2(new_n670), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(G229));
  NOR2_X1   g260(.A1(G5), .A2(G16), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G171), .B2(G16), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT94), .Z(new_n688));
  INV_X1    g263(.A(G1961), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(G27), .A2(G29), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G164), .B2(G29), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n690), .B1(G2078), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G29), .A2(G35), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G162), .B2(G29), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT29), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(G2090), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n692), .A2(G2078), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n696), .B2(G2090), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G20), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT23), .ZN(new_n702));
  INV_X1    g277(.A(G299), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n700), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1956), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n689), .B2(new_n688), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n693), .A2(new_n697), .A3(new_n699), .A4(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G21), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G168), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT91), .ZN(new_n710));
  INV_X1    g285(.A(G1966), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT93), .Z(new_n713));
  NAND2_X1  g288(.A1(G160), .A2(G29), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  AND2_X1   g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  NOR2_X1   g291(.A1(KEYINPUT24), .A2(G34), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G2084), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n707), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n598), .A2(new_n602), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G4), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1348), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n715), .A2(G32), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT89), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT26), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n488), .A2(G129), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n486), .A2(G141), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n478), .A2(G105), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n729), .B1(new_n737), .B2(new_n715), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n728), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n715), .A2(G26), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n486), .A2(G140), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n488), .A2(G128), .ZN(new_n745));
  MUX2_X1   g320(.A(G104), .B(G116), .S(G2105), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G2104), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n749), .B2(new_n715), .ZN(new_n750));
  INV_X1    g325(.A(G2067), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n710), .A2(new_n711), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT31), .B(G11), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT92), .B(G28), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT30), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n754), .B1(new_n756), .B2(new_n715), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n629), .B2(new_n715), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n726), .B2(new_n727), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n741), .A2(new_n752), .A3(new_n753), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n700), .A2(G19), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n547), .B2(new_n700), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1341), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n723), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n719), .A2(new_n720), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n738), .A2(new_n740), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n465), .A2(new_n471), .A3(G127), .ZN(new_n769));
  NAND2_X1  g344(.A1(G115), .A2(G2104), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n462), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT87), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n773), .A2(KEYINPUT87), .A3(G2105), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n478), .A2(G103), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT86), .B(KEYINPUT25), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G139), .B2(new_n486), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n772), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G29), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n715), .A2(G33), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n782), .B2(G2072), .ZN(new_n784));
  AND3_X1   g359(.A1(new_n782), .A2(new_n783), .A3(G2072), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n768), .B1(G2072), .B2(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n765), .A2(new_n788), .A3(KEYINPUT95), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n723), .A2(new_n789), .A3(new_n764), .ZN(new_n792));
  INV_X1    g367(.A(new_n788), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G25), .A2(G29), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n486), .A2(G131), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n488), .A2(G119), .ZN(new_n797));
  MUX2_X1   g372(.A(G95), .B(G107), .S(G2105), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G2104), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT35), .B(G1991), .Z(new_n803));
  XOR2_X1   g378(.A(new_n802), .B(new_n803), .Z(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G24), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n594), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1986), .ZN(new_n807));
  MUX2_X1   g382(.A(G6), .B(G305), .S(G16), .Z(new_n808));
  XOR2_X1   g383(.A(KEYINPUT32), .B(G1981), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G16), .A2(G22), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G166), .B2(G16), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT83), .B(G1971), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n700), .A2(G23), .ZN(new_n815));
  INV_X1    g390(.A(G288), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n700), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT33), .B(G1976), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT82), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n810), .A2(new_n814), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT34), .ZN(new_n822));
  AOI211_X1 g397(.A(new_n804), .B(new_n807), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT84), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(KEYINPUT84), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT85), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n827), .A2(new_n828), .A3(KEYINPUT36), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n823), .B(new_n830), .C1(new_n825), .C2(new_n826), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n790), .A2(new_n794), .B1(new_n829), .B2(new_n831), .ZN(G311));
  NAND2_X1  g407(.A1(new_n790), .A2(new_n794), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n829), .A2(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(G150));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n504), .A2(new_n836), .B1(new_n506), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(new_n510), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n610), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n724), .A2(G559), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n838), .A2(new_n840), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n546), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n841), .A2(new_n531), .A3(new_n538), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(KEYINPUT97), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n841), .B1(new_n540), .B2(new_n545), .ZN(new_n852));
  NOR4_X1   g427(.A1(new_n544), .A2(new_n543), .A3(new_n838), .A4(new_n840), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n846), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n846), .A2(new_n855), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT39), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n858), .B2(KEYINPUT98), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(KEYINPUT98), .B2(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT39), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT99), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n843), .B1(new_n860), .B2(new_n862), .ZN(G145));
  XNOR2_X1  g438(.A(new_n619), .B(new_n800), .ZN(new_n864));
  MUX2_X1   g439(.A(G106), .B(G118), .S(G2105), .Z(new_n865));
  AOI22_X1  g440(.A1(new_n488), .A2(G130), .B1(G2104), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G142), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n481), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT101), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n864), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(G164), .B(new_n748), .ZN(new_n871));
  INV_X1    g446(.A(new_n737), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(G126), .B1(new_n463), .B2(new_n464), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n462), .B1(new_n874), .B2(new_n496), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT4), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n500), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(KEYINPUT4), .A2(G138), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n485), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n494), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n462), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n748), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n737), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n873), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n779), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n779), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n779), .A2(new_n886), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n873), .A2(new_n888), .A3(new_n884), .A4(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n887), .A2(KEYINPUT103), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT103), .B1(new_n887), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n870), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(G160), .B(G162), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n629), .ZN(new_n897));
  INV_X1    g472(.A(new_n870), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n887), .A2(new_n890), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g475(.A(KEYINPUT104), .B(new_n870), .C1(new_n891), .C2(new_n892), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n895), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT102), .B1(new_n899), .B2(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(new_n898), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n887), .A2(new_n905), .A3(new_n870), .A4(new_n890), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G37), .B1(new_n907), .B2(new_n897), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g485(.A1(new_n847), .A2(new_n604), .ZN(new_n911));
  XNOR2_X1  g486(.A(G305), .B(G166), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n594), .B(G288), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(KEYINPUT107), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n912), .A2(new_n913), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT108), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n603), .A2(G559), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n850), .A2(new_n927), .A3(new_n854), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n850), .B2(new_n854), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n724), .B2(G299), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n603), .A3(KEYINPUT105), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n724), .A2(G299), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(KEYINPUT41), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n932), .A2(new_n939), .A3(new_n933), .A4(new_n934), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n938), .B(new_n940), .C1(new_n928), .C2(new_n929), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n936), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n941), .A2(new_n937), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT109), .B1(new_n926), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n921), .A2(new_n925), .ZN(new_n947));
  OAI221_X1 g522(.A(new_n946), .B1(new_n942), .B2(new_n943), .C1(new_n947), .C2(new_n924), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n926), .A2(new_n944), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n911), .B1(new_n950), .B2(new_n604), .ZN(G295));
  OAI21_X1  g526(.A(new_n911), .B1(new_n950), .B2(new_n604), .ZN(G331));
  NAND3_X1  g527(.A1(new_n563), .A2(G168), .A3(new_n565), .ZN(new_n953));
  NAND2_X1  g528(.A1(G286), .A2(G171), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n850), .A3(new_n854), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n955), .B1(new_n850), .B2(new_n854), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n938), .B(new_n940), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n954), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n855), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n935), .A3(new_n956), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n921), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  INV_X1    g540(.A(G37), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n959), .A2(new_n920), .A3(new_n962), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT110), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n967), .A2(new_n966), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n965), .A4(new_n964), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n966), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n920), .B1(new_n959), .B2(new_n962), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(KEYINPUT44), .A3(new_n968), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(G397));
  NAND2_X1  g555(.A1(new_n872), .A2(G1996), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n737), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n748), .B(new_n751), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n472), .A2(new_n473), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n476), .B1(new_n986), .B2(new_n462), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n483), .B1(new_n474), .B2(KEYINPUT68), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(G40), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(G164), .B2(G1384), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n985), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT112), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n800), .B(new_n803), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n992), .ZN(new_n998));
  NAND2_X1  g573(.A1(G290), .A2(G1986), .ZN(new_n999));
  OR2_X1    g574(.A1(G290), .A2(G1986), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT111), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(G160), .A2(new_n991), .A3(G40), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1971), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n987), .A2(new_n988), .A3(G40), .ZN(new_n1009));
  INV_X1    g584(.A(G2090), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n882), .A2(new_n1004), .A3(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(G8), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n877), .B2(new_n881), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1022), .A2(new_n987), .A3(new_n988), .A4(G40), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n816), .A2(G1976), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(G8), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT114), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1028), .A3(KEYINPUT52), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1023), .A2(G8), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n580), .A2(new_n583), .A3(new_n587), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT115), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT72), .B1(new_n586), .B2(G651), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n581), .B(new_n510), .C1(new_n584), .C2(new_n585), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1032), .A4(new_n580), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n580), .B1(new_n510), .B2(new_n582), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G1981), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1031), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AND4_X1   g620(.A1(KEYINPUT116), .A2(new_n1040), .A3(KEYINPUT49), .A4(new_n1042), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1034), .A2(new_n1039), .B1(G1981), .B2(new_n1041), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT116), .B1(new_n1047), .B2(KEYINPUT49), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1045), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n816), .A2(G1976), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n1025), .A2(KEYINPUT52), .A3(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1021), .A2(new_n1030), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n689), .B1(new_n1053), .B2(new_n989), .ZN(new_n1054));
  NOR4_X1   g629(.A1(G164), .A2(KEYINPUT121), .A3(new_n990), .A4(G1384), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n1022), .B2(KEYINPUT45), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1009), .B(new_n991), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G2078), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT53), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1054), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1009), .A2(new_n1059), .A3(new_n1005), .A4(new_n991), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(KEYINPUT124), .A3(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1012), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(G164), .B2(G1384), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n1071));
  AND4_X1   g646(.A1(KEYINPUT120), .A2(new_n882), .A3(new_n1071), .A4(new_n1004), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT120), .B1(new_n1022), .B2(new_n1071), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1009), .B(new_n1070), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1008), .B1(new_n1074), .B2(G2090), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1020), .B1(new_n1075), .B2(G8), .ZN(new_n1076));
  NOR4_X1   g651(.A1(new_n1052), .A2(new_n1068), .A3(new_n1076), .A4(G301), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1058), .A2(new_n711), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1009), .A2(new_n720), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(G168), .ZN(new_n1080));
  AOI21_X1  g655(.A(G168), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  OAI211_X1 g657(.A(G8), .B(new_n1080), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1005), .A2(KEYINPUT121), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1022), .A2(new_n1056), .A3(KEYINPUT45), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT45), .B1(new_n882), .B2(new_n1004), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n989), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1966), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1079), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1089), .A2(new_n1090), .A3(G286), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT51), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1083), .A2(KEYINPUT62), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT62), .B1(new_n1083), .B2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1077), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1031), .B(KEYINPUT117), .ZN(new_n1098));
  NOR2_X1   g673(.A1(G288), .A2(G1976), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT118), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1049), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1101), .B2(new_n1040), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n1092), .B(new_n1019), .C1(new_n1008), .C2(new_n1014), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n1103), .A2(new_n1030), .A3(new_n1051), .A4(new_n1049), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1097), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1103), .A2(new_n1030), .A3(new_n1051), .A4(new_n1049), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1049), .A2(new_n1100), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1106), .B(KEYINPUT119), .C1(new_n1107), .C2(new_n1098), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(G8), .B(G168), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1052), .A2(new_n1110), .A3(new_n1076), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1110), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1092), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1112), .B(KEYINPUT63), .C1(new_n1113), .C2(new_n1020), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1111), .A2(KEYINPUT63), .B1(new_n1052), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1096), .A2(new_n1109), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1009), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1117));
  AOI211_X1 g692(.A(new_n990), .B(G1384), .C1(new_n877), .C2(new_n881), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1087), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G40), .ZN(new_n1120));
  NOR4_X1   g695(.A1(new_n474), .A2(new_n483), .A3(new_n1120), .A4(new_n1060), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1117), .A2(new_n689), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1067), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT124), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1124));
  OAI211_X1 g699(.A(G301), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1068), .B2(G301), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G171), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1068), .A2(G301), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(KEYINPUT54), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1052), .A2(new_n1076), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1083), .A2(new_n1093), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1128), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1956), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1137));
  NAND3_X1  g712(.A1(G160), .A2(new_n1070), .A3(G40), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n989), .A2(new_n1087), .A3(new_n1118), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT56), .B(G2072), .Z(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G299), .B(KEYINPUT57), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1139), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT122), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1074), .A2(new_n1136), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(new_n1149), .A3(new_n1145), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n727), .B1(new_n1053), .B2(new_n989), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1023), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n751), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n603), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n882), .A2(new_n1071), .A3(new_n1004), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1022), .A2(KEYINPUT120), .A3(new_n1071), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1022), .A2(new_n1012), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n989), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(G1956), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NOR4_X1   g738(.A1(new_n989), .A2(new_n1087), .A3(new_n1118), .A4(new_n1141), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1144), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1147), .A2(new_n1150), .B1(new_n1155), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1149), .B1(new_n1148), .B2(new_n1145), .ZN(new_n1167));
  NOR4_X1   g742(.A1(new_n1163), .A2(new_n1164), .A3(KEYINPUT122), .A4(new_n1144), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(KEYINPUT58), .B(G1341), .Z(new_n1172));
  AOI22_X1  g747(.A1(new_n1140), .A2(new_n982), .B1(new_n1023), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT59), .B1(new_n1173), .B2(new_n546), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1006), .A2(G1996), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1023), .A2(new_n1172), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1175), .B(new_n547), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1165), .A2(new_n1146), .A3(KEYINPUT61), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1117), .A2(new_n727), .B1(new_n1152), .B2(new_n751), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n603), .B(KEYINPUT60), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1154), .A2(KEYINPUT60), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1179), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1166), .B1(new_n1171), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1135), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1003), .B1(new_n1116), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n997), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT127), .B1(new_n994), .B2(new_n996), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n998), .A2(new_n1000), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT48), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT46), .ZN(new_n1194));
  OAI22_X1  g769(.A1(new_n998), .A2(G1996), .B1(KEYINPUT126), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1195), .B1(new_n1196), .B2(KEYINPUT46), .ZN(new_n1197));
  OAI211_X1 g772(.A(KEYINPUT126), .B(new_n1194), .C1(new_n998), .C2(G1996), .ZN(new_n1198));
  INV_X1    g773(.A(new_n984), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n992), .B1(new_n1199), .B2(new_n872), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT47), .Z(new_n1202));
  NAND2_X1  g777(.A1(new_n801), .A2(new_n803), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT125), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n994), .A2(new_n1204), .B1(new_n751), .B2(new_n749), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1205), .A2(new_n998), .ZN(new_n1206));
  NOR3_X1   g781(.A1(new_n1193), .A2(new_n1202), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1187), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g783(.A1(new_n460), .A2(G229), .A3(G227), .A4(G401), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n1210), .B1(new_n902), .B2(new_n908), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n976), .A2(new_n1211), .ZN(G225));
  INV_X1    g786(.A(G225), .ZN(G308));
endmodule


