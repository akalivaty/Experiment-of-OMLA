//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT64), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  OR4_X1    g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(G101), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI22_X1  g045(.A1(new_n464), .A2(new_n465), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n469), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n467), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n462), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n477), .A2(G124), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n470), .A2(KEYINPUT69), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n470), .A2(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT70), .Z(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G138), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n476), .B2(new_n492), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n493), .A2(G2105), .B1(G102), .B2(new_n463), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT71), .B1(new_n499), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(new_n497), .A3(KEYINPUT5), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n506), .A2(new_n510), .ZN(G166));
  NAND2_X1  g086(.A1(new_n503), .A2(new_n508), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n514));
  AND3_X1   g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n513), .A2(G89), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT72), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n519), .A2(G651), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n522), .A2(G51), .A3(G543), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n527), .B2(new_n528), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n518), .B1(new_n531), .B2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND3_X1  g109(.A1(new_n522), .A2(G543), .A3(new_n526), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n512), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n503), .A2(G64), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n505), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND4_X1  g117(.A1(new_n522), .A2(G43), .A3(G543), .A4(new_n526), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n500), .A2(new_n502), .ZN(new_n544));
  INV_X1    g119(.A(new_n498), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n544), .A2(G81), .A3(new_n545), .A4(new_n508), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n501), .B1(KEYINPUT5), .B2(new_n497), .ZN(new_n548));
  NOR3_X1   g123(.A1(new_n499), .A2(KEYINPUT71), .A3(G543), .ZN(new_n549));
  OAI211_X1 g124(.A(G56), .B(new_n545), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n505), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n522), .A2(G53), .A3(G543), .A4(new_n526), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n503), .A2(G91), .A3(new_n508), .ZN(new_n563));
  INV_X1    g138(.A(G78), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n497), .ZN(new_n565));
  AND2_X1   g140(.A1(KEYINPUT75), .A2(G65), .ZN(new_n566));
  NOR2_X1   g141(.A1(KEYINPUT75), .A2(G65), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n565), .B1(new_n503), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n563), .B1(new_n569), .B2(new_n505), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n560), .B1(new_n562), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n525), .B1(new_n523), .B2(new_n524), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n575), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n561), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g154(.A1(new_n579), .A2(KEYINPUT76), .A3(new_n570), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  OR2_X1    g158(.A1(new_n506), .A2(new_n510), .ZN(G303));
  OAI21_X1  g159(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI221_X1 g162(.A(new_n585), .B1(new_n512), .B2(new_n586), .C1(new_n587), .C2(new_n535), .ZN(G288));
  AOI22_X1  g163(.A1(new_n503), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n505), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n503), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n509), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT77), .ZN(G305));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n535), .A2(new_n595), .B1(new_n512), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n505), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n535), .B(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G54), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n513), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n512), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n503), .A2(G66), .ZN(new_n609));
  INV_X1    g184(.A(G79), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n497), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n605), .A2(new_n608), .B1(G651), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n602), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n602), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  MUX2_X1   g192(.A(G286), .B(G299), .S(new_n617), .Z(G297));
  MUX2_X1   g193(.A(G286), .B(G299), .S(new_n617), .Z(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n614), .B1(new_n620), .B2(G860), .ZN(G148));
  NOR2_X1   g196(.A1(new_n613), .A2(G559), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT79), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g201(.A1(new_n464), .A2(new_n476), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n477), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n632), .B1(new_n633), .B2(new_n634), .C1(new_n484), .C2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n631), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2435), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2438), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT81), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n650), .B(new_n651), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(KEYINPUT82), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n658), .A3(new_n666), .ZN(new_n667));
  OAI221_X1 g242(.A(new_n661), .B1(new_n662), .B2(new_n663), .C1(new_n665), .C2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2096), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2100), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n673), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  AOI22_X1  g254(.A1(new_n677), .A2(KEYINPUT20), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n681), .A2(new_n673), .A3(new_n676), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n680), .B(new_n682), .C1(KEYINPUT20), .C2(new_n677), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G229));
  NAND2_X1  g264(.A1(new_n477), .A2(G119), .ZN(new_n690));
  OR2_X1    g265(.A1(G95), .A2(G2105), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n462), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI221_X1 g268(.A(new_n693), .B1(new_n692), .B2(new_n691), .C1(G107), .C2(new_n467), .ZN(new_n694));
  INV_X1    g269(.A(G131), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n690), .B(new_n694), .C1(new_n484), .C2(new_n695), .ZN(new_n696));
  MUX2_X1   g271(.A(G25), .B(new_n696), .S(G29), .Z(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT35), .B(G1991), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n600), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n700), .B2(G24), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n699), .B1(G1986), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G6), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G16), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G305), .B2(G16), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n710), .A2(new_n711), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n707), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n714), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n716), .A2(new_n706), .A3(new_n712), .ZN(new_n717));
  MUX2_X1   g292(.A(G23), .B(G288), .S(G16), .Z(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT33), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT33), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n719), .A2(G1976), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n700), .A2(G22), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G166), .B2(new_n700), .ZN(new_n723));
  MUX2_X1   g298(.A(new_n722), .B(new_n723), .S(KEYINPUT85), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G1971), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(G1976), .B1(new_n719), .B2(new_n720), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n724), .A2(G1971), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n715), .A2(new_n717), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n705), .B1(new_n730), .B2(KEYINPUT34), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n717), .A2(new_n728), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT34), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n732), .A2(new_n733), .A3(new_n729), .A4(new_n715), .ZN(new_n734));
  INV_X1    g309(.A(G1986), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n702), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n731), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(KEYINPUT36), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n731), .A2(new_n734), .A3(new_n739), .A4(new_n736), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n700), .A2(KEYINPUT23), .A3(G20), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n743));
  INV_X1    g318(.A(G20), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G16), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n742), .B(new_n745), .C1(new_n581), .C2(new_n700), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1956), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n748), .ZN(new_n750));
  MUX2_X1   g325(.A(new_n749), .B(new_n750), .S(KEYINPUT94), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT29), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n747), .B1(new_n752), .B2(G2090), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G2090), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n614), .A2(new_n700), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G4), .B2(new_n700), .ZN(new_n756));
  INV_X1    g331(.A(G1348), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  NAND2_X1  g334(.A1(G168), .A2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G16), .B2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G5), .A2(G16), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G171), .B2(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n748), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n748), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n764), .A2(G1961), .B1(new_n766), .B2(G2078), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n767), .B1(G1961), .B2(new_n764), .C1(new_n756), .C2(new_n757), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n766), .A2(G2078), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n762), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G29), .A2(G32), .ZN(new_n771));
  INV_X1    g346(.A(new_n464), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n772), .A2(G105), .B1(G129), .B2(new_n477), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT26), .Z(new_n775));
  NAND3_X1  g350(.A1(new_n482), .A2(G141), .A3(new_n483), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT87), .B1(G29), .B2(G33), .ZN(new_n782));
  OR3_X1    g357(.A1(KEYINPUT87), .A2(G29), .A3(G33), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n482), .A2(G139), .A3(new_n483), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n463), .A2(G103), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n784), .A2(KEYINPUT89), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT89), .B1(new_n784), .B2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  INV_X1    g365(.A(G127), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n476), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT90), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n788), .A2(new_n789), .B1(new_n467), .B2(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n782), .B(new_n783), .C1(new_n794), .C2(new_n748), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2072), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n748), .A2(G26), .ZN(new_n797));
  OR2_X1    g372(.A1(G104), .A2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT86), .Z(new_n800));
  NAND3_X1  g375(.A1(new_n482), .A2(G140), .A3(new_n483), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n477), .A2(G128), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n748), .ZN(new_n804));
  MUX2_X1   g379(.A(new_n797), .B(new_n804), .S(KEYINPUT28), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2067), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n700), .A2(G19), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n553), .B2(new_n700), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1341), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G34), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(G29), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G160), .B2(G29), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(G2084), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT30), .B(G28), .Z(new_n815));
  MUX2_X1   g390(.A(new_n815), .B(new_n636), .S(G29), .Z(new_n816));
  XOR2_X1   g391(.A(KEYINPUT31), .B(G11), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT92), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n813), .A2(G2084), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n814), .A2(new_n816), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n806), .A2(new_n809), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n770), .A2(new_n781), .A3(new_n796), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n754), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n761), .A2(new_n759), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT93), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n741), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(G311));
  NAND2_X1  g402(.A1(new_n826), .A2(KEYINPUT95), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n741), .A2(new_n823), .A3(new_n829), .A4(new_n825), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(G150));
  NAND4_X1  g406(.A1(new_n522), .A2(G55), .A3(G543), .A4(new_n526), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n503), .A2(G93), .A3(new_n508), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n505), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n614), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT39), .ZN(new_n840));
  INV_X1    g415(.A(new_n551), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n503), .B2(G56), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n543), .B(new_n546), .C1(new_n842), .C2(new_n505), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n503), .A2(G67), .ZN(new_n844));
  AND2_X1   g419(.A1(G80), .A2(G543), .ZN(new_n845));
  OAI21_X1  g420(.A(G651), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n832), .A2(new_n833), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n553), .A2(new_n835), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n851));
  XOR2_X1   g426(.A(new_n850), .B(new_n851), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n840), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n838), .B1(new_n853), .B2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT98), .Z(G145));
  INV_X1    g430(.A(new_n629), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n803), .A2(new_n495), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G164), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n778), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n857), .A2(new_n777), .A3(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n794), .A2(KEYINPUT99), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n477), .A2(G130), .ZN(new_n867));
  NOR2_X1   g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(new_n467), .B2(G118), .ZN(new_n869));
  INV_X1    g444(.A(G142), .ZN(new_n870));
  OAI221_X1 g445(.A(new_n867), .B1(new_n868), .B2(new_n869), .C1(new_n484), .C2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(new_n696), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n794), .A2(KEYINPUT99), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n861), .A2(new_n864), .A3(new_n873), .A4(new_n862), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n866), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n872), .B1(new_n866), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n856), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n629), .A3(new_n875), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT101), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G162), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT101), .A4(new_n487), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n636), .B(G160), .Z(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(KEYINPUT100), .B(G37), .Z(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g467(.A1(new_n835), .A2(new_n617), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n623), .B(new_n850), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n613), .B(KEYINPUT102), .C1(new_n572), .C2(new_n580), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT102), .B1(new_n572), .B2(new_n580), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n562), .A2(new_n560), .A3(new_n571), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT76), .B1(new_n579), .B2(new_n570), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n614), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n894), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n895), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n905), .A3(new_n895), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n894), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n902), .B1(new_n909), .B2(KEYINPUT103), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(KEYINPUT103), .B2(new_n902), .ZN(new_n911));
  XNOR2_X1  g486(.A(G303), .B(G288), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G305), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n912), .A2(G305), .ZN(new_n915));
  OAI21_X1  g490(.A(G290), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n915), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n600), .A3(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT42), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n911), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n893), .B1(new_n921), .B2(new_n617), .ZN(G295));
  OAI21_X1  g497(.A(new_n893), .B1(new_n921), .B2(new_n617), .ZN(G331));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n553), .A2(new_n835), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n843), .A2(new_n846), .A3(new_n847), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT105), .B1(new_n538), .B2(new_n541), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n926), .B2(new_n927), .ZN(new_n930));
  INV_X1    g505(.A(new_n541), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n513), .A2(G90), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n573), .A2(new_n574), .A3(new_n497), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G52), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n532), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n530), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n938), .A3(new_n518), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n929), .A2(new_n930), .A3(new_n939), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n538), .A2(new_n541), .A3(KEYINPUT105), .ZN(new_n941));
  NOR2_X1   g516(.A1(G286), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n928), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n848), .B2(new_n849), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n925), .B1(new_n947), .B2(new_n903), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n939), .B1(new_n929), .B2(new_n930), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n942), .A3(new_n945), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(KEYINPUT106), .A3(new_n895), .A4(new_n901), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n906), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n905), .B1(new_n901), .B2(new_n895), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n947), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n919), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n924), .B1(new_n957), .B2(G37), .ZN(new_n958));
  INV_X1    g533(.A(G37), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n907), .A2(new_n947), .B1(new_n948), .B2(new_n952), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT107), .B(new_n959), .C1(new_n960), .C2(new_n919), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n919), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n955), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n947), .B(new_n968), .C1(new_n907), .C2(new_n967), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n951), .A2(new_n895), .A3(new_n901), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n919), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n888), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n964), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n962), .A3(new_n974), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n965), .A2(new_n966), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n972), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n889), .A3(new_n962), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n958), .A2(new_n961), .A3(new_n962), .A4(new_n974), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n966), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT109), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n980), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n973), .B2(new_n962), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT44), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n965), .A2(new_n975), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n986), .B(new_n987), .C1(KEYINPUT44), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n989), .ZN(G397));
  AOI21_X1  g565(.A(G1384), .B1(new_n490), .B2(new_n494), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G40), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n471), .A2(new_n994), .A3(new_n474), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1996), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n998), .A2(new_n999), .A3(new_n778), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  INV_X1    g578(.A(G2067), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n858), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G1996), .B2(new_n777), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n1002), .B(new_n1003), .C1(new_n997), .C2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n696), .B(new_n698), .Z(new_n1008));
  OAI21_X1  g583(.A(new_n1007), .B1(new_n998), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n600), .B(new_n735), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n997), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n995), .B1(new_n991), .B2(KEYINPUT45), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n759), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n495), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(G2084), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n991), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1019), .A2(new_n1020), .A3(new_n995), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1012), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(KEYINPUT123), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT123), .ZN(new_n1026));
  AOI211_X1 g601(.A(new_n1026), .B(new_n1012), .C1(new_n1016), .C2(new_n1023), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G168), .A2(new_n1012), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1025), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1029), .B1(new_n1036), .B2(KEYINPUT51), .ZN(new_n1037));
  OAI22_X1  g612(.A1(new_n1032), .A2(new_n1033), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1028), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT62), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n1028), .B(new_n1034), .C1(new_n1024), .C2(new_n1033), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1036), .A2(new_n1026), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1031), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1024), .A2(KEYINPUT123), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1045), .B2(KEYINPUT51), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT62), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1039), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1040), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT127), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n996), .A2(new_n1018), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(new_n1012), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G288), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT52), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n593), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(G1981), .B1(new_n590), .B2(new_n592), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT49), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(KEYINPUT49), .A3(new_n1060), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1053), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1053), .B(new_n1066), .C1(new_n1055), .C2(G288), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1057), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(G166), .B2(new_n1012), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT55), .B(G8), .C1(new_n506), .C2(new_n510), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT112), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1075), .A3(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1013), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n991), .A2(KEYINPUT111), .A3(KEYINPUT45), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1015), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1019), .A2(new_n995), .A3(new_n1022), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1081), .A2(G1971), .B1(new_n1082), .B2(G2090), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1077), .A2(new_n1083), .A3(G8), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1077), .A2(new_n1083), .A3(KEYINPUT113), .A4(G8), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1068), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1019), .A2(new_n1089), .A3(new_n995), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n995), .B1(new_n991), .B2(new_n1021), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT116), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1092), .A3(new_n1022), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G2090), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1081), .A2(G1971), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1088), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  OR4_X1    g676(.A1(new_n1101), .A2(new_n1014), .A3(new_n1015), .A4(G2078), .ZN(new_n1102));
  INV_X1    g677(.A(G1961), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1082), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT125), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1015), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1101), .B1(new_n1109), .B2(G2078), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1102), .A2(new_n1111), .A3(new_n1104), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1106), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1050), .A2(new_n1051), .A3(new_n1100), .A4(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1100), .B(new_n1114), .C1(new_n1040), .C2(new_n1049), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT127), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n1068), .ZN(new_n1120));
  NOR2_X1   g695(.A1(G288), .A2(G1976), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1065), .A2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1059), .B(KEYINPUT114), .Z(new_n1124));
  AOI21_X1  g699(.A(new_n1054), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1126), .B(new_n1068), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1024), .A2(G168), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT117), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1083), .A2(G8), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1097), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1120), .B(new_n1125), .C1(new_n1132), .C2(KEYINPUT63), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT118), .B(G1956), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n1093), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1081), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT120), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n562), .A2(new_n571), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n570), .B2(KEYINPUT119), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1140), .B(new_n1142), .Z(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1082), .A2(new_n757), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1052), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1146), .B1(G2067), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1148), .A2(new_n614), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1135), .A2(new_n1143), .A3(new_n1137), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(KEYINPUT61), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n613), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT58), .B(G1341), .Z(new_n1156));
  NAND2_X1  g731(.A1(new_n1147), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1109), .B2(G1996), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n553), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1081), .A2(new_n999), .B1(new_n1147), .B2(new_n1156), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n553), .A2(new_n1159), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT59), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1155), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1135), .A2(new_n1143), .A3(new_n1137), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1143), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1148), .A2(new_n614), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT60), .B1(new_n1149), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1165), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1145), .B(new_n1151), .C1(new_n1154), .C2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(G171), .B(KEYINPUT54), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n1113), .A2(new_n1174), .ZN(new_n1175));
  OR4_X1    g750(.A1(new_n1101), .A2(new_n992), .A3(G2078), .A4(new_n474), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n994), .B1(new_n471), .B2(KEYINPUT126), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(KEYINPUT126), .B2(new_n471), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1174), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1181), .A2(new_n1104), .A3(new_n1110), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1175), .B(new_n1182), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1173), .A2(new_n1184), .B1(new_n1129), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1133), .B1(new_n1186), .B2(new_n1099), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1011), .B1(new_n1118), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n997), .A2(new_n735), .A3(new_n600), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT48), .Z(new_n1190));
  NOR2_X1   g765(.A1(new_n1009), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n696), .A2(new_n698), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1007), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n803), .A2(new_n1004), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n998), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OR3_X1    g770(.A1(new_n998), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1196));
  OAI21_X1  g771(.A(KEYINPUT46), .B1(new_n998), .B2(G1996), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1005), .A2(new_n778), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1196), .A2(new_n1197), .B1(new_n997), .B2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT47), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1191), .A2(new_n1195), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1188), .A2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g777(.A1(G229), .A2(new_n460), .ZN(new_n1204));
  NOR2_X1   g778(.A1(G401), .A2(G227), .ZN(new_n1205));
  NAND4_X1  g779(.A1(new_n891), .A2(new_n988), .A3(new_n1204), .A4(new_n1205), .ZN(G225));
  INV_X1    g780(.A(G225), .ZN(G308));
endmodule


