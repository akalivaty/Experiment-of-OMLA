

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U545 ( .A(n522), .B(n521), .ZN(n600) );
  XNOR2_X2 U546 ( .A(n754), .B(KEYINPUT98), .ZN(n760) );
  AND2_X2 U547 ( .A1(n753), .A2(n514), .ZN(n754) );
  AND2_X1 U548 ( .A1(n958), .A2(n818), .ZN(n805) );
  AND2_X2 U549 ( .A1(G2105), .A2(G2104), .ZN(n871) );
  NOR2_X1 U550 ( .A1(n770), .A2(n771), .ZN(n512) );
  OR2_X2 U551 ( .A1(n512), .A2(n513), .ZN(n821) );
  OR2_X1 U552 ( .A1(n805), .A2(n804), .ZN(n513) );
  XNOR2_X1 U553 ( .A(n519), .B(n518), .ZN(n601) );
  INV_X1 U554 ( .A(KEYINPUT17), .ZN(n518) );
  NOR2_X1 U555 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  BUF_X1 U556 ( .A(n714), .Z(n700) );
  BUF_X1 U557 ( .A(n601), .Z(n875) );
  NAND2_X1 U558 ( .A1(n601), .A2(G137), .ZN(n530) );
  NAND2_X1 U559 ( .A1(n752), .A2(n751), .ZN(n514) );
  AND2_X1 U560 ( .A1(n871), .A2(G114), .ZN(n515) );
  INV_X1 U561 ( .A(KEYINPUT92), .ZN(n684) );
  NOR2_X1 U562 ( .A1(n725), .A2(n724), .ZN(n726) );
  INV_X1 U563 ( .A(KEYINPUT32), .ZN(n737) );
  XNOR2_X1 U564 ( .A(n738), .B(n737), .ZN(n746) );
  INV_X1 U565 ( .A(KEYINPUT90), .ZN(n680) );
  INV_X1 U566 ( .A(KEYINPUT69), .ZN(n565) );
  INV_X1 U567 ( .A(KEYINPUT99), .ZN(n768) );
  XNOR2_X1 U568 ( .A(n566), .B(n565), .ZN(n567) );
  NOR2_X1 U569 ( .A1(G164), .A2(G1384), .ZN(n772) );
  INV_X1 U570 ( .A(KEYINPUT65), .ZN(n521) );
  BUF_X1 U571 ( .A(n600), .Z(n878) );
  NOR2_X1 U572 ( .A1(G543), .A2(G651), .ZN(n636) );
  NOR2_X1 U573 ( .A1(n652), .A2(n545), .ZN(n639) );
  NOR2_X1 U574 ( .A1(n652), .A2(G651), .ZN(n646) );
  INV_X1 U575 ( .A(KEYINPUT84), .ZN(n525) );
  XNOR2_X1 U576 ( .A(n526), .B(n525), .ZN(n527) );
  AND2_X1 U577 ( .A1(n528), .A2(n527), .ZN(G164) );
  XOR2_X2 U578 ( .A(G2104), .B(KEYINPUT64), .Z(n520) );
  AND2_X1 U579 ( .A1(n520), .A2(G2105), .ZN(n870) );
  NAND2_X1 U580 ( .A1(G126), .A2(n870), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(KEYINPUT83), .ZN(n517) );
  NOR2_X1 U582 ( .A1(n517), .A2(n515), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n601), .A2(G138), .ZN(n524) );
  NOR2_X2 U584 ( .A1(n520), .A2(G2105), .ZN(n522) );
  NAND2_X1 U585 ( .A1(n600), .A2(G102), .ZN(n523) );
  NAND2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n526) );
  NAND2_X1 U587 ( .A1(n871), .A2(G113), .ZN(n529) );
  XNOR2_X1 U588 ( .A(n529), .B(KEYINPUT66), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U590 ( .A(n532), .B(KEYINPUT67), .ZN(n534) );
  NAND2_X1 U591 ( .A1(G125), .A2(n870), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n538) );
  AND2_X2 U593 ( .A1(G101), .A2(n600), .ZN(n536) );
  INV_X1 U594 ( .A(KEYINPUT23), .ZN(n535) );
  XNOR2_X1 U595 ( .A(n536), .B(n535), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n538), .A2(n537), .ZN(n679) );
  BUF_X1 U597 ( .A(n679), .Z(G160) );
  NAND2_X1 U598 ( .A1(n636), .A2(G89), .ZN(n540) );
  XNOR2_X1 U599 ( .A(KEYINPUT4), .B(n540), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT0), .B(G543), .Z(n652) );
  INV_X1 U601 ( .A(G651), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n639), .A2(G76), .ZN(n541) );
  XOR2_X1 U603 ( .A(KEYINPUT73), .B(n541), .Z(n542) );
  NAND2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U605 ( .A(KEYINPUT5), .B(n544), .ZN(n552) );
  NOR2_X1 U606 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U607 ( .A(KEYINPUT1), .B(n546), .Z(n650) );
  NAND2_X1 U608 ( .A1(G63), .A2(n650), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G51), .A2(n646), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n550) );
  XOR2_X1 U611 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n549) );
  XNOR2_X1 U612 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U614 ( .A(KEYINPUT7), .B(n553), .ZN(G168) );
  XNOR2_X1 U615 ( .A(G168), .B(KEYINPUT8), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U617 ( .A1(G64), .A2(n650), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G52), .A2(n646), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G90), .A2(n636), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G77), .A2(n639), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U624 ( .A1(n561), .A2(n560), .ZN(G171) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U629 ( .A(G223), .ZN(n823) );
  NAND2_X1 U630 ( .A1(n823), .A2(G567), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U632 ( .A1(G56), .A2(n650), .ZN(n564) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n564), .Z(n572) );
  NAND2_X1 U634 ( .A1(G81), .A2(n636), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G68), .A2(n639), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(n570), .Z(n571) );
  NOR2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n646), .A2(G43), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n947) );
  INV_X1 U642 ( .A(G860), .ZN(n613) );
  OR2_X1 U643 ( .A1(n947), .A2(n613), .ZN(G153) );
  XOR2_X1 U644 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U645 ( .A1(G92), .A2(n636), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G66), .A2(n650), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G79), .A2(n639), .ZN(n578) );
  NAND2_X1 U649 ( .A1(G54), .A2(n646), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U652 ( .A(KEYINPUT15), .B(n581), .Z(n944) );
  NOR2_X1 U653 ( .A1(n944), .A2(G868), .ZN(n582) );
  XOR2_X1 U654 ( .A(KEYINPUT72), .B(n582), .Z(n585) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n583) );
  XOR2_X1 U656 ( .A(KEYINPUT71), .B(n583), .Z(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G65), .A2(n650), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G53), .A2(n646), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G91), .A2(n636), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G78), .A2(n639), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n954) );
  INV_X1 U665 ( .A(n954), .ZN(G299) );
  INV_X1 U666 ( .A(G868), .ZN(n663) );
  NOR2_X1 U667 ( .A1(G286), .A2(n663), .ZN(n593) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n592) );
  NOR2_X1 U669 ( .A1(n593), .A2(n592), .ZN(G297) );
  NAND2_X1 U670 ( .A1(G559), .A2(n613), .ZN(n594) );
  XNOR2_X1 U671 ( .A(KEYINPUT76), .B(n594), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n595), .A2(n944), .ZN(n596) );
  XNOR2_X1 U673 ( .A(KEYINPUT16), .B(n596), .ZN(G148) );
  NOR2_X1 U674 ( .A1(G868), .A2(n947), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G868), .A2(n944), .ZN(n597) );
  NOR2_X1 U676 ( .A1(G559), .A2(n597), .ZN(n598) );
  NOR2_X1 U677 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G111), .A2(n871), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G99), .A2(n878), .ZN(n603) );
  NAND2_X1 U680 ( .A1(G135), .A2(n875), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n870), .A2(G123), .ZN(n604) );
  XOR2_X1 U683 ( .A(KEYINPUT18), .B(n604), .Z(n605) );
  NOR2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U686 ( .A(n609), .B(KEYINPUT77), .ZN(n979) );
  XNOR2_X1 U687 ( .A(G2096), .B(n979), .ZN(n611) );
  INV_X1 U688 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U690 ( .A1(G559), .A2(n944), .ZN(n612) );
  XOR2_X1 U691 ( .A(n947), .B(n612), .Z(n660) );
  NAND2_X1 U692 ( .A1(n613), .A2(n660), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G67), .A2(n650), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G55), .A2(n646), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n636), .A2(G93), .ZN(n616) );
  XOR2_X1 U697 ( .A(KEYINPUT78), .B(n616), .Z(n617) );
  NOR2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n639), .A2(G80), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n662) );
  XNOR2_X1 U701 ( .A(n621), .B(n662), .ZN(G145) );
  NAND2_X1 U702 ( .A1(G75), .A2(n639), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G50), .A2(n646), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G88), .A2(n636), .ZN(n624) );
  XNOR2_X1 U706 ( .A(KEYINPUT81), .B(n624), .ZN(n625) );
  NOR2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n650), .A2(G62), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(G303) );
  INV_X1 U710 ( .A(G303), .ZN(G166) );
  NAND2_X1 U711 ( .A1(G60), .A2(n650), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G47), .A2(n646), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G85), .A2(n636), .ZN(n631) );
  XOR2_X1 U715 ( .A(KEYINPUT68), .B(n631), .Z(n632) );
  NOR2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n639), .A2(G72), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(G290) );
  NAND2_X1 U719 ( .A1(G86), .A2(n636), .ZN(n638) );
  NAND2_X1 U720 ( .A1(G61), .A2(n650), .ZN(n637) );
  NAND2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n639), .A2(G73), .ZN(n640) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n640), .Z(n641) );
  NOR2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n646), .A2(G48), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G651), .A2(G74), .ZN(n645) );
  XOR2_X1 U728 ( .A(KEYINPUT79), .B(n645), .Z(n648) );
  NAND2_X1 U729 ( .A1(n646), .A2(G49), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U732 ( .A(n651), .B(KEYINPUT80), .ZN(n654) );
  NAND2_X1 U733 ( .A1(G87), .A2(n652), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(G288) );
  XNOR2_X1 U735 ( .A(G166), .B(KEYINPUT19), .ZN(n656) );
  XNOR2_X1 U736 ( .A(G290), .B(n954), .ZN(n655) );
  XNOR2_X1 U737 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U738 ( .A(n657), .B(G305), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n658), .B(n662), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n659), .B(G288), .ZN(n896) );
  XNOR2_X1 U741 ( .A(n660), .B(n896), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n661), .A2(G868), .ZN(n665) );
  NAND2_X1 U743 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U744 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U751 ( .A1(G132), .A2(G82), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(KEYINPUT22), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n671), .B(KEYINPUT82), .ZN(n672) );
  NOR2_X1 U754 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U755 ( .A1(G96), .A2(n673), .ZN(n827) );
  NAND2_X1 U756 ( .A1(n827), .A2(G2106), .ZN(n677) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U758 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U759 ( .A1(G108), .A2(n675), .ZN(n828) );
  NAND2_X1 U760 ( .A1(n828), .A2(G567), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n829) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U763 ( .A1(n829), .A2(n678), .ZN(n826) );
  NAND2_X1 U764 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U765 ( .A1(n679), .A2(G40), .ZN(n773) );
  XNOR2_X2 U766 ( .A(n773), .B(n680), .ZN(n681) );
  NAND2_X2 U767 ( .A1(n772), .A2(n681), .ZN(n692) );
  NAND2_X1 U768 ( .A1(G8), .A2(n692), .ZN(n764) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n682) );
  XOR2_X1 U770 ( .A(n682), .B(KEYINPUT24), .Z(n683) );
  NOR2_X1 U771 ( .A1(n764), .A2(n683), .ZN(n771) );
  XNOR2_X2 U772 ( .A(n692), .B(n684), .ZN(n714) );
  NAND2_X1 U773 ( .A1(n714), .A2(G2072), .ZN(n685) );
  XNOR2_X1 U774 ( .A(n685), .B(KEYINPUT27), .ZN(n687) );
  INV_X1 U775 ( .A(G1956), .ZN(n999) );
  NOR2_X1 U776 ( .A1(n700), .A2(n999), .ZN(n686) );
  NOR2_X1 U777 ( .A1(n687), .A2(n686), .ZN(n707) );
  NOR2_X1 U778 ( .A1(n954), .A2(n707), .ZN(n689) );
  INV_X1 U779 ( .A(KEYINPUT28), .ZN(n688) );
  XNOR2_X1 U780 ( .A(n689), .B(n688), .ZN(n711) );
  INV_X1 U781 ( .A(G1996), .ZN(n920) );
  NOR2_X2 U782 ( .A1(n692), .A2(n920), .ZN(n691) );
  INV_X1 U783 ( .A(KEYINPUT26), .ZN(n690) );
  XNOR2_X1 U784 ( .A(n691), .B(n690), .ZN(n694) );
  BUF_X2 U785 ( .A(n692), .Z(n729) );
  NAND2_X1 U786 ( .A1(n729), .A2(G1341), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X2 U788 ( .A1(n695), .A2(n947), .ZN(n698) );
  NOR2_X1 U789 ( .A1(n698), .A2(n944), .ZN(n697) );
  INV_X1 U790 ( .A(KEYINPUT94), .ZN(n696) );
  XNOR2_X1 U791 ( .A(n697), .B(n696), .ZN(n706) );
  BUF_X1 U792 ( .A(n698), .Z(n699) );
  NAND2_X1 U793 ( .A1(n944), .A2(n699), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n700), .ZN(n702) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n729), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n954), .A2(n707), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n713) );
  XNOR2_X1 U802 ( .A(KEYINPUT29), .B(KEYINPUT95), .ZN(n712) );
  XNOR2_X1 U803 ( .A(n713), .B(n712), .ZN(n719) );
  XNOR2_X1 U804 ( .A(KEYINPUT25), .B(G2078), .ZN(n919) );
  NAND2_X1 U805 ( .A1(n919), .A2(n714), .ZN(n716) );
  XNOR2_X1 U806 ( .A(KEYINPUT91), .B(G1961), .ZN(n1011) );
  NAND2_X1 U807 ( .A1(n1011), .A2(n729), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U809 ( .A(KEYINPUT93), .B(n717), .Z(n723) );
  NAND2_X1 U810 ( .A1(n723), .A2(G171), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n719), .A2(n718), .ZN(n728) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n764), .ZN(n744) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n729), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n744), .A2(n740), .ZN(n720) );
  NAND2_X1 U815 ( .A1(G8), .A2(n720), .ZN(n721) );
  XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n721), .ZN(n722) );
  NOR2_X1 U817 ( .A1(G168), .A2(n722), .ZN(n725) );
  NOR2_X1 U818 ( .A1(G171), .A2(n723), .ZN(n724) );
  XOR2_X1 U819 ( .A(KEYINPUT31), .B(n726), .Z(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n739) );
  NAND2_X1 U821 ( .A1(n739), .A2(G286), .ZN(n735) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n729), .ZN(n731) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n764), .ZN(n730) );
  NOR2_X1 U824 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U825 ( .A1(n732), .A2(G303), .ZN(n733) );
  XNOR2_X1 U826 ( .A(n733), .B(KEYINPUT96), .ZN(n734) );
  NAND2_X1 U827 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U828 ( .A1(n736), .A2(G8), .ZN(n738) );
  BUF_X1 U829 ( .A(n739), .Z(n742) );
  NAND2_X1 U830 ( .A1(G8), .A2(n740), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X2 U833 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U834 ( .A(n747), .B(KEYINPUT97), .ZN(n761) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n755) );
  NOR2_X1 U836 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U837 ( .A1(n755), .A2(n748), .ZN(n959) );
  INV_X1 U838 ( .A(KEYINPUT33), .ZN(n752) );
  AND2_X1 U839 ( .A1(n959), .A2(n752), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n761), .A2(n749), .ZN(n753) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n945) );
  INV_X1 U842 ( .A(n764), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n945), .A2(n750), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U845 ( .A1(n764), .A2(n756), .ZN(n758) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n941) );
  INV_X1 U847 ( .A(n941), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n767) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n761), .A2(n763), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n769) );
  XNOR2_X1 U855 ( .A(n769), .B(n768), .ZN(n770) );
  NOR2_X1 U856 ( .A1(n772), .A2(n773), .ZN(n818) );
  NAND2_X1 U857 ( .A1(G104), .A2(n878), .ZN(n775) );
  NAND2_X1 U858 ( .A1(G140), .A2(n875), .ZN(n774) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n776), .ZN(n782) );
  NAND2_X1 U861 ( .A1(G128), .A2(n870), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G116), .A2(n871), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U864 ( .A(KEYINPUT85), .B(n779), .ZN(n780) );
  XNOR2_X1 U865 ( .A(KEYINPUT35), .B(n780), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n783), .ZN(n892) );
  XNOR2_X1 U868 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  NOR2_X1 U869 ( .A1(n892), .A2(n816), .ZN(n974) );
  NAND2_X1 U870 ( .A1(n818), .A2(n974), .ZN(n814) );
  NAND2_X1 U871 ( .A1(G105), .A2(n878), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT38), .ZN(n791) );
  NAND2_X1 U873 ( .A1(G141), .A2(n875), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G117), .A2(n871), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n870), .A2(G129), .ZN(n787) );
  XOR2_X1 U877 ( .A(KEYINPUT88), .B(n787), .Z(n788) );
  NOR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n891) );
  NAND2_X1 U880 ( .A1(G1996), .A2(n891), .ZN(n801) );
  NAND2_X1 U881 ( .A1(n870), .A2(G119), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G131), .A2(n875), .ZN(n793) );
  NAND2_X1 U883 ( .A1(G107), .A2(n871), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n878), .A2(G95), .ZN(n794) );
  XOR2_X1 U886 ( .A(KEYINPUT86), .B(n794), .Z(n795) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U889 ( .A(KEYINPUT87), .B(n799), .Z(n885) );
  NAND2_X1 U890 ( .A1(G1991), .A2(n885), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U892 ( .A(KEYINPUT89), .B(n802), .ZN(n986) );
  INV_X1 U893 ( .A(n986), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n803), .A2(n818), .ZN(n809) );
  NAND2_X1 U895 ( .A1(n814), .A2(n809), .ZN(n804) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n958) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n891), .ZN(n982) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n885), .ZN(n806) );
  XOR2_X1 U899 ( .A(KEYINPUT101), .B(n806), .Z(n973) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n807) );
  XNOR2_X1 U901 ( .A(KEYINPUT100), .B(n807), .ZN(n808) );
  NOR2_X1 U902 ( .A1(n973), .A2(n808), .ZN(n811) );
  INV_X1 U903 ( .A(n809), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n982), .A2(n812), .ZN(n813) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n813), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n892), .A2(n816), .ZN(n977) );
  NAND2_X1 U909 ( .A1(n817), .A2(n977), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U912 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U915 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U919 ( .A(G132), .ZN(G219) );
  INV_X1 U920 ( .A(G120), .ZN(G236) );
  INV_X1 U921 ( .A(G82), .ZN(G220) );
  INV_X1 U922 ( .A(G69), .ZN(G235) );
  NOR2_X1 U923 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  INV_X1 U925 ( .A(n829), .ZN(G319) );
  XOR2_X1 U926 ( .A(KEYINPUT105), .B(G1976), .Z(n831) );
  XNOR2_X1 U927 ( .A(G1986), .B(G1971), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U929 ( .A(n832), .B(G2474), .Z(n834) );
  XNOR2_X1 U930 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U932 ( .A(G1961), .B(G1956), .Z(n836) );
  XNOR2_X1 U933 ( .A(G1981), .B(G1966), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U938 ( .A(G2096), .B(KEYINPUT43), .Z(n842) );
  XNOR2_X1 U939 ( .A(G2090), .B(G2678), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(n843), .B(KEYINPUT42), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U944 ( .A(KEYINPUT104), .B(G2100), .Z(n847) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(G227) );
  NAND2_X1 U948 ( .A1(G124), .A2(n870), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n850), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U950 ( .A1(G136), .A2(n875), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G112), .A2(n871), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G100), .A2(n878), .ZN(n853) );
  XNOR2_X1 U954 ( .A(KEYINPUT107), .B(n853), .ZN(n854) );
  NOR2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(KEYINPUT108), .B(n858), .Z(G162) );
  XNOR2_X1 U958 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n860) );
  XNOR2_X1 U959 ( .A(G162), .B(KEYINPUT112), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n889) );
  XNOR2_X1 U961 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G106), .A2(n878), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G142), .A2(n875), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n863), .B(KEYINPUT45), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G130), .A2(n870), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G118), .A2(n871), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n883) );
  NAND2_X1 U971 ( .A1(G127), .A2(n870), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G115), .A2(n871), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n874), .B(KEYINPUT47), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G139), .A2(n875), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G103), .A2(n878), .ZN(n879) );
  XNOR2_X1 U978 ( .A(KEYINPUT111), .B(n879), .ZN(n880) );
  NOR2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n969) );
  XNOR2_X1 U980 ( .A(n969), .B(n979), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n887) );
  XNOR2_X1 U983 ( .A(G164), .B(G160), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U985 ( .A(n889), .B(n888), .Z(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n893) );
  XOR2_X1 U987 ( .A(n893), .B(n892), .Z(n894) );
  NOR2_X1 U988 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U989 ( .A(n944), .B(G286), .Z(n895) );
  XNOR2_X1 U990 ( .A(n947), .B(n895), .ZN(n898) );
  XOR2_X1 U991 ( .A(G171), .B(n896), .Z(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U993 ( .A1(G37), .A2(n899), .ZN(G397) );
  XNOR2_X1 U994 ( .A(G2454), .B(G2443), .ZN(n909) );
  XOR2_X1 U995 ( .A(G2430), .B(KEYINPUT102), .Z(n901) );
  XNOR2_X1 U996 ( .A(G2446), .B(KEYINPUT103), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U998 ( .A(G2451), .B(G2427), .Z(n903) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1001 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G2435), .B(G2438), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  NAND2_X1 U1005 ( .A1(n910), .A2(G14), .ZN(n916) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n916), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n916), .ZN(G401) );
  XNOR2_X1 U1016 ( .A(G2067), .B(G26), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(G2072), .B(G33), .ZN(n917) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(n919), .B(G27), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n920), .B(G32), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n926) );
  XOR2_X1 U1022 ( .A(G1991), .B(G25), .Z(n923) );
  NAND2_X1 U1023 ( .A1(n923), .A2(G28), .ZN(n924) );
  XOR2_X1 U1024 ( .A(KEYINPUT117), .B(n924), .Z(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(KEYINPUT53), .B(n929), .ZN(n933) );
  XOR2_X1 U1028 ( .A(G34), .B(KEYINPUT118), .Z(n931) );
  XNOR2_X1 U1029 ( .A(G2084), .B(KEYINPUT54), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(n931), .B(n930), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT116), .B(G2090), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(G35), .B(n934), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(n937), .B(KEYINPUT55), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G29), .B(KEYINPUT119), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(G11), .A2(n940), .ZN(n967) );
  XOR2_X1 U1039 ( .A(G16), .B(KEYINPUT56), .Z(n964) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G168), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(n943), .B(KEYINPUT57), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(n944), .B(G1348), .ZN(n946) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n951) );
  XOR2_X1 U1045 ( .A(n947), .B(G1341), .Z(n949) );
  XNOR2_X1 U1046 ( .A(G171), .B(G1961), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n962) );
  XNOR2_X1 U1050 ( .A(n954), .B(G1956), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(G1971), .A2(G303), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(n965), .B(KEYINPUT120), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n997) );
  XNOR2_X1 U1059 ( .A(G164), .B(G2078), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n968), .B(KEYINPUT115), .ZN(n971) );
  XOR2_X1 U1061 ( .A(G2072), .B(n969), .Z(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1063 ( .A(KEYINPUT50), .B(n972), .Z(n991) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n981) );
  XOR2_X1 U1065 ( .A(G160), .B(G2084), .Z(n975) );
  XNOR2_X1 U1066 ( .A(KEYINPUT113), .B(n975), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n988) );
  XOR2_X1 U1070 ( .A(G2090), .B(G162), .Z(n983) );
  NOR2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1072 ( .A(KEYINPUT51), .B(n984), .Z(n985) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1075 ( .A(KEYINPUT114), .B(n989), .Z(n990) );
  NOR2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1077 ( .A(KEYINPUT52), .B(n992), .ZN(n994) );
  INV_X1 U1078 ( .A(KEYINPUT55), .ZN(n993) );
  NAND2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1080 ( .A1(n995), .A2(G29), .ZN(n996) );
  NAND2_X1 U1081 ( .A1(n997), .A2(n996), .ZN(n1026) );
  XNOR2_X1 U1082 ( .A(KEYINPUT59), .B(G1348), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(n998), .B(G4), .ZN(n1005) );
  XOR2_X1 U1084 ( .A(G1981), .B(G6), .Z(n1001) );
  XNOR2_X1 U1085 ( .A(n999), .B(G20), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XNOR2_X1 U1087 ( .A(G19), .B(G1341), .ZN(n1002) );
  NOR2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1089 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1090 ( .A(KEYINPUT121), .B(KEYINPUT60), .Z(n1006) );
  XNOR2_X1 U1091 ( .A(n1007), .B(n1006), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1008) );
  NOR2_X1 U1093 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(KEYINPUT122), .B(n1010), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(n1011), .B(G5), .ZN(n1012) );
  NAND2_X1 U1096 ( .A1(n1013), .A2(n1012), .ZN(n1022) );
  XNOR2_X1 U1097 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(n1014), .B(KEYINPUT58), .ZN(n1020) );
  XOR2_X1 U1099 ( .A(G1986), .B(G24), .Z(n1018) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(n1020), .B(n1019), .Z(n1021) );
  NOR2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1023), .Z(n1024) );
  NOR2_X1 U1107 ( .A1(G16), .A2(n1024), .ZN(n1025) );
  NOR2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XOR2_X1 U1109 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n1027) );
  XNOR2_X1 U1110 ( .A(n1028), .B(n1027), .ZN(G311) );
  XOR2_X1 U1111 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

