//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT95), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT96), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G134gat), .B(G162gat), .Z(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT41), .ZN(new_n208));
  INV_X1    g007(.A(G232gat), .ZN(new_n209));
  INV_X1    g008(.A(G233gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n207), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT83), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT83), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n219), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT84), .ZN(new_n223));
  NAND2_X1  g022(.A1(G29gat), .A2(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G43gat), .B(G50gat), .Z(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(new_n227), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n217), .B(KEYINPUT86), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n221), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n224), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G99gat), .B(G106gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT92), .ZN(new_n240));
  NAND2_X1  g039(.A1(G99gat), .A2(G106gat), .ZN(new_n241));
  INV_X1    g040(.A(G85gat), .ZN(new_n242));
  INV_X1    g041(.A(G92gat), .ZN(new_n243));
  AOI22_X1  g042(.A1(KEYINPUT8), .A2(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT7), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT92), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n239), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n244), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT93), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n240), .A2(KEYINPUT93), .A3(new_n244), .A4(new_n246), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n229), .A2(KEYINPUT17), .A3(new_n235), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n238), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT94), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n236), .A2(new_n255), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n238), .A2(KEYINPUT94), .A3(new_n256), .A4(new_n257), .ZN(new_n262));
  NAND3_X1  g061(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n260), .A2(new_n261), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n203), .A2(new_n204), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n213), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n266), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT91), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n212), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT16), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(G1gat), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(G1gat), .B2(new_n275), .ZN(new_n278));
  INV_X1    g077(.A(G8gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G57gat), .B(G64gat), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G78gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n281), .B1(KEYINPUT21), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G231gat), .A2(G233gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n288), .B(KEYINPUT90), .Z(new_n289));
  XOR2_X1   g088(.A(new_n289), .B(KEYINPUT19), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n287), .B(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G127gat), .B(G155gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n286), .A2(KEYINPUT21), .ZN(new_n294));
  XNOR2_X1  g093(.A(G183gat), .B(G211gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n293), .B(new_n298), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n274), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT18), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n302), .A2(new_n303), .B1(G229gat), .B2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n238), .A2(new_n305), .A3(new_n280), .A4(new_n257), .ZN(new_n306));
  INV_X1    g105(.A(new_n257), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT17), .B1(new_n229), .B2(new_n235), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n307), .A2(new_n308), .A3(new_n281), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n280), .B1(new_n229), .B2(new_n235), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(KEYINPUT87), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n304), .B(new_n306), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n302), .A2(new_n303), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n238), .A2(new_n280), .A3(new_n257), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(KEYINPUT87), .B2(new_n310), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n317), .A2(new_n313), .A3(new_n304), .A4(new_n306), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n236), .B(new_n281), .ZN(new_n319));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n320), .B(KEYINPUT13), .Z(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n315), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G113gat), .B(G141gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(G197gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(KEYINPUT11), .ZN(new_n326));
  INV_X1    g125(.A(G169gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT12), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n315), .A2(new_n318), .A3(new_n329), .A4(new_n322), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n335), .B(KEYINPUT99), .Z(new_n336));
  AND3_X1   g135(.A1(new_n247), .A2(KEYINPUT97), .A3(new_n251), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n251), .B1(new_n247), .B2(KEYINPUT97), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n286), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n286), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n253), .A2(new_n342), .A3(new_n254), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n286), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n336), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n339), .B2(new_n343), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G120gat), .B(G148gat), .ZN(new_n350));
  INV_X1    g149(.A(G176gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G204gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n349), .B(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n334), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT0), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G57gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(new_n242), .ZN(new_n362));
  INV_X1    g161(.A(G134gat), .ZN(new_n363));
  INV_X1    g162(.A(G127gat), .ZN(new_n364));
  INV_X1    g163(.A(G120gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G113gat), .ZN(new_n366));
  INV_X1    g165(.A(G113gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G120gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n364), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g170(.A(KEYINPUT1), .B(G127gat), .C1(new_n366), .C2(new_n368), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n363), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G141gat), .B(G148gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT2), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(G155gat), .B2(G162gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n376), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G141gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G148gat), .ZN(new_n382));
  INV_X1    g181(.A(G148gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G141gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G155gat), .B(G162gat), .ZN(new_n386));
  INV_X1    g185(.A(G155gat), .ZN(new_n387));
  INV_X1    g186(.A(G162gat), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT2), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n380), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G113gat), .B(G120gat), .ZN(new_n392));
  OAI21_X1  g191(.A(G127gat), .B1(new_n392), .B2(KEYINPUT1), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n369), .A2(new_n370), .A3(new_n364), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(G134gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n373), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT71), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT71), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n396), .A2(new_n399), .A3(KEYINPUT4), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n373), .A2(new_n391), .A3(new_n401), .A4(new_n395), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT72), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n393), .A2(new_n394), .A3(G134gat), .ZN(new_n404));
  AOI21_X1  g203(.A(G134gat), .B1(new_n393), .B2(new_n394), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT72), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n401), .A4(new_n391), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n398), .A2(new_n400), .A3(new_n403), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n373), .A2(new_n395), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n380), .A2(new_n390), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n409), .A2(new_n410), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n414), .B1(new_n404), .B2(new_n405), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n396), .ZN(new_n419));
  INV_X1    g218(.A(new_n410), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT73), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n410), .B1(new_n418), .B2(new_n396), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n417), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n420), .A2(KEYINPUT5), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT74), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n402), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n397), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n402), .B2(new_n430), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n402), .A2(new_n430), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT75), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n397), .B1(new_n438), .B2(new_n432), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n416), .B(new_n429), .C1(new_n436), .C2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n362), .B1(new_n428), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT6), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT25), .ZN(new_n445));
  NOR2_X1   g244(.A1(G169gat), .A2(G176gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT23), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT24), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(G183gat), .A3(G190gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(G169gat), .A2(G176gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT24), .ZN(new_n452));
  NOR2_X1   g251(.A1(G183gat), .A2(G190gat), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n449), .B(new_n450), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n445), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT23), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n446), .B(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n449), .A2(new_n450), .ZN(new_n458));
  INV_X1    g257(.A(new_n453), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(KEYINPUT24), .A3(new_n451), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT25), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT64), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n327), .A2(new_n351), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(KEYINPUT26), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(KEYINPUT26), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT26), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n446), .A2(KEYINPUT64), .A3(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n465), .A2(new_n450), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT27), .B(G183gat), .ZN(new_n470));
  INV_X1    g269(.A(G190gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT28), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT28), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n470), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n469), .A2(new_n473), .A3(new_n451), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n462), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(G226gat), .A2(G233gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(G211gat), .A2(G218gat), .ZN(new_n480));
  INV_X1    g279(.A(G211gat), .ZN(new_n481));
  INV_X1    g280(.A(G218gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(G197gat), .B(G204gat), .Z(new_n484));
  INV_X1    g283(.A(KEYINPUT22), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n480), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT68), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n483), .A2(new_n485), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(G211gat), .B2(G218gat), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n490), .A2(new_n484), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n487), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT29), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n462), .B2(new_n476), .ZN(new_n495));
  OR3_X1    g294(.A1(new_n479), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n479), .B2(new_n495), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT37), .ZN(new_n499));
  XNOR2_X1  g298(.A(G8gat), .B(G36gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT69), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n501), .B(G64gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(new_n243), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n498), .A2(KEYINPUT37), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n504), .A2(KEYINPUT38), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n498), .A2(new_n503), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509));
  AOI211_X1 g308(.A(new_n509), .B(new_n362), .C1(new_n428), .C2(new_n440), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n428), .A2(new_n440), .A3(new_n362), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(new_n441), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n512), .B2(new_n509), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n444), .B(new_n508), .C1(new_n513), .C2(new_n443), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT80), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT81), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n505), .B1(new_n504), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n517), .B2(new_n504), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT38), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n428), .A2(new_n440), .ZN(new_n521));
  INV_X1    g320(.A(new_n362), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n428), .A2(new_n440), .A3(new_n362), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n509), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n442), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT79), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n527), .A2(KEYINPUT80), .A3(new_n444), .A4(new_n508), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n516), .A2(new_n520), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G78gat), .B(G106gat), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(G22gat), .Z(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT29), .B1(new_n391), .B2(new_n412), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n493), .A2(KEYINPUT77), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT77), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n533), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT29), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT3), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n535), .B(new_n538), .C1(new_n540), .C2(new_n391), .ZN(new_n541));
  INV_X1    g340(.A(G228gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n210), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G50gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT29), .B1(new_n491), .B2(new_n486), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n414), .B1(new_n547), .B2(KEYINPUT3), .ZN(new_n548));
  OAI221_X1 g347(.A(new_n548), .B1(new_n542), .B2(new_n210), .C1(new_n533), .C2(new_n537), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n546), .B1(new_n544), .B2(new_n549), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n532), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n531), .A3(new_n550), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n416), .B1(new_n436), .B2(new_n439), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n420), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n558), .B(KEYINPUT39), .C1(new_n420), .C2(new_n419), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n559), .B(new_n362), .C1(KEYINPUT39), .C2(new_n558), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT40), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n523), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n507), .A2(KEYINPUT30), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n503), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n565), .A2(KEYINPUT30), .A3(new_n497), .A4(new_n496), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n498), .A2(new_n503), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n560), .A2(new_n561), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n556), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n529), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n553), .A2(new_n555), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT70), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n568), .B(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n526), .A2(new_n578), .A3(new_n564), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n563), .B1(new_n525), .B2(new_n442), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(KEYINPUT76), .A3(new_n578), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n576), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G227gat), .A2(G233gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n477), .A2(new_n411), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n406), .A2(new_n462), .A3(new_n476), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT32), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT65), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n585), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n477), .A2(new_n411), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n462), .A2(new_n476), .B1(new_n373), .B2(new_n395), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT65), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT32), .ZN(new_n596));
  XNOR2_X1  g395(.A(G15gat), .B(G43gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G71gat), .ZN(new_n598));
  INV_X1    g397(.A(G99gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n590), .A2(new_n596), .A3(new_n600), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n594), .A2(KEYINPUT32), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT67), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n603), .B2(new_n605), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n592), .A2(new_n591), .A3(new_n593), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT34), .B1(new_n591), .B2(KEYINPUT66), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n603), .A2(new_n605), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n613), .A2(new_n606), .A3(new_n611), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT36), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT78), .B1(new_n584), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n582), .A2(KEYINPUT76), .A3(new_n578), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT76), .B1(new_n582), .B2(new_n578), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n556), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT78), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n608), .A2(new_n611), .ZN(new_n622));
  INV_X1    g421(.A(new_n607), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n613), .A2(new_n606), .A3(new_n611), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT36), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n620), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n575), .A2(new_n617), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT82), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(new_n615), .B2(new_n556), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(KEYINPUT82), .A3(new_n576), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n581), .A2(new_n631), .A3(new_n632), .A4(new_n583), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT35), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n570), .B1(new_n527), .B2(new_n444), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT35), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n615), .A2(new_n556), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  AOI211_X1 g438(.A(new_n301), .B(new_n358), .C1(new_n629), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n513), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g441(.A1(new_n276), .A2(new_n279), .ZN(new_n643));
  NAND2_X1  g442(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n644));
  AND4_X1   g443(.A1(new_n570), .A2(new_n640), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n279), .B1(new_n640), .B2(new_n570), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT42), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(KEYINPUT42), .B2(new_n645), .ZN(G1325gat));
  AOI21_X1  g447(.A(G15gat), .B1(new_n640), .B2(new_n626), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n616), .B(KEYINPUT100), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n651), .A2(G15gat), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n640), .B2(new_n652), .ZN(G1326gat));
  NAND2_X1  g452(.A1(new_n640), .A2(new_n556), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT43), .B(G22gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n629), .A2(new_n639), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n269), .A2(new_n273), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n584), .A2(new_n616), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n575), .A2(new_n661), .B1(new_n634), .B2(new_n638), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n663));
  NOR3_X1   g462(.A1(new_n662), .A2(new_n274), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n358), .A2(new_n300), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(G29gat), .B1(new_n667), .B2(new_n526), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n658), .A2(new_n659), .A3(new_n666), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(new_n215), .A3(new_n513), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT45), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(G1328gat));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n216), .A3(new_n570), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT46), .Z(new_n674));
  OAI21_X1  g473(.A(G36gat), .B1(new_n667), .B2(new_n571), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(G1329gat));
  INV_X1    g475(.A(G43gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n669), .A2(new_n677), .A3(new_n626), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT102), .Z(new_n679));
  OAI21_X1  g478(.A(G43gat), .B1(new_n667), .B2(new_n627), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(KEYINPUT47), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G43gat), .B1(new_n667), .B2(new_n650), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n683), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g483(.A(G50gat), .B1(new_n667), .B2(new_n576), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT48), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(G50gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n688), .A3(new_n556), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n685), .B(new_n689), .C1(new_n686), .C2(KEYINPUT48), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1331gat));
  INV_X1    g492(.A(new_n356), .ZN(new_n694));
  NOR4_X1   g493(.A1(new_n662), .A2(new_n301), .A3(new_n333), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n513), .B(KEYINPUT104), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(new_n570), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT105), .Z(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1333gat));
  NAND2_X1  g502(.A1(new_n695), .A2(new_n651), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n615), .A2(G71gat), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n704), .A2(G71gat), .B1(new_n695), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g506(.A1(new_n695), .A2(new_n556), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT106), .B(G78gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1335gat));
  NOR2_X1   g509(.A1(new_n300), .A2(new_n333), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n694), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n665), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G85gat), .B1(new_n714), .B2(new_n526), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n575), .A2(new_n661), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n274), .B1(new_n717), .B2(new_n639), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n718), .B2(new_n711), .ZN(new_n719));
  NOR4_X1   g518(.A1(new_n662), .A2(KEYINPUT51), .A3(new_n274), .A4(new_n712), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n356), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n513), .A2(new_n242), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n715), .B1(new_n725), .B2(new_n726), .ZN(G1336gat));
  OAI21_X1  g526(.A(G92gat), .B1(new_n714), .B2(new_n571), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n620), .A2(new_n627), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n574), .B2(new_n529), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n634), .A2(new_n638), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n659), .B(new_n711), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n719), .B2(new_n720), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(KEYINPUT108), .A3(new_n716), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n694), .A2(new_n571), .A3(G92gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n728), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT52), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(new_n721), .B2(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(G1337gat));
  OAI21_X1  g541(.A(G99gat), .B1(new_n714), .B2(new_n650), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n626), .A2(new_n599), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n725), .B2(new_n744), .ZN(G1338gat));
  NOR3_X1   g544(.A1(new_n694), .A2(new_n576), .A3(G106gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n734), .A2(new_n735), .A3(new_n746), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n556), .B(new_n713), .C1(new_n660), .C2(new_n664), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G106gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT53), .B1(new_n721), .B2(new_n746), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n752), .A2(new_n749), .A3(KEYINPUT109), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT109), .B1(new_n752), .B2(new_n749), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT110), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n751), .B(new_n757), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1339gat));
  NAND2_X1  g558(.A1(new_n344), .A2(new_n345), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n347), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n344), .A2(new_n336), .A3(new_n345), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(KEYINPUT54), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n355), .B1(new_n346), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n766), .A2(KEYINPUT112), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT112), .B1(new_n766), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n763), .A2(new_n765), .A3(KEYINPUT55), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n349), .A2(new_n355), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n763), .A2(new_n765), .A3(KEYINPUT111), .A4(KEYINPUT55), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n333), .A2(new_n770), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n320), .B1(new_n317), .B2(new_n306), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n319), .A2(new_n321), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n328), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n332), .A2(new_n780), .A3(new_n356), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n659), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n332), .A2(new_n780), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n659), .A2(new_n783), .A3(new_n770), .A4(new_n776), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n299), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n274), .A2(new_n300), .A3(new_n334), .A4(new_n694), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n786), .B2(new_n787), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n526), .A2(new_n570), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n637), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n334), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n367), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT114), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n795), .A2(KEYINPUT114), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n791), .A2(new_n696), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n631), .A2(new_n632), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n571), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n333), .A2(new_n367), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT115), .Z(new_n803));
  OAI22_X1  g602(.A1(new_n797), .A2(new_n798), .B1(new_n801), .B2(new_n803), .ZN(G1340gat));
  OAI21_X1  g603(.A(G120gat), .B1(new_n793), .B2(new_n694), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n356), .A2(new_n365), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n801), .B2(new_n806), .ZN(G1341gat));
  NOR3_X1   g606(.A1(new_n793), .A2(new_n364), .A3(new_n299), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n801), .A2(new_n299), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n364), .ZN(G1342gat));
  OAI21_X1  g609(.A(G134gat), .B1(new_n793), .B2(new_n274), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n801), .A2(G134gat), .ZN(new_n812));
  XNOR2_X1  g611(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n812), .A2(new_n659), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n812), .B2(new_n659), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(G1343gat));
  NAND2_X1  g615(.A1(new_n766), .A2(new_n767), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n333), .A2(new_n776), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n783), .A2(new_n819), .A3(new_n356), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n781), .A2(KEYINPUT117), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n818), .A2(new_n820), .A3(KEYINPUT118), .A4(new_n821), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n274), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n300), .B1(new_n826), .B2(new_n784), .ZN(new_n827));
  INV_X1    g626(.A(new_n787), .ZN(new_n828));
  OAI211_X1 g627(.A(KEYINPUT57), .B(new_n556), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n789), .A2(new_n790), .A3(new_n576), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(KEYINPUT57), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n784), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n299), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n576), .B1(new_n834), .B2(new_n787), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n627), .A2(new_n792), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n832), .A2(new_n836), .A3(new_n333), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G141gat), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n651), .A2(new_n576), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n791), .A2(new_n696), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n334), .A2(G141gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n571), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT58), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT58), .B1(new_n838), .B2(G141gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n799), .A2(KEYINPUT120), .A3(new_n840), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n847), .A2(new_n571), .A3(new_n842), .A4(new_n849), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n846), .A2(KEYINPUT121), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT121), .B1(new_n846), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n845), .B1(new_n851), .B2(new_n852), .ZN(G1344gat));
  NOR2_X1   g652(.A1(new_n694), .A2(G148gat), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n847), .A2(new_n571), .A3(new_n849), .A4(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n832), .A2(new_n836), .A3(new_n837), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT59), .B(new_n383), .C1(new_n856), .C2(new_n356), .ZN(new_n857));
  XOR2_X1   g656(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n858));
  OR2_X1    g657(.A1(new_n835), .A2(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n831), .A2(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n356), .A3(new_n837), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n858), .B1(new_n862), .B2(G148gat), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n855), .B1(new_n857), .B2(new_n863), .ZN(G1345gat));
  NAND4_X1  g663(.A1(new_n847), .A2(new_n300), .A3(new_n571), .A4(new_n849), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n300), .A2(G155gat), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT123), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n865), .A2(new_n387), .B1(new_n856), .B2(new_n867), .ZN(G1346gat));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n571), .A3(new_n849), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n869), .A2(G162gat), .A3(new_n274), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n388), .B1(new_n856), .B2(new_n659), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n870), .A2(new_n871), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n696), .A2(new_n571), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT125), .Z(new_n874));
  NAND3_X1  g673(.A1(new_n791), .A2(new_n637), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G169gat), .B1(new_n875), .B2(new_n334), .ZN(new_n876));
  INV_X1    g675(.A(new_n790), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n879), .A2(KEYINPUT124), .A3(new_n513), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT124), .B1(new_n879), .B2(new_n513), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n800), .A3(new_n881), .A4(new_n570), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n333), .A2(new_n327), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(G1348gat));
  NOR3_X1   g683(.A1(new_n875), .A2(new_n351), .A3(new_n694), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n880), .A2(new_n570), .A3(new_n881), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n356), .A3(new_n800), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n885), .B1(new_n887), .B2(new_n351), .ZN(G1349gat));
  OAI21_X1  g687(.A(G183gat), .B1(new_n875), .B2(new_n299), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n300), .A2(new_n470), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n875), .B2(new_n274), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT61), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n882), .A2(G190gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n659), .ZN(new_n897));
  NOR4_X1   g696(.A1(new_n882), .A2(KEYINPUT126), .A3(G190gat), .A4(new_n274), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(G1351gat));
  AOI21_X1  g698(.A(new_n651), .B1(new_n859), .B2(new_n860), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n874), .ZN(new_n901));
  OAI21_X1  g700(.A(G197gat), .B1(new_n901), .B2(new_n334), .ZN(new_n902));
  AND4_X1   g701(.A1(new_n570), .A2(new_n880), .A3(new_n840), .A4(new_n881), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n334), .A2(G197gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(G1352gat));
  NAND4_X1  g705(.A1(new_n861), .A2(new_n356), .A3(new_n650), .A4(new_n874), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT127), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n900), .A2(KEYINPUT127), .A3(new_n356), .A4(new_n874), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(G204gat), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n903), .A2(new_n353), .A3(new_n356), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT62), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n903), .A2(new_n914), .A3(new_n353), .A4(new_n356), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n913), .A3(new_n915), .ZN(G1353gat));
  NAND3_X1  g715(.A1(new_n903), .A2(new_n481), .A3(new_n300), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n861), .A2(new_n300), .A3(new_n650), .A4(new_n874), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT63), .B1(new_n918), .B2(G211gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1354gat));
  NOR3_X1   g720(.A1(new_n901), .A2(new_n482), .A3(new_n274), .ZN(new_n922));
  AOI21_X1  g721(.A(G218gat), .B1(new_n903), .B2(new_n659), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1355gat));
endmodule


