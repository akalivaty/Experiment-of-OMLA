

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U326 ( .A(n438), .B(n300), .ZN(n301) );
  XNOR2_X1 U327 ( .A(n311), .B(n310), .ZN(n531) );
  XOR2_X1 U328 ( .A(n354), .B(n353), .Z(n294) );
  AND2_X1 U329 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U330 ( .A(n383), .B(KEYINPUT45), .ZN(n384) );
  XNOR2_X1 U331 ( .A(n385), .B(n384), .ZN(n403) );
  XNOR2_X1 U332 ( .A(n352), .B(n295), .ZN(n300) );
  INV_X1 U333 ( .A(n387), .ZN(n304) );
  XNOR2_X1 U334 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U335 ( .A(n355), .B(n294), .ZN(n360) );
  XNOR2_X1 U336 ( .A(n471), .B(KEYINPUT37), .ZN(n472) );
  XNOR2_X1 U337 ( .A(n307), .B(n306), .ZN(n309) );
  XNOR2_X1 U338 ( .A(n360), .B(n359), .ZN(n365) );
  XNOR2_X1 U339 ( .A(n473), .B(n472), .ZN(n516) );
  INV_X1 U340 ( .A(G43GAT), .ZN(n475) );
  XNOR2_X1 U341 ( .A(n474), .B(KEYINPUT38), .ZN(n502) );
  XNOR2_X1 U342 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U343 ( .A(n475), .B(KEYINPUT40), .ZN(n476) );
  XNOR2_X1 U344 ( .A(n453), .B(n452), .ZN(G1349GAT) );
  XNOR2_X1 U345 ( .A(n477), .B(n476), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(KEYINPUT78), .Z(n297) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(G15GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n311) );
  XOR2_X1 U349 ( .A(G183GAT), .B(KEYINPUT17), .Z(n299) );
  XNOR2_X1 U350 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n438) );
  XOR2_X1 U352 ( .A(G190GAT), .B(G134GAT), .Z(n352) );
  XNOR2_X1 U353 ( .A(n301), .B(G176GAT), .ZN(n307) );
  XOR2_X1 U354 ( .A(G127GAT), .B(KEYINPUT77), .Z(n303) );
  XNOR2_X1 U355 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n346) );
  XOR2_X1 U357 ( .A(n346), .B(KEYINPUT79), .Z(n305) );
  XOR2_X1 U358 ( .A(G120GAT), .B(G71GAT), .Z(n387) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G99GAT), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U361 ( .A(G211GAT), .B(KEYINPUT21), .Z(n313) );
  XNOR2_X1 U362 ( .A(G197GAT), .B(KEYINPUT82), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n430) );
  XOR2_X1 U364 ( .A(KEYINPUT23), .B(KEYINPUT83), .Z(n315) );
  XNOR2_X1 U365 ( .A(KEYINPUT22), .B(G204GAT), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n319) );
  XOR2_X1 U367 ( .A(G218GAT), .B(G162GAT), .Z(n356) );
  XOR2_X1 U368 ( .A(KEYINPUT81), .B(n356), .Z(n317) );
  XOR2_X1 U369 ( .A(G141GAT), .B(G22GAT), .Z(n408) );
  XNOR2_X1 U370 ( .A(G50GAT), .B(n408), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n321) );
  NAND2_X1 U373 ( .A1(G228GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n323) );
  INV_X1 U375 ( .A(KEYINPUT24), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n326) );
  XNOR2_X1 U377 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n324), .B(KEYINPUT2), .ZN(n345) );
  XNOR2_X1 U379 ( .A(n345), .B(KEYINPUT80), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n430), .B(n327), .ZN(n329) );
  XOR2_X1 U382 ( .A(G106GAT), .B(G78GAT), .Z(n328) );
  XOR2_X1 U383 ( .A(G148GAT), .B(n328), .Z(n393) );
  XOR2_X1 U384 ( .A(n329), .B(n393), .Z(n464) );
  XOR2_X1 U385 ( .A(G85GAT), .B(G162GAT), .Z(n331) );
  XNOR2_X1 U386 ( .A(G29GAT), .B(G134GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U388 ( .A(KEYINPUT4), .B(G148GAT), .Z(n333) );
  XNOR2_X1 U389 ( .A(G141GAT), .B(G120GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U391 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U392 ( .A(KEYINPUT84), .B(G57GAT), .Z(n337) );
  NAND2_X1 U393 ( .A1(G225GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U395 ( .A(KEYINPUT1), .B(n338), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U397 ( .A(KEYINPUT6), .B(KEYINPUT85), .Z(n342) );
  XNOR2_X1 U398 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(n344), .B(n343), .Z(n348) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n518) );
  XOR2_X1 U403 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n350) );
  XNOR2_X1 U404 ( .A(KEYINPUT70), .B(KEYINPUT9), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n355) );
  XOR2_X1 U407 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n354) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(G92GAT), .ZN(n353) );
  XOR2_X1 U409 ( .A(G99GAT), .B(G85GAT), .Z(n386) );
  XNOR2_X1 U410 ( .A(n386), .B(n356), .ZN(n358) );
  AND2_X1 U411 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U413 ( .A(G29GAT), .B(KEYINPUT8), .Z(n362) );
  XNOR2_X1 U414 ( .A(G43GAT), .B(G36GAT), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U416 ( .A(G50GAT), .B(KEYINPUT7), .Z(n363) );
  XNOR2_X1 U417 ( .A(n364), .B(n363), .ZN(n410) );
  XOR2_X1 U418 ( .A(n365), .B(n410), .Z(n559) );
  INV_X1 U419 ( .A(n559), .ZN(n565) );
  XOR2_X1 U420 ( .A(KEYINPUT36), .B(n565), .Z(n587) );
  XOR2_X1 U421 ( .A(G155GAT), .B(G183GAT), .Z(n367) );
  XNOR2_X1 U422 ( .A(G71GAT), .B(G127GAT), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U424 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n369) );
  XNOR2_X1 U425 ( .A(G64GAT), .B(KEYINPUT73), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U427 ( .A(n371), .B(n370), .Z(n373) );
  XOR2_X1 U428 ( .A(G15GAT), .B(G1GAT), .Z(n415) );
  XOR2_X1 U429 ( .A(G57GAT), .B(KEYINPUT13), .Z(n398) );
  XNOR2_X1 U430 ( .A(n415), .B(n398), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U432 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n375) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U435 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U436 ( .A(G78GAT), .B(G211GAT), .Z(n379) );
  XNOR2_X1 U437 ( .A(G8GAT), .B(G22GAT), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n380), .B(KEYINPUT14), .ZN(n381) );
  XOR2_X1 U440 ( .A(n382), .B(n381), .Z(n579) );
  INV_X1 U441 ( .A(n579), .ZN(n555) );
  NOR2_X1 U442 ( .A1(n587), .A2(n555), .ZN(n385) );
  INV_X1 U443 ( .A(KEYINPUT64), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n402) );
  XOR2_X1 U445 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n389) );
  NAND2_X1 U446 ( .A1(G230GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U448 ( .A(n390), .B(KEYINPUT68), .Z(n395) );
  XOR2_X1 U449 ( .A(G64GAT), .B(G92GAT), .Z(n392) );
  XNOR2_X1 U450 ( .A(G176GAT), .B(G204GAT), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n429) );
  XNOR2_X1 U452 ( .A(n393), .B(n429), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n397) );
  INV_X1 U454 ( .A(KEYINPUT32), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n398), .B(KEYINPUT31), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n576) );
  NOR2_X1 U459 ( .A1(n403), .A2(n576), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n404), .B(KEYINPUT114), .ZN(n418) );
  XOR2_X1 U461 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n406) );
  NAND2_X1 U462 ( .A1(G229GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U464 ( .A(n408), .B(n407), .Z(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U466 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n412) );
  XNOR2_X1 U467 ( .A(G113GAT), .B(G197GAT), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U469 ( .A(n414), .B(n413), .Z(n417) );
  XOR2_X1 U470 ( .A(G169GAT), .B(G8GAT), .Z(n434) );
  XNOR2_X1 U471 ( .A(n434), .B(n415), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n573) );
  XNOR2_X1 U473 ( .A(KEYINPUT67), .B(n573), .ZN(n561) );
  INV_X1 U474 ( .A(n561), .ZN(n533) );
  NAND2_X1 U475 ( .A1(n418), .A2(n533), .ZN(n427) );
  XOR2_X1 U476 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n419) );
  XNOR2_X1 U477 ( .A(KEYINPUT47), .B(n419), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n576), .B(KEYINPUT41), .ZN(n551) );
  NOR2_X1 U479 ( .A1(n573), .A2(n551), .ZN(n421) );
  XNOR2_X1 U480 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n422) );
  NAND2_X1 U482 ( .A1(n422), .A2(n555), .ZN(n423) );
  NOR2_X1 U483 ( .A1(n565), .A2(n423), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  NAND2_X1 U485 ( .A1(n427), .A2(n426), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n428), .B(KEYINPUT48), .ZN(n529) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n442) );
  XOR2_X1 U488 ( .A(KEYINPUT87), .B(G218GAT), .Z(n432) );
  XNOR2_X1 U489 ( .A(G36GAT), .B(G190GAT), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U491 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U492 ( .A1(G226GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U494 ( .A(n437), .B(KEYINPUT86), .Z(n440) );
  XNOR2_X1 U495 ( .A(n438), .B(KEYINPUT88), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U497 ( .A(n442), .B(n441), .Z(n521) );
  INV_X1 U498 ( .A(n521), .ZN(n443) );
  NAND2_X1 U499 ( .A1(n529), .A2(n443), .ZN(n445) );
  XOR2_X1 U500 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U502 ( .A1(n518), .A2(n446), .ZN(n572) );
  NOR2_X1 U503 ( .A1(n464), .A2(n572), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n447), .B(KEYINPUT55), .ZN(n448) );
  NOR2_X1 U505 ( .A1(n531), .A2(n448), .ZN(n449) );
  XOR2_X1 U506 ( .A(KEYINPUT119), .B(n449), .Z(n566) );
  XOR2_X1 U507 ( .A(KEYINPUT104), .B(n551), .Z(n536) );
  NAND2_X1 U508 ( .A1(n566), .A2(n536), .ZN(n453) );
  XOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT57), .Z(n451) );
  XOR2_X1 U510 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n450) );
  XNOR2_X1 U511 ( .A(n521), .B(KEYINPUT27), .ZN(n463) );
  XOR2_X1 U512 ( .A(KEYINPUT90), .B(KEYINPUT26), .Z(n455) );
  AND2_X1 U513 ( .A1(n464), .A2(n531), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n455), .B(n454), .ZN(n571) );
  OR2_X1 U515 ( .A1(n463), .A2(n571), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n531), .A2(n521), .ZN(n456) );
  NOR2_X1 U517 ( .A1(n456), .A2(n464), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n457), .B(KEYINPUT25), .ZN(n459) );
  INV_X1 U519 ( .A(KEYINPUT91), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n461), .A2(n460), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n462), .A2(n518), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n518), .A2(n463), .ZN(n547) );
  INV_X1 U524 ( .A(KEYINPUT28), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(n464), .ZN(n526) );
  NAND2_X1 U526 ( .A1(n547), .A2(n526), .ZN(n530) );
  XNOR2_X1 U527 ( .A(n530), .B(KEYINPUT89), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n466), .A2(n531), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n480) );
  NAND2_X1 U530 ( .A1(n480), .A2(n555), .ZN(n469) );
  XNOR2_X1 U531 ( .A(KEYINPUT98), .B(n469), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n587), .A2(n470), .ZN(n473) );
  XNOR2_X1 U533 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n471) );
  NOR2_X1 U534 ( .A1(n533), .A2(n576), .ZN(n482) );
  NAND2_X1 U535 ( .A1(n516), .A2(n482), .ZN(n474) );
  NOR2_X1 U536 ( .A1(n502), .A2(n531), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(KEYINPUT76), .Z(n479) );
  NAND2_X1 U538 ( .A1(n579), .A2(n559), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(n481) );
  AND2_X1 U540 ( .A1(n481), .A2(n480), .ZN(n506) );
  NAND2_X1 U541 ( .A1(n482), .A2(n506), .ZN(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT92), .B(n483), .ZN(n493) );
  NOR2_X1 U543 ( .A1(n518), .A2(n493), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT94), .B(KEYINPUT34), .Z(n485) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U547 ( .A(n487), .B(n486), .Z(G1324GAT) );
  NOR2_X1 U548 ( .A1(n493), .A2(n521), .ZN(n489) );
  XNOR2_X1 U549 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1325GAT) );
  NOR2_X1 U551 ( .A1(n493), .A2(n531), .ZN(n491) );
  XNOR2_X1 U552 ( .A(KEYINPUT35), .B(KEYINPUT96), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(n492), .ZN(G1326GAT) );
  NOR2_X1 U555 ( .A1(n493), .A2(n526), .ZN(n494) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT97), .B(KEYINPUT39), .Z(n496) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n498) );
  NOR2_X1 U560 ( .A1(n518), .A2(n502), .ZN(n497) );
  XOR2_X1 U561 ( .A(n498), .B(n497), .Z(G1328GAT) );
  NOR2_X1 U562 ( .A1(n502), .A2(n521), .ZN(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  NOR2_X1 U566 ( .A1(n502), .A2(n526), .ZN(n503) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n505) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n508) );
  AND2_X1 U571 ( .A1(n573), .A2(n536), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n517), .A2(n506), .ZN(n512) );
  NOR2_X1 U573 ( .A1(n518), .A2(n512), .ZN(n507) );
  XOR2_X1 U574 ( .A(n508), .B(n507), .Z(G1332GAT) );
  NOR2_X1 U575 ( .A1(n521), .A2(n512), .ZN(n509) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n509), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n531), .A2(n512), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U580 ( .A1(n526), .A2(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n525) );
  NOR2_X1 U585 ( .A1(n518), .A2(n525), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U589 ( .A(KEYINPUT110), .B(n522), .Z(n523) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U591 ( .A1(n531), .A2(n525), .ZN(n524) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n527), .Z(n528) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  BUF_X1 U596 ( .A(n529), .Z(n549) );
  NOR2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U598 ( .A1(n549), .A2(n532), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n533), .A2(n535), .ZN(n534) );
  XOR2_X1 U600 ( .A(G113GAT), .B(n534), .Z(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  INV_X1 U602 ( .A(n535), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n542), .A2(n536), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n540) );
  NAND2_X1 U606 ( .A1(n542), .A2(n579), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n544) );
  NAND2_X1 U610 ( .A1(n542), .A2(n565), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(n545), .ZN(G1343GAT) );
  INV_X1 U613 ( .A(n571), .ZN(n546) );
  AND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n573), .A2(n558), .ZN(n550) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n558), .ZN(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n558), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n566), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT120), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n579), .A2(n566), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n568), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n570) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n575) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n580) );
  INV_X1 U639 ( .A(n580), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n573), .A2(n586), .ZN(n574) );
  XOR2_X1 U641 ( .A(n575), .B(n574), .Z(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U643 ( .A1(n580), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n585) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n589) );
  NOR2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U653 ( .A(n589), .B(n588), .Z(G1355GAT) );
endmodule

