//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n637,
    new_n638, new_n641, new_n643, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1220, new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(new_n439), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n468), .A2(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n475), .B2(G112), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n468), .B2(G2105), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(KEYINPUT68), .A3(new_n475), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  OAI221_X1 g063(.A(new_n480), .B1(new_n481), .B2(new_n482), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n464), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NOR2_X1   g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(new_n475), .B2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n497), .B2(new_n494), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n485), .A2(G126), .A3(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n475), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n485), .A2(KEYINPUT4), .A3(G138), .A4(new_n475), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n499), .A2(new_n500), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT70), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(G651), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(new_n511), .B1(KEYINPUT6), .B2(new_n507), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n512), .A2(G50), .A3(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(KEYINPUT72), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT5), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(new_n507), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n509), .B1(new_n510), .B2(G651), .ZN(new_n524));
  NOR3_X1   g099(.A1(new_n507), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n517), .A2(new_n519), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n514), .A2(new_n522), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND2_X1  g106(.A1(new_n508), .A2(new_n511), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n532), .A2(new_n533), .A3(new_n523), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n533), .B1(new_n532), .B2(new_n523), .ZN(new_n535));
  NOR3_X1   g110(.A1(new_n534), .A2(new_n535), .A3(new_n515), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n512), .A2(G89), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n520), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n537), .A2(new_n540), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n527), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT74), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n549), .B(new_n545), .C1(new_n527), .C2(new_n546), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(G651), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n526), .A2(KEYINPUT73), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n532), .A2(new_n533), .A3(new_n523), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n553), .A2(G52), .A3(G543), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n528), .A2(G90), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n555), .A2(KEYINPUT75), .A3(new_n556), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n552), .B1(new_n559), .B2(new_n560), .ZN(G171));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n517), .B2(new_n519), .ZN(new_n563));
  AND2_X1   g138(.A1(G68), .A2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(KEYINPUT76), .B(G81), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n512), .A2(new_n520), .A3(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n553), .A2(G43), .A3(G543), .A4(new_n554), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  AND3_X1   g147(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G36), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(G188));
  NAND4_X1  g152(.A1(new_n553), .A2(G53), .A3(G543), .A4(new_n554), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G78), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n527), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(G91), .A2(new_n528), .B1(new_n585), .B2(G651), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n534), .A2(new_n535), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n587), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n578), .A2(new_n579), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n582), .A2(new_n586), .A3(new_n591), .ZN(G299));
  AND3_X1   g167(.A1(new_n555), .A2(KEYINPUT75), .A3(new_n556), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT75), .B1(new_n555), .B2(new_n556), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n551), .B1(new_n593), .B2(new_n594), .ZN(G301));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n536), .A2(new_n596), .A3(G49), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n553), .A2(G543), .A3(new_n554), .ZN(new_n598));
  INV_X1    g173(.A(G49), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT78), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n520), .A2(G74), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n528), .A2(G87), .B1(new_n601), .B2(G651), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(G288));
  AND3_X1   g178(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n604));
  INV_X1    g179(.A(G61), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n527), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G73), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n520), .A2(new_n608), .A3(G61), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n604), .B1(new_n610), .B2(G651), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n528), .A2(G86), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(G305));
  NAND2_X1  g188(.A1(new_n536), .A2(G47), .ZN(new_n614));
  NAND2_X1  g189(.A1(G72), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G60), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n527), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(G85), .A2(new_n528), .B1(new_n617), .B2(G651), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n587), .A2(G54), .A3(G543), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n512), .A2(new_n520), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g200(.A1(new_n512), .A2(KEYINPUT10), .A3(G92), .A4(new_n520), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(new_n507), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n621), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT80), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n620), .B1(new_n632), .B2(G868), .ZN(G284));
  OAI21_X1  g208(.A(new_n620), .B1(new_n632), .B2(G868), .ZN(G321));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  OR3_X1    g210(.A1(G168), .A2(KEYINPUT81), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(G299), .A2(new_n635), .ZN(new_n637));
  OAI21_X1  g212(.A(KEYINPUT81), .B1(G168), .B2(new_n635), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(G297));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(G280));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n632), .B1(new_n641), .B2(G860), .ZN(G148));
  AND3_X1   g217(.A1(new_n632), .A2(KEYINPUT82), .A3(new_n641), .ZN(new_n643));
  AOI21_X1  g218(.A(KEYINPUT82), .B1(new_n632), .B2(new_n641), .ZN(new_n644));
  OAI21_X1  g219(.A(G868), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(G868), .B2(new_n571), .ZN(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n479), .A2(G123), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n484), .A2(new_n486), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G135), .ZN(new_n651));
  NOR2_X1   g226(.A1(G99), .A2(G2105), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n649), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n466), .A2(new_n464), .A3(G2105), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n656), .B(new_n657), .Z(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT13), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(new_n660), .ZN(G156));
  XNOR2_X1  g236(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT86), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2451), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2454), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT15), .B(G2435), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT87), .B(G2438), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2427), .B(G2430), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT14), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n665), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1341), .B(G1348), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G14), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G401));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  XOR2_X1   g254(.A(G2067), .B(G2678), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n679), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2096), .B(G2100), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n681), .A2(new_n682), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n689), .A2(new_n683), .A3(KEYINPUT17), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n690), .A2(new_n684), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n688), .B(new_n691), .Z(G227));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(new_n694), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n696), .A2(new_n698), .A3(new_n700), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n703), .B(new_n704), .C1(new_n702), .C2(new_n701), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n705), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT89), .B(G1986), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(G229));
  AND3_X1   g287(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G16), .B2(G23), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT33), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT33), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G1976), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n716), .A2(G1976), .A3(new_n717), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G22), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G166), .B2(new_n723), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT92), .B(G1971), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G6), .B(G305), .S(G16), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT91), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT32), .B(G1981), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n722), .A2(new_n727), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT34), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT34), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n722), .A2(new_n734), .A3(new_n727), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n723), .A2(G24), .ZN(new_n740));
  INV_X1    g315(.A(G290), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(new_n723), .ZN(new_n742));
  INV_X1    g317(.A(G1986), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G25), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n479), .A2(G119), .ZN(new_n747));
  OR2_X1    g322(.A1(G95), .A2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n749));
  INV_X1    g324(.A(G131), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n749), .C1(new_n487), .C2(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(KEYINPUT90), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(KEYINPUT90), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n746), .B1(new_n755), .B2(new_n745), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT35), .B(G1991), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n756), .B(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n737), .A2(new_n739), .A3(new_n744), .A4(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n732), .A2(KEYINPUT34), .B1(KEYINPUT93), .B2(KEYINPUT36), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n761), .A2(new_n744), .A3(new_n735), .A4(new_n759), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(new_n738), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT96), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G2105), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n650), .A2(G139), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  AND3_X1   g345(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G29), .B2(G33), .ZN(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n745), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n745), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT99), .Z(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT29), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(KEYINPUT29), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(G2090), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT100), .ZN(new_n783));
  INV_X1    g358(.A(G2090), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n779), .A2(new_n783), .A3(new_n784), .A4(new_n780), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n723), .A2(G4), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n632), .B2(new_n723), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G1348), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AND3_X1   g364(.A1(new_n723), .A2(KEYINPUT23), .A3(G20), .ZN(new_n790));
  AOI21_X1  g365(.A(KEYINPUT23), .B1(new_n723), .B2(G20), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n790), .B(new_n791), .C1(G299), .C2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1956), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n782), .A2(new_n785), .A3(new_n789), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(G171), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G5), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n787), .ZN(new_n799));
  INV_X1    g374(.A(G1348), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n571), .A2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G16), .B2(G19), .ZN(new_n804));
  INV_X1    g379(.A(G1341), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT100), .B1(new_n781), .B2(G2090), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n654), .A2(new_n745), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT24), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n745), .B1(new_n809), .B2(G34), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(G34), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(new_n811), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n477), .B2(new_n745), .ZN(new_n816));
  INV_X1    g391(.A(G2084), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n745), .A2(G27), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G164), .B2(new_n745), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2078), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT31), .B(G11), .Z(new_n822));
  XOR2_X1   g397(.A(KEYINPUT98), .B(G28), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT30), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n816), .A2(new_n817), .B1(G29), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n807), .A2(new_n808), .A3(new_n818), .A4(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n802), .A2(new_n806), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n796), .A2(new_n797), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(G168), .A2(G16), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G16), .B2(G21), .ZN(new_n833));
  INV_X1    g408(.A(G1966), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n773), .A2(new_n774), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n804), .A2(new_n805), .ZN(new_n837));
  NOR2_X1   g412(.A1(G29), .A2(G32), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n475), .A2(G105), .A3(G2104), .ZN(new_n839));
  NAND3_X1  g414(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT26), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n839), .B(new_n841), .C1(G129), .C2(new_n479), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n650), .A2(G141), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n838), .B1(new_n845), .B2(G29), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT27), .B(G1996), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n833), .A2(new_n834), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n829), .A2(new_n831), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n745), .A2(G26), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n479), .A2(G128), .ZN(new_n854));
  NOR2_X1   g429(.A1(G104), .A2(G2105), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(new_n475), .B2(G116), .ZN(new_n856));
  INV_X1    g431(.A(G140), .ZN(new_n857));
  OAI221_X1 g432(.A(new_n854), .B1(new_n855), .B2(new_n856), .C1(new_n487), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT94), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n853), .B1(new_n860), .B2(new_n745), .ZN(new_n861));
  MUX2_X1   g436(.A(new_n853), .B(new_n861), .S(KEYINPUT28), .Z(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT95), .B(G2067), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n764), .A2(new_n852), .A3(new_n864), .ZN(G311));
  NAND4_X1  g440(.A1(new_n802), .A2(new_n851), .A3(new_n806), .A4(new_n828), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n866), .A2(new_n830), .A3(new_n849), .ZN(new_n867));
  INV_X1    g442(.A(new_n864), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n867), .A2(new_n868), .A3(new_n763), .A4(new_n760), .ZN(G150));
  INV_X1    g444(.A(G67), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n517), .B2(new_n519), .ZN(new_n871));
  AND2_X1   g446(.A1(G80), .A2(G543), .ZN(new_n872));
  OAI21_X1  g447(.A(G651), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n512), .A2(G93), .A3(new_n520), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n553), .A2(G55), .A3(G543), .A4(new_n554), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n632), .A2(G559), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n569), .A3(new_n568), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n570), .A2(new_n876), .A3(new_n875), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n880), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n879), .B1(new_n886), .B2(G860), .ZN(G145));
  XNOR2_X1  g462(.A(new_n654), .B(G160), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(G162), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n771), .A2(new_n505), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G164), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n859), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n859), .B1(new_n891), .B2(new_n893), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n844), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n845), .A3(new_n894), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n903), .B(new_n904), .C1(G118), .C2(new_n475), .ZN(new_n905));
  INV_X1    g480(.A(new_n479), .ZN(new_n906));
  INV_X1    g481(.A(G130), .ZN(new_n907));
  INV_X1    g482(.A(G142), .ZN(new_n908));
  OAI221_X1 g483(.A(new_n905), .B1(new_n906), .B2(new_n907), .C1(new_n487), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n755), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n754), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n658), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n658), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT102), .B1(new_n900), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n899), .A4(new_n897), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n900), .A2(new_n917), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n890), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n889), .B1(new_n923), .B2(KEYINPUT103), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n900), .A2(new_n926), .A3(new_n917), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT104), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n922), .A2(new_n925), .A3(new_n930), .A4(new_n927), .ZN(new_n931));
  AOI211_X1 g506(.A(G37), .B(new_n924), .C1(new_n929), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(G395));
  INV_X1    g509(.A(new_n644), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n632), .A2(KEYINPUT82), .A3(new_n641), .ZN(new_n936));
  INV_X1    g511(.A(new_n883), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n883), .B1(new_n643), .B2(new_n644), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n588), .A2(new_n590), .A3(new_n589), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n590), .B1(new_n588), .B2(new_n589), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n944), .B2(new_n586), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n582), .A2(new_n941), .A3(new_n586), .A4(new_n591), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n621), .A2(new_n627), .A3(new_n629), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(G299), .A2(KEYINPUT105), .A3(new_n630), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n940), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT41), .B1(new_n949), .B2(new_n951), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(G299), .A2(KEYINPUT105), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n947), .A3(new_n946), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT41), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n950), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n957), .A2(new_n958), .A3(new_n950), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n940), .ZN(new_n964));
  XNOR2_X1  g539(.A(G288), .B(G290), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  XOR2_X1   g543(.A(G303), .B(G305), .Z(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n965), .A2(new_n966), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT42), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n974), .A2(KEYINPUT42), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n953), .A2(new_n964), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n974), .B(KEYINPUT42), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n960), .A2(new_n962), .B1(new_n939), .B2(new_n938), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n940), .A2(new_n952), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n981), .A3(G868), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT108), .B1(new_n877), .B2(new_n635), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n977), .A2(new_n981), .A3(KEYINPUT108), .A4(G868), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(KEYINPUT109), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(G295));
  INV_X1    g565(.A(new_n986), .ZN(G331));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g567(.A1(G171), .A2(KEYINPUT110), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n883), .B(G286), .C1(G171), .C2(KEYINPUT110), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g571(.A1(G301), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n883), .B1(new_n997), .B2(G286), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n993), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(G286), .B1(G171), .B2(KEYINPUT110), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n937), .ZN(new_n1001));
  INV_X1    g576(.A(new_n993), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n994), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n952), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n958), .B1(new_n957), .B2(new_n950), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n961), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1007), .B2(new_n1004), .ZN(new_n1008));
  AOI21_X1  g583(.A(G37), .B1(new_n1008), .B2(new_n974), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1004), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n960), .A2(new_n962), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n974), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1005), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1004), .A2(KEYINPUT111), .A3(new_n952), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1009), .A2(new_n1016), .A3(KEYINPUT112), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n992), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1016), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1004), .A2(KEYINPUT111), .A3(new_n952), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT111), .B1(new_n1004), .B2(new_n952), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1012), .B1(new_n1025), .B2(new_n1011), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G37), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT43), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT44), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1011), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n974), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(new_n1028), .A3(new_n1016), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT43), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1009), .A2(new_n1016), .A3(new_n992), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1030), .A2(new_n1039), .ZN(G397));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n611), .A2(new_n1041), .A3(new_n612), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT119), .B(G86), .Z(new_n1043));
  NAND2_X1  g618(.A1(new_n528), .A2(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n611), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n1045), .B2(new_n1041), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1384), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n505), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n471), .A2(new_n476), .A3(G40), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT116), .B(G8), .Z(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT49), .B(new_n1042), .C1(new_n1045), .C2(new_n1041), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1048), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT120), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1048), .A2(new_n1059), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT45), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1051), .B1(new_n1050), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n1049), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1051), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n505), .A2(KEYINPUT50), .A3(new_n1049), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT50), .B1(new_n505), .B2(new_n1049), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT114), .B(G2090), .Z(new_n1070));
  OAI22_X1  g645(.A1(new_n1065), .A2(G1971), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(G8), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(G303), .B2(G8), .ZN(new_n1075));
  INV_X1    g650(.A(G8), .ZN(new_n1076));
  NOR2_X1   g651(.A1(G166), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1055), .B1(G288), .B2(new_n719), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT52), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT117), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n1084), .A3(KEYINPUT52), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n713), .B2(G1976), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1081), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1083), .A2(new_n1085), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1065), .A2(G1966), .B1(G2084), .B2(new_n1069), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1053), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G286), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1061), .A2(new_n1080), .A3(new_n1091), .A4(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1061), .A2(new_n1091), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1079), .A2(G8), .A3(new_n1071), .ZN(new_n1097));
  OR3_X1    g672(.A1(new_n1093), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1079), .B1(new_n1071), .B2(new_n1053), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g675(.A1(KEYINPUT63), .A2(new_n1095), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(G1976), .B(G288), .C1(new_n1058), .C2(new_n1060), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1042), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1055), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT121), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1095), .A2(KEYINPUT63), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1107));
  AND4_X1   g682(.A1(KEYINPUT121), .A2(new_n1104), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1099), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1069), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1111), .A2(new_n817), .B1(new_n834), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G168), .A2(new_n1054), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT123), .B1(new_n1113), .B2(new_n1076), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1115), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1113), .A2(KEYINPUT123), .A3(new_n1076), .ZN(new_n1118));
  OAI221_X1 g693(.A(KEYINPUT51), .B1(new_n1113), .B2(new_n1115), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1093), .A2(new_n1120), .A3(new_n1115), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1063), .A2(KEYINPUT124), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1064), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(G2078), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1063), .A2(KEYINPUT124), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1123), .A2(KEYINPUT53), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1127), .A2(KEYINPUT125), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1063), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n1069), .B2(new_n797), .ZN(new_n1131));
  XNOR2_X1  g706(.A(G171), .B(KEYINPUT54), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1127), .A2(KEYINPUT125), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1131), .B1(new_n1130), .B2(new_n1129), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1132), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1050), .A2(new_n1051), .A3(G2067), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1138), .B(new_n947), .C1(new_n1069), .C2(new_n800), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1069), .A2(new_n800), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1138), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n630), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT60), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n630), .A2(KEYINPUT60), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT58), .B(G1341), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n1112), .A2(G1996), .B1(new_n1052), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1147), .A2(new_n1148), .A3(new_n571), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1147), .B2(new_n571), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1143), .B(new_n1145), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT56), .B(G2072), .ZN(new_n1152));
  INV_X1    g727(.A(G1956), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1065), .A2(new_n1152), .B1(new_n1069), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n588), .A2(new_n589), .A3(new_n1156), .A4(new_n586), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT61), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1154), .A2(new_n1155), .A3(new_n1160), .A4(new_n1157), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1151), .A2(new_n1162), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1142), .A2(KEYINPUT122), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1142), .A2(KEYINPUT122), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n1158), .A3(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1167), .B2(new_n1154), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1134), .B(new_n1137), .C1(new_n1163), .C2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1135), .A2(new_n1170), .A3(G171), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1122), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1135), .A2(G171), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1170), .B(new_n1173), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1097), .B(new_n1110), .C1(new_n1172), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1096), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1109), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(G2067), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n859), .B(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(G1996), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n844), .B(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n757), .B2(new_n754), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n755), .A2(new_n758), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(G290), .A2(G1986), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT113), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(G1986), .B2(G290), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1050), .A2(new_n1062), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1190), .A2(new_n1051), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1177), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1191), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1194), .B1(new_n1179), .B2(new_n845), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT46), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1195), .B1(KEYINPUT127), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1191), .A2(new_n1180), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1196), .A2(KEYINPUT127), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1198), .B(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT47), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1184), .B(KEYINPUT126), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1203), .A2(new_n1182), .B1(G2067), .B2(new_n859), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1191), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1206), .B(KEYINPUT48), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1207), .B1(new_n1185), .B2(new_n1194), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1202), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1193), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g786(.A(new_n1036), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n1213), .B1(KEYINPUT43), .B2(new_n1034), .ZN(new_n1214));
  NOR2_X1   g788(.A1(G229), .A2(new_n461), .ZN(new_n1215));
  INV_X1    g789(.A(new_n1215), .ZN(new_n1216));
  INV_X1    g790(.A(G227), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n677), .A2(new_n1217), .ZN(new_n1218));
  NOR4_X1   g792(.A1(new_n1214), .A2(new_n932), .A3(new_n1216), .A4(new_n1218), .ZN(G308));
  INV_X1    g793(.A(new_n932), .ZN(new_n1220));
  INV_X1    g794(.A(new_n1218), .ZN(new_n1221));
  NAND4_X1  g795(.A1(new_n1220), .A2(new_n1037), .A3(new_n1215), .A4(new_n1221), .ZN(G225));
endmodule


