//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1347, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1352, new_n1353, new_n1354, new_n1355, new_n1356, new_n1357,
    new_n1358, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  OR2_X1    g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n201), .A2(G77), .A3(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(new_n202), .A2(G50), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n206), .A2(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT66), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G116), .A2(G270), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n221), .ZN(new_n224));
  INV_X1    g0024(.A(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  OAI22_X1  g0028(.A1(new_n225), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(G77), .B2(G244), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(new_n211), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT67), .B(KEYINPUT1), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n215), .B(new_n234), .C1(new_n214), .C2(new_n213), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT68), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT69), .B(G50), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT73), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n253), .B1(new_n211), .B2(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(KEYINPUT73), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(new_n207), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT24), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT82), .B(G33), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n208), .B(new_n260), .C1(new_n261), .C2(new_n259), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT22), .B1(new_n262), .B2(new_n218), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT3), .B(G33), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT88), .B(KEYINPUT22), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n264), .A2(new_n265), .A3(new_n208), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G87), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G107), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT23), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n261), .A2(new_n208), .A3(G116), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n258), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  AOI211_X1 g0076(.A(KEYINPUT24), .B(new_n274), .C1(new_n263), .C2(new_n267), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n257), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT82), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n254), .A2(KEYINPUT82), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT3), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G257), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n219), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n284), .A2(new_n260), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n261), .A2(G294), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n280), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT5), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n280), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(KEYINPUT70), .A2(G41), .ZN(new_n297));
  NOR2_X1   g0097(.A1(KEYINPUT70), .A2(G41), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT5), .ZN(new_n299));
  INV_X1    g0099(.A(G45), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT85), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT70), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(KEYINPUT70), .A2(G41), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(new_n292), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT85), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n309), .A3(new_n301), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n296), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n293), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(new_n301), .A3(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n313), .A2(G264), .A3(new_n280), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n291), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G190), .ZN(new_n316));
  INV_X1    g0116(.A(new_n257), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n254), .A2(G1), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G13), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n320), .A2(new_n208), .A3(G1), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n317), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n269), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n269), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT25), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n289), .A2(new_n290), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n279), .ZN(new_n329));
  INV_X1    g0129(.A(new_n314), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n279), .A2(new_n294), .A3(new_n293), .ZN(new_n331));
  INV_X1    g0131(.A(new_n310), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n309), .B1(new_n308), .B2(new_n301), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G200), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n278), .A2(new_n316), .A3(new_n327), .A4(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n284), .A2(new_n208), .A3(G87), .A4(new_n260), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(KEYINPUT22), .B1(new_n266), .B2(G87), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT24), .B1(new_n340), .B2(new_n274), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n268), .A2(new_n258), .A3(new_n275), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n317), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n327), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT89), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT89), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n278), .A2(new_n346), .A3(new_n327), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n315), .A2(G179), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n335), .A2(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n338), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n254), .A2(KEYINPUT82), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n281), .A2(G33), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n259), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n260), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT83), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(KEYINPUT7), .A2(G20), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT83), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n260), .C1(new_n261), .C2(new_n259), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n353), .A2(new_n354), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n356), .B1(new_n362), .B2(KEYINPUT3), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(G20), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(G68), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT74), .B(G58), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n202), .B1(new_n366), .B2(new_n227), .ZN(new_n367));
  NOR2_X1   g0167(.A1(G20), .A2(G33), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n367), .A2(G20), .B1(G159), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n365), .A2(KEYINPUT16), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n260), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n358), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n353), .A2(new_n354), .A3(new_n259), .ZN(new_n374));
  AOI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n371), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  OAI211_X1 g0176(.A(G68), .B(new_n373), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n369), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n370), .A2(new_n257), .A3(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(KEYINPUT8), .A2(G58), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT8), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n366), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n322), .ZN(new_n385));
  INV_X1    g0185(.A(G1), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n257), .B1(new_n386), .B2(G20), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(new_n387), .B2(new_n384), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n226), .A2(G1698), .ZN(new_n390));
  OR2_X1    g0190(.A1(G223), .A2(G1698), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n284), .A2(new_n260), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n280), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n386), .B1(G41), .B2(G45), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n280), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G232), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n300), .B1(new_n297), .B2(new_n298), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(new_n386), .A3(G274), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n394), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G179), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n389), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT18), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n389), .A2(KEYINPUT18), .A3(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT84), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n392), .A2(new_n393), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n401), .B1(new_n412), .B2(new_n279), .ZN(new_n413));
  INV_X1    g0213(.A(new_n398), .ZN(new_n414));
  AOI21_X1  g0214(.A(G200), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n394), .A2(new_n398), .A3(G190), .A4(new_n401), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n279), .ZN(new_n418));
  INV_X1    g0218(.A(G190), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(new_n414), .A4(new_n400), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n420), .B(KEYINPUT84), .C1(new_n402), .C2(G200), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n381), .A2(new_n388), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT17), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n410), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(G20), .B1(new_n201), .B2(new_n202), .ZN(new_n430));
  INV_X1    g0230(.A(G150), .ZN(new_n431));
  INV_X1    g0231(.A(new_n368), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n208), .A2(G33), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n430), .B1(new_n431), .B2(new_n432), .C1(new_n384), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n257), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n321), .A2(new_n225), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n387), .A2(G50), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT9), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n400), .B1(new_n396), .B2(new_n226), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT71), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(KEYINPUT72), .A2(G223), .ZN(new_n443));
  NOR2_X1   g0243(.A1(KEYINPUT72), .A2(G223), .ZN(new_n444));
  OAI21_X1  g0244(.A(G1698), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n287), .A2(G222), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n264), .A3(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(new_n279), .C1(G77), .C2(new_n264), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n440), .A2(new_n441), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n442), .A2(G190), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n440), .B(KEYINPUT71), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n453), .A2(KEYINPUT77), .A3(G190), .A4(new_n448), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n448), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n439), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT10), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n439), .A2(new_n455), .A3(KEYINPUT10), .A4(new_n457), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n438), .B1(new_n456), .B2(G179), .ZN(new_n462));
  AOI21_X1  g0262(.A(G169), .B1(new_n453), .B2(new_n448), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n226), .A2(new_n287), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n397), .A2(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n260), .A2(new_n466), .A3(new_n371), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G97), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT78), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n468), .A2(new_n472), .A3(new_n469), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n471), .A2(new_n279), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n280), .A2(G238), .A3(new_n395), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n400), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n399), .A2(KEYINPUT79), .A3(new_n386), .A4(G274), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  XOR2_X1   g0280(.A(KEYINPUT80), .B(KEYINPUT13), .Z(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n481), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n474), .A2(new_n483), .A3(new_n475), .A4(new_n479), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(KEYINPUT81), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n480), .A2(new_n486), .A3(new_n481), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(G200), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n227), .A2(G20), .ZN(new_n489));
  INV_X1    g0289(.A(G77), .ZN(new_n490));
  OAI221_X1 g0290(.A(new_n489), .B1(new_n433), .B2(new_n490), .C1(new_n432), .C2(new_n225), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n491), .A2(new_n257), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT11), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n492), .A2(KEYINPUT11), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n387), .A2(G68), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n321), .A2(new_n227), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n496), .B(KEYINPUT12), .ZN(new_n497));
  AND4_X1   g0297(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n480), .A2(KEYINPUT13), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(G190), .A3(new_n484), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n488), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n485), .A2(G169), .A3(new_n487), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT14), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n499), .A2(G179), .A3(new_n484), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT14), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n485), .A2(new_n506), .A3(G169), .A4(new_n487), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n498), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n321), .A2(new_n490), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n387), .A2(G77), .ZN(new_n512));
  XOR2_X1   g0312(.A(KEYINPUT8), .B(G58), .Z(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n368), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n208), .B2(new_n490), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT75), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g0317(.A(KEYINPUT15), .B(G87), .Z(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n208), .A3(G33), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n514), .B(KEYINPUT75), .C1(new_n208), .C2(new_n490), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n521), .A2(KEYINPUT76), .A3(new_n257), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT76), .B1(new_n521), .B2(new_n257), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n511), .B(new_n512), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n372), .B1(G232), .B2(new_n287), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n228), .B2(new_n287), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(new_n279), .C1(G107), .C2(new_n264), .ZN(new_n527));
  INV_X1    g0327(.A(G244), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n400), .C1(new_n528), .C2(new_n396), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n404), .ZN(new_n530));
  OR2_X1    g0330(.A1(new_n529), .A2(G179), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n524), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(G200), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n419), .B2(new_n529), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n524), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n429), .A2(new_n465), .A3(new_n510), .A4(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n313), .A2(G270), .A3(new_n280), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G264), .A2(G1698), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n285), .B2(G1698), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n260), .B(new_n541), .C1(new_n261), .C2(new_n259), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n372), .A2(G303), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n280), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n311), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G190), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G20), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G283), .ZN(new_n549));
  INV_X1    g0349(.A(G97), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n208), .C1(G33), .C2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n257), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT20), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n257), .A2(KEYINPUT20), .A3(new_n548), .A4(new_n551), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n322), .A2(G116), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n257), .A2(new_n318), .A3(new_n321), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(G116), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G200), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n546), .B(new_n561), .C1(new_n562), .C2(new_n545), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n545), .A2(new_n560), .A3(G179), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n545), .A2(new_n404), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(new_n560), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n313), .A2(G270), .A3(new_n280), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n542), .A2(new_n543), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n334), .B(new_n568), .C1(new_n569), .C2(new_n280), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n565), .A2(new_n570), .A3(new_n560), .A4(G169), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n563), .B(new_n564), .C1(new_n567), .C2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n313), .A2(G257), .A3(new_n280), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n334), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n260), .A2(new_n371), .A3(G250), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n287), .B1(new_n575), .B2(KEYINPUT4), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n549), .B1(new_n372), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n260), .B1(new_n261), .B2(new_n259), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n528), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n280), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(G169), .B1(new_n574), .B2(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n313), .A2(G257), .A3(new_n280), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n311), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT4), .B1(new_n363), .B2(G244), .ZN(new_n587));
  INV_X1    g0387(.A(new_n549), .ZN(new_n588));
  INV_X1    g0388(.A(new_n577), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n264), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n580), .B1(new_n264), .B2(G250), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n287), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n279), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n586), .A2(new_n593), .A3(G179), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(G107), .B(new_n373), .C1(new_n375), .C2(new_n376), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n550), .A2(new_n269), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G97), .A2(G107), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n269), .A2(KEYINPUT6), .A3(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(G20), .B1(G77), .B2(new_n368), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n257), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n322), .A2(G97), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n323), .B2(new_n550), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n595), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n604), .B2(new_n257), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n574), .A2(new_n583), .A3(G190), .ZN(new_n613));
  AOI21_X1  g0413(.A(G200), .B1(new_n586), .B2(new_n593), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n572), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT86), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n228), .A2(new_n287), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n528), .A2(G1698), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n355), .A2(new_n356), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n261), .A2(G116), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n618), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(KEYINPUT86), .B(new_n623), .C1(new_n581), .C2(new_n621), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n279), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n279), .B1(new_n294), .B2(new_n301), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(G250), .B2(new_n301), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(G200), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT19), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(new_n208), .A3(G33), .A4(G97), .ZN(new_n633));
  NOR2_X1   g0433(.A1(G87), .A2(G97), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n269), .B1(new_n469), .B2(new_n208), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(new_n632), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n262), .B2(new_n227), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n257), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n322), .B2(new_n518), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n323), .A2(new_n218), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n631), .A2(KEYINPUT87), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT87), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n562), .B1(new_n627), .B2(new_n629), .ZN(new_n644));
  OAI221_X1 g0444(.A(new_n638), .B1(new_n218), .B2(new_n323), .C1(new_n322), .C2(new_n518), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n627), .A2(G190), .A3(new_n629), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n642), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n518), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n323), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n639), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n404), .B1(new_n627), .B2(new_n629), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n627), .A2(G179), .A3(new_n629), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n352), .A2(new_n538), .A3(new_n617), .A4(new_n655), .ZN(G372));
  INV_X1    g0456(.A(new_n464), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n508), .A2(new_n509), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT93), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n532), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n524), .A2(KEYINPUT93), .A3(new_n530), .A4(new_n531), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n427), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT17), .B1(new_n422), .B2(new_n423), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n665), .A3(new_n501), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n410), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n460), .A2(new_n461), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n657), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT91), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT90), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n653), .A2(new_n652), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n630), .A2(G169), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n627), .A2(G179), .A3(new_n629), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT90), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n651), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n644), .A2(new_n645), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n647), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n337), .A2(new_n611), .A3(new_n615), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n670), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n564), .B1(new_n567), .B2(new_n571), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n278), .A2(new_n327), .B1(new_n350), .B2(new_n349), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n671), .B1(new_n653), .B2(new_n652), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n673), .A2(KEYINPUT90), .A3(new_n674), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n687), .A2(new_n651), .B1(new_n647), .B2(new_n677), .ZN(new_n688));
  INV_X1    g0488(.A(new_n680), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(KEYINPUT91), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n681), .A2(new_n684), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n612), .B1(new_n584), .B2(new_n594), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n648), .A2(new_n692), .A3(new_n654), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT26), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n584), .A2(KEYINPUT92), .A3(new_n594), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT92), .B1(new_n584), .B2(new_n594), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n696), .A2(new_n697), .A3(new_n612), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT26), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n676), .A2(new_n698), .A3(new_n699), .A4(new_n678), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n694), .A2(new_n700), .A3(new_n676), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n691), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n669), .B1(new_n537), .B2(new_n702), .ZN(G369));
  INV_X1    g0503(.A(new_n564), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n566), .A2(new_n565), .A3(new_n560), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n570), .A2(new_n560), .A3(G169), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT21), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n704), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n320), .A2(G20), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n386), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G343), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n708), .B(new_n563), .C1(new_n561), .C2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n682), .A2(new_n560), .A3(new_n715), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n348), .A2(new_n715), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n345), .A2(new_n347), .B1(new_n350), .B2(new_n349), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n352), .A2(new_n721), .B1(new_n722), .B2(new_n715), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n683), .A2(new_n716), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n343), .A2(KEYINPUT89), .A3(new_n344), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n346), .B1(new_n278), .B2(new_n327), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n351), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n721), .A2(new_n730), .A3(new_n337), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(new_n715), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT94), .B1(new_n708), .B2(new_n715), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT94), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n682), .A2(new_n735), .A3(new_n716), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n727), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n725), .A2(new_n738), .ZN(G399));
  NAND2_X1  g0539(.A1(new_n306), .A2(new_n307), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n212), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n634), .A2(new_n269), .A3(new_n547), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n743), .A2(new_n386), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT95), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  INV_X1    g0548(.A(new_n743), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n747), .B(new_n748), .C1(new_n205), .C2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  INV_X1    g0551(.A(G330), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n352), .A2(new_n655), .A3(new_n617), .A4(new_n716), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT31), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n315), .A2(G179), .A3(new_n629), .A4(new_n627), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n539), .A2(new_n544), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n586), .A2(new_n593), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(KEYINPUT30), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n586), .A2(new_n593), .A3(new_n756), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT30), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n653), .A2(new_n759), .A3(new_n760), .A4(new_n315), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT96), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n315), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n586), .A2(new_n593), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n764), .A2(new_n765), .A3(new_n570), .A4(new_n630), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n762), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n762), .B2(new_n766), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n715), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n754), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n674), .A2(new_n335), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n760), .B1(new_n772), .B2(new_n759), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n674), .A2(new_n757), .A3(KEYINPUT30), .A4(new_n335), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n766), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(KEYINPUT31), .A3(new_n715), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n752), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n730), .A2(new_n708), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n586), .A2(new_n593), .A3(new_n419), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n562), .B1(new_n574), .B2(new_n583), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n610), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(KEYINPUT98), .B1(new_n782), .B2(new_n692), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT98), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n611), .A2(new_n615), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n338), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n779), .A2(new_n786), .A3(new_n688), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n648), .A2(new_n699), .A3(new_n692), .A4(new_n654), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n788), .A2(new_n676), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n676), .A2(new_n698), .A3(new_n678), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT26), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n787), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(KEYINPUT29), .A3(new_n716), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n715), .B1(new_n691), .B2(new_n701), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n778), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n751), .B1(new_n798), .B2(G1), .ZN(G364));
  NAND2_X1  g0599(.A1(new_n709), .A2(G45), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT99), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(KEYINPUT99), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n801), .A2(G1), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n749), .ZN(new_n805));
  AND3_X1   g0605(.A1(KEYINPUT100), .A2(G20), .A3(G179), .ZN(new_n806));
  AOI21_X1  g0606(.A(KEYINPUT100), .B1(G20), .B2(G179), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n809), .A2(new_n419), .A3(new_n562), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n419), .A2(G200), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n811), .A2(new_n225), .B1(new_n814), .B2(new_n366), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n808), .A2(new_n419), .A3(G200), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n815), .B1(G68), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n208), .A2(G179), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n819), .A2(G190), .A3(G200), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n264), .B1(new_n820), .B2(new_n218), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G190), .A2(G200), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n824));
  INV_X1    g0624(.A(G159), .ZN(new_n825));
  OR3_X1    g0625(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n819), .A2(new_n419), .A3(G200), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G107), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n826), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G179), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n812), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G20), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n821), .B(new_n831), .C1(G97), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n808), .A2(new_n822), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n818), .B(new_n835), .C1(new_n490), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT102), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n264), .B1(new_n834), .B2(G294), .ZN(new_n839));
  INV_X1    g0639(.A(new_n823), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G329), .ZN(new_n841));
  INV_X1    g0641(.A(G303), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n839), .B(new_n841), .C1(new_n842), .C2(new_n820), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G322), .B2(new_n813), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n810), .A2(G326), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n828), .A2(G283), .ZN(new_n846));
  XOR2_X1   g0646(.A(KEYINPUT33), .B(G317), .Z(new_n847));
  INV_X1    g0647(.A(G311), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n816), .A2(new_n847), .B1(new_n836), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n838), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n207), .B1(G20), .B2(new_n404), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n805), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n264), .A2(G355), .A3(new_n212), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n357), .A2(new_n360), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(new_n742), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n248), .B2(new_n300), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n206), .A2(G45), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n855), .B1(G116), .B2(new_n212), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(G13), .A2(G33), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(G20), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(new_n853), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n863), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n854), .B(new_n865), .C1(new_n719), .C2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n719), .A2(G330), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n720), .A2(new_n805), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(G396));
  NAND2_X1  g0670(.A1(new_n524), .A2(new_n715), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n535), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n871), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n660), .A2(new_n661), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n794), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n874), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n715), .B(new_n877), .C1(new_n691), .C2(new_n701), .ZN(new_n878));
  OR3_X1    g0678(.A1(new_n778), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n778), .B1(new_n876), .B2(new_n878), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n805), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n828), .A2(G68), .ZN(new_n882));
  INV_X1    g0682(.A(G132), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(new_n823), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n834), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n885), .B(new_n856), .C1(new_n366), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n813), .A2(G143), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n431), .B2(new_n816), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(G137), .B2(new_n810), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n825), .B2(new_n836), .ZN(new_n891));
  XNOR2_X1  g0691(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n893), .B1(new_n225), .B2(new_n820), .C1(new_n892), .C2(new_n891), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n827), .A2(new_n218), .ZN(new_n895));
  INV_X1    g0695(.A(new_n820), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(G107), .B2(new_n896), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n897), .B1(new_n848), .B2(new_n823), .C1(new_n836), .C2(new_n547), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n372), .B1(new_n886), .B2(new_n550), .ZN(new_n899));
  INV_X1    g0699(.A(G294), .ZN(new_n900));
  XNOR2_X1  g0700(.A(KEYINPUT103), .B(G283), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n814), .A2(new_n900), .B1(new_n816), .B2(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n842), .B2(new_n811), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n894), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n805), .B1(new_n906), .B2(new_n853), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n853), .A2(new_n861), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n907), .B1(G77), .B2(new_n909), .C1(new_n875), .C2(new_n862), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n881), .A2(new_n910), .ZN(G384));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n365), .A2(new_n369), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n379), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n257), .A3(new_n370), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n713), .B1(new_n915), .B2(new_n388), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n665), .B2(new_n410), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n389), .B1(new_n417), .B2(new_n421), .ZN(new_n919));
  NOR4_X1   g0719(.A1(new_n394), .A2(new_n398), .A3(new_n832), .A4(new_n401), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n413), .A2(new_n414), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(G169), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n388), .A2(new_n915), .B1(new_n922), .B2(new_n713), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT37), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT37), .ZN(new_n925));
  INV_X1    g0725(.A(new_n713), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n389), .B1(new_n405), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n424), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n912), .B1(new_n918), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n426), .A2(new_n427), .ZN(new_n932));
  INV_X1    g0732(.A(new_n409), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT18), .B1(new_n389), .B2(new_n405), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n916), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(KEYINPUT38), .A3(new_n929), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n762), .A2(new_n763), .A3(new_n766), .ZN(new_n940));
  AND4_X1   g0740(.A1(KEYINPUT31), .A2(new_n939), .A3(new_n715), .A4(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n771), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n509), .A2(new_n715), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n658), .A2(new_n501), .A3(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n509), .B(new_n715), .C1(new_n508), .C2(new_n502), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n938), .A2(new_n943), .A3(new_n875), .A4(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n941), .B1(new_n754), .B2(new_n770), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n945), .A2(new_n946), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n950), .A2(new_n877), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n389), .A2(new_n926), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n665), .B2(new_n410), .ZN(new_n954));
  INV_X1    g0754(.A(new_n928), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n925), .B1(new_n424), .B2(new_n927), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n912), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n949), .B1(new_n958), .B2(new_n937), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n948), .A2(new_n949), .B1(new_n952), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT105), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n950), .A2(new_n537), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n961), .B(new_n962), .Z(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(G330), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n532), .A2(new_n715), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n938), .B(new_n947), .C1(new_n878), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n410), .A2(new_n926), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT39), .ZN(new_n969));
  AOI221_X4 g0769(.A(new_n912), .B1(new_n924), .B2(new_n928), .C1(new_n428), .C2(new_n916), .ZN(new_n970));
  INV_X1    g0770(.A(new_n953), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n428), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n956), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n928), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT38), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n969), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n658), .A2(new_n715), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n931), .A2(new_n937), .A3(KEYINPUT39), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n966), .A2(new_n968), .A3(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n538), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n669), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n980), .B(new_n982), .Z(new_n983));
  XNOR2_X1  g0783(.A(new_n964), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n386), .B2(new_n709), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n547), .B1(new_n602), .B2(KEYINPUT35), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(new_n209), .C1(KEYINPUT35), .C2(new_n602), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT36), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n366), .A2(new_n227), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n989), .A2(new_n490), .A3(new_n205), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n201), .A2(new_n227), .ZN(new_n991));
  OAI211_X1 g0791(.A(G1), .B(new_n320), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n985), .A2(new_n988), .A3(new_n992), .ZN(G367));
  NAND2_X1  g0793(.A1(new_n645), .A2(new_n715), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n676), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n688), .B2(new_n994), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n783), .A2(new_n785), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n612), .A2(new_n716), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT106), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT106), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1004), .B(new_n1001), .C1(new_n783), .C2(new_n785), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n698), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n1003), .A2(new_n1005), .B1(new_n1006), .B2(new_n716), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n724), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1006), .A2(new_n716), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n782), .A2(new_n692), .A3(KEYINPUT98), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n784), .B1(new_n611), .B2(new_n615), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1002), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n1004), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1000), .A2(KEYINPUT106), .A3(new_n1002), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n733), .A2(new_n737), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n1015), .A2(new_n1016), .A3(KEYINPUT42), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT42), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n692), .B1(new_n1007), .B2(new_n722), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1017), .B(new_n1018), .C1(new_n715), .C2(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n996), .A2(new_n997), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1008), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1020), .A2(new_n1008), .A3(new_n1021), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n999), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AND3_X1   g0825(.A1(new_n1020), .A2(new_n1008), .A3(new_n1021), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1026), .A2(new_n1022), .A3(new_n998), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n743), .B(KEYINPUT41), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n734), .A2(new_n736), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n726), .B1(new_n723), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(KEYINPUT107), .B1(new_n1032), .B2(new_n1015), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT107), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n738), .A2(new_n1034), .A3(new_n1007), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1035), .A3(KEYINPUT45), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT44), .B1(new_n738), .B2(new_n1007), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n738), .A2(new_n1007), .A3(KEYINPUT44), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT45), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1032), .A2(new_n1015), .A3(KEYINPUT107), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1034), .B1(new_n738), .B2(new_n1007), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n725), .A3(new_n1039), .A4(new_n1043), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1043), .A2(new_n1039), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n724), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n720), .B(new_n723), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(new_n1031), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n797), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1044), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1030), .B1(new_n1050), .B2(new_n798), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1028), .B1(new_n1051), .B2(new_n803), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n814), .A2(new_n431), .B1(new_n825), .B2(new_n816), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n827), .A2(new_n490), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G68), .B2(new_n834), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n264), .C1(new_n366), .C2(new_n820), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G143), .B2(new_n810), .ZN(new_n1057));
  INV_X1    g0857(.A(G137), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n823), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n836), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1053), .B(new_n1059), .C1(new_n201), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n840), .A2(G317), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n810), .A2(G311), .B1(new_n817), .B2(G294), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n836), .B2(new_n902), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n856), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n842), .B2(new_n814), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n827), .A2(new_n550), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G107), .B2(new_n834), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n896), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT46), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n820), .B2(new_n547), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1064), .A2(new_n1066), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1061), .B1(new_n1062), .B2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT47), .Z(new_n1075));
  AOI21_X1  g0875(.A(new_n805), .B1(new_n1075), .B2(new_n853), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n857), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n864), .B1(new_n212), .B2(new_n649), .C1(new_n243), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n996), .A2(new_n863), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1052), .A2(new_n1080), .ZN(G387));
  NOR2_X1   g0881(.A1(new_n733), .A2(new_n866), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n813), .A2(G317), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n842), .B2(new_n836), .C1(new_n848), .C2(new_n816), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G322), .B2(new_n810), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT48), .Z(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n900), .B2(new_n820), .C1(new_n886), .C2(new_n902), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT49), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n828), .A2(G116), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n856), .B1(G326), .B2(new_n840), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n816), .A2(new_n384), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n811), .A2(new_n825), .B1(new_n814), .B2(new_n225), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n886), .A2(new_n649), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1067), .B(new_n1097), .C1(G150), .C2(new_n840), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n820), .A2(new_n490), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1065), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1060), .A2(G68), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1093), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n805), .B(new_n1082), .C1(new_n1103), .C2(new_n853), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n513), .A2(new_n225), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n744), .B1(new_n1105), .B2(KEYINPUT50), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n300), .C1(KEYINPUT50), .C2(new_n1105), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G68), .B2(G77), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n857), .B1(new_n239), .B2(new_n300), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n264), .A2(new_n744), .A3(new_n212), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n212), .A2(G107), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n864), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1104), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1049), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n743), .B(KEYINPUT108), .Z(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1048), .A2(new_n797), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1114), .B1(new_n804), .B2(new_n1048), .C1(new_n1118), .C2(new_n1119), .ZN(G393));
  NAND3_X1  g0920(.A1(new_n1044), .A2(new_n1046), .A3(new_n803), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n896), .A2(new_n901), .B1(new_n834), .B2(G116), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n840), .A2(G322), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(new_n842), .C2(new_n816), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n264), .B(new_n1124), .C1(G294), .C2(new_n1060), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n810), .A2(G317), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n848), .B2(new_n814), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1125), .A2(new_n829), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT111), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n811), .A2(new_n431), .B1(new_n814), .B2(new_n825), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT51), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n896), .A2(G68), .B1(new_n840), .B2(G143), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT109), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n895), .B(new_n1065), .C1(G77), .C2(new_n834), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n201), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1136), .A2(KEYINPUT109), .B1(new_n1139), .B2(new_n816), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n513), .B2(new_n1060), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1133), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT112), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n805), .B1(new_n1144), .B2(new_n853), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n864), .B1(new_n550), .B2(new_n212), .C1(new_n1077), .C2(new_n251), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1015), .A2(new_n863), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT113), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(new_n1115), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1117), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1049), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1050), .B1(new_n1153), .B2(new_n1150), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1121), .B(new_n1148), .C1(new_n1152), .C2(new_n1154), .ZN(G390));
  NAND2_X1  g0955(.A1(new_n962), .A2(G330), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT117), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n950), .A2(KEYINPUT117), .A3(new_n537), .A4(new_n752), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n982), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(KEYINPUT31), .A2(new_n753), .B1(new_n769), .B2(new_n715), .ZN(new_n1161));
  OAI211_X1 g0961(.A(G330), .B(new_n875), .C1(new_n1161), .C2(new_n941), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT114), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n947), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n945), .A2(KEYINPUT114), .A3(new_n946), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n792), .A2(new_n716), .A3(new_n875), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n965), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT116), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n777), .A2(new_n1172), .A3(new_n875), .A4(new_n947), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n776), .ZN(new_n1174));
  OAI211_X1 g0974(.A(G330), .B(new_n875), .C1(new_n1161), .C2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(KEYINPUT116), .B1(new_n1175), .B2(new_n951), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1171), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n965), .B1(new_n794), .B2(new_n875), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n877), .B1(new_n771), .B2(new_n942), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(G330), .A3(new_n947), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n951), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1160), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n976), .A2(new_n978), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n794), .A2(new_n875), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n951), .B1(new_n1185), .B2(new_n1169), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1186), .B2(new_n977), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n1165), .A3(new_n1164), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT115), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n977), .B1(new_n958), .B2(new_n937), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1190), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1187), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1180), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1176), .A2(new_n1173), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n1187), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1183), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT118), .B1(new_n1198), .B2(new_n1116), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1191), .B1(new_n1170), .B2(new_n1166), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT115), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1178), .A2(new_n951), .B1(new_n658), .B2(new_n715), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1201), .A2(new_n1202), .B1(new_n1184), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1180), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1197), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT117), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n962), .B2(G330), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n669), .B(new_n981), .C1(new_n1208), .C2(new_n1158), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1182), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1176), .A2(new_n1173), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1188), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1209), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1206), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT118), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1117), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1195), .A2(new_n1183), .A3(new_n1197), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1199), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n853), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n816), .A2(new_n1058), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n820), .A2(new_n431), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT53), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n372), .B1(new_n828), .B2(new_n201), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n825), .C2(new_n886), .ZN(new_n1225));
  XOR2_X1   g1025(.A(KEYINPUT54), .B(G143), .Z(new_n1226));
  AOI211_X1 g1026(.A(new_n1221), .B(new_n1225), .C1(new_n1060), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n840), .A2(G125), .ZN(new_n1228));
  INV_X1    g1028(.A(G128), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n811), .A2(new_n1229), .B1(new_n814), .B2(new_n883), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT120), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1227), .A2(new_n1228), .A3(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n882), .B1(new_n900), .B2(new_n823), .C1(new_n886), .C2(new_n490), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G283), .B2(new_n810), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n814), .A2(new_n547), .B1(new_n269), .B2(new_n816), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1060), .A2(G97), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n264), .B1(new_n896), .B2(G87), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1234), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1220), .B1(new_n1232), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n805), .B1(new_n384), .B2(new_n908), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT119), .Z(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(new_n1184), .C2(new_n861), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1206), .B2(new_n803), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1219), .A2(new_n1244), .ZN(G378));
  INV_X1    g1045(.A(KEYINPUT57), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1209), .B1(new_n1206), .B2(new_n1214), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n875), .B(new_n947), .C1(new_n1161), .C2(new_n941), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT38), .B1(new_n936), .B2(new_n929), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n970), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n949), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n959), .A2(new_n1179), .A3(new_n947), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(G330), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1253), .A2(new_n968), .A3(new_n966), .A4(new_n979), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n980), .A2(new_n960), .A3(G330), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT55), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n465), .B(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n438), .A2(new_n926), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n465), .B(KEYINPUT55), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(new_n1258), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1264), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1254), .A2(new_n1255), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1246), .B1(new_n1247), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1268), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1254), .A2(new_n1255), .A3(new_n1268), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1277), .B(KEYINPUT57), .C1(new_n1198), .C2(new_n1209), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1272), .A2(new_n1278), .A3(new_n1117), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1268), .A2(new_n861), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n908), .A2(new_n1139), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n814), .A2(new_n1229), .B1(new_n883), .B2(new_n816), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1060), .A2(G137), .B1(new_n896), .B2(new_n1226), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(new_n431), .C2(new_n886), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(G125), .B2(new_n810), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1287), .A2(KEYINPUT59), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n840), .A2(G124), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(KEYINPUT59), .ZN(new_n1290));
  AOI211_X1 g1090(.A(G33), .B(G41), .C1(new_n828), .C2(G159), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  OAI221_X1 g1092(.A(new_n225), .B1(G33), .B2(G41), .C1(new_n856), .C2(new_n741), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n811), .A2(new_n547), .ZN(new_n1294));
  INV_X1    g1094(.A(G283), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n886), .A2(new_n227), .B1(new_n1295), .B2(new_n823), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n827), .A2(new_n366), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(new_n1294), .A2(new_n1099), .A3(new_n1296), .A4(new_n1297), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n814), .A2(new_n269), .B1(new_n550), .B2(new_n816), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n518), .B2(new_n1060), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1298), .A2(new_n740), .A3(new_n1065), .A4(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT58), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1292), .A2(new_n1293), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n805), .B1(new_n1303), .B2(new_n853), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1280), .A2(new_n1281), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1277), .B2(new_n803), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1279), .A2(KEYINPUT122), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT122), .B1(new_n1279), .B2(new_n1307), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(G375));
  NAND3_X1  g1111(.A1(new_n1213), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1183), .A2(new_n1029), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n804), .B1(new_n1213), .B2(new_n1210), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n908), .A2(new_n227), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n862), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1097), .B1(G97), .B2(new_n896), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n842), .B2(new_n823), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n816), .A2(new_n547), .ZN(new_n1319));
  NOR4_X1   g1119(.A1(new_n1318), .A2(new_n1319), .A3(new_n264), .A4(new_n1054), .ZN(new_n1320));
  OAI22_X1  g1120(.A1(new_n811), .A2(new_n900), .B1(new_n836), .B2(new_n269), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1320), .B(new_n1322), .C1(new_n1295), .C2(new_n814), .ZN(new_n1323));
  XOR2_X1   g1123(.A(new_n1323), .B(KEYINPUT123), .Z(new_n1324));
  OAI22_X1  g1124(.A1(new_n811), .A2(new_n883), .B1(new_n814), .B2(new_n1058), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1325), .B1(new_n817), .B2(new_n1226), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1060), .A2(G150), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1065), .B1(G50), .B2(new_n834), .ZN(new_n1328));
  OAI22_X1  g1128(.A1(new_n820), .A2(new_n825), .B1(new_n823), .B2(new_n1229), .ZN(new_n1329));
  XOR2_X1   g1129(.A(new_n1329), .B(KEYINPUT124), .Z(new_n1330));
  NOR2_X1   g1130(.A1(new_n1330), .A2(new_n1297), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1326), .A2(new_n1327), .A3(new_n1328), .A4(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1220), .B1(new_n1324), .B2(new_n1332), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1316), .A2(new_n805), .A3(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1314), .B1(new_n1315), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1313), .A2(new_n1335), .ZN(G381));
  NOR3_X1   g1136(.A1(new_n1308), .A2(new_n1309), .A3(G378), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1148), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1154), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1116), .B1(new_n1153), .B2(new_n1150), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1338), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1341), .A2(new_n1080), .A3(new_n1052), .A4(new_n1121), .ZN(new_n1342));
  OR2_X1    g1142(.A1(G393), .A2(G396), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(G381), .A2(G384), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1337), .A2(new_n1344), .A3(new_n1345), .ZN(G407));
  AND3_X1   g1146(.A1(new_n1337), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1279), .A2(new_n1307), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT122), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  AND2_X1   g1150(.A1(new_n1219), .A2(new_n1244), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1279), .A2(KEYINPUT122), .A3(new_n1307), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1350), .A2(new_n1351), .A3(new_n1352), .ZN(new_n1353));
  OAI21_X1  g1153(.A(G213), .B1(new_n1353), .B2(G343), .ZN(new_n1354));
  OAI21_X1  g1154(.A(KEYINPUT125), .B1(new_n1347), .B2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1354), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT125), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1356), .A2(G407), .A3(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1358), .ZN(G409));
  NAND2_X1  g1159(.A1(new_n1348), .A2(G378), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n714), .A2(G213), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1277), .B(new_n1029), .C1(new_n1198), .C2(new_n1209), .ZN(new_n1362));
  NAND4_X1  g1162(.A1(new_n1219), .A2(new_n1244), .A3(new_n1307), .A4(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT60), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1312), .A2(new_n1364), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1213), .A2(new_n1209), .A3(new_n1210), .A4(KEYINPUT60), .ZN(new_n1366));
  NAND4_X1  g1166(.A1(new_n1365), .A2(new_n1117), .A3(new_n1183), .A4(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(new_n1335), .ZN(new_n1368));
  INV_X1    g1168(.A(G384), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1368), .A2(new_n1369), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1370), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1367), .A2(G384), .A3(new_n1335), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1372), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1371), .A2(new_n1373), .ZN(new_n1374));
  NAND4_X1  g1174(.A1(new_n1360), .A2(new_n1361), .A3(new_n1363), .A4(new_n1374), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1375), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1363), .A2(new_n1361), .ZN(new_n1377));
  AOI22_X1  g1177(.A1(new_n1279), .A2(new_n1307), .B1(new_n1219), .B2(new_n1244), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1380));
  OR2_X1    g1180(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1381));
  NAND4_X1  g1181(.A1(new_n1379), .A2(new_n1374), .A3(new_n1380), .A4(new_n1381), .ZN(new_n1382));
  INV_X1    g1182(.A(new_n1307), .ZN(new_n1383));
  OAI21_X1  g1183(.A(new_n1277), .B1(new_n1198), .B2(new_n1209), .ZN(new_n1384));
  AOI21_X1  g1184(.A(new_n1116), .B1(new_n1384), .B2(new_n1246), .ZN(new_n1385));
  AOI21_X1  g1185(.A(new_n1383), .B1(new_n1385), .B2(new_n1278), .ZN(new_n1386));
  OAI211_X1 g1186(.A(new_n1361), .B(new_n1363), .C1(new_n1386), .C2(new_n1351), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n714), .A2(G213), .A3(G2897), .ZN(new_n1388));
  AND3_X1   g1188(.A1(new_n1370), .A2(new_n1372), .A3(new_n1388), .ZN(new_n1389));
  AOI21_X1  g1189(.A(new_n1388), .B1(new_n1370), .B2(new_n1372), .ZN(new_n1390));
  NOR2_X1   g1190(.A1(new_n1389), .A2(new_n1390), .ZN(new_n1391));
  AOI21_X1  g1191(.A(KEYINPUT61), .B1(new_n1387), .B2(new_n1391), .ZN(new_n1392));
  NAND3_X1  g1192(.A1(new_n1376), .A2(new_n1382), .A3(new_n1392), .ZN(new_n1393));
  XNOR2_X1  g1193(.A(G393), .B(G396), .ZN(new_n1394));
  INV_X1    g1194(.A(new_n1394), .ZN(new_n1395));
  AND2_X1   g1195(.A1(G387), .A2(G390), .ZN(new_n1396));
  NOR2_X1   g1196(.A1(G387), .A2(G390), .ZN(new_n1397));
  OAI21_X1  g1197(.A(new_n1395), .B1(new_n1396), .B2(new_n1397), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(G387), .A2(G390), .ZN(new_n1399));
  NAND3_X1  g1199(.A1(new_n1342), .A2(new_n1394), .A3(new_n1399), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1398), .A2(new_n1400), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1393), .A2(new_n1401), .ZN(new_n1402));
  INV_X1    g1202(.A(KEYINPUT61), .ZN(new_n1403));
  NAND3_X1  g1203(.A1(new_n1398), .A2(new_n1403), .A3(new_n1400), .ZN(new_n1404));
  XNOR2_X1  g1204(.A(new_n1404), .B(KEYINPUT126), .ZN(new_n1405));
  OAI21_X1  g1205(.A(new_n1391), .B1(new_n1377), .B2(new_n1378), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1406), .A2(KEYINPUT63), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(new_n1407), .A2(new_n1375), .ZN(new_n1408));
  NAND3_X1  g1208(.A1(new_n1379), .A2(KEYINPUT63), .A3(new_n1374), .ZN(new_n1409));
  NAND3_X1  g1209(.A1(new_n1405), .A2(new_n1408), .A3(new_n1409), .ZN(new_n1410));
  NAND2_X1  g1210(.A1(new_n1402), .A2(new_n1410), .ZN(G405));
  AND3_X1   g1211(.A1(new_n1353), .A2(new_n1401), .A3(new_n1360), .ZN(new_n1412));
  AOI21_X1  g1212(.A(new_n1401), .B1(new_n1353), .B2(new_n1360), .ZN(new_n1413));
  INV_X1    g1213(.A(new_n1374), .ZN(new_n1414));
  NOR3_X1   g1214(.A1(new_n1412), .A2(new_n1413), .A3(new_n1414), .ZN(new_n1415));
  INV_X1    g1215(.A(new_n1401), .ZN(new_n1416));
  OAI21_X1  g1216(.A(new_n1416), .B1(new_n1337), .B2(new_n1378), .ZN(new_n1417));
  NAND3_X1  g1217(.A1(new_n1353), .A2(new_n1401), .A3(new_n1360), .ZN(new_n1418));
  AOI21_X1  g1218(.A(new_n1374), .B1(new_n1417), .B2(new_n1418), .ZN(new_n1419));
  NOR2_X1   g1219(.A1(new_n1415), .A2(new_n1419), .ZN(G402));
endmodule


