

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759;

  INV_X1 U368 ( .A(G953), .ZN(n750) );
  OR2_X2 U369 ( .A1(n758), .A2(n577), .ZN(n378) );
  XNOR2_X2 U370 ( .A(n550), .B(KEYINPUT32), .ZN(n758) );
  NAND2_X2 U371 ( .A1(n582), .A2(n508), .ZN(n436) );
  AND2_X2 U372 ( .A1(n555), .A2(n695), .ZN(n562) );
  XNOR2_X2 U373 ( .A(n433), .B(n362), .ZN(n757) );
  NAND2_X1 U374 ( .A1(n692), .A2(n691), .ZN(n689) );
  NAND2_X1 U375 ( .A1(n555), .A2(n599), .ZN(n556) );
  INV_X1 U376 ( .A(n585), .ZN(n692) );
  XNOR2_X1 U377 ( .A(KEYINPUT69), .B(KEYINPUT94), .ZN(n412) );
  AND2_X1 U378 ( .A1(n415), .A2(KEYINPUT89), .ZN(n401) );
  XNOR2_X1 U379 ( .A(n386), .B(KEYINPUT110), .ZN(n576) );
  NAND2_X1 U380 ( .A1(n435), .A2(n434), .ZN(n433) );
  AND2_X1 U381 ( .A1(n417), .A2(n416), .ZN(n419) );
  NOR2_X1 U382 ( .A1(n623), .A2(n620), .ZN(n603) );
  NAND2_X1 U383 ( .A1(n426), .A2(n425), .ZN(n424) );
  AND2_X1 U384 ( .A1(n369), .A2(n368), .ZN(n367) );
  XNOR2_X1 U385 ( .A(n695), .B(n398), .ZN(n599) );
  XNOR2_X1 U386 ( .A(n468), .B(n388), .ZN(n585) );
  XNOR2_X1 U387 ( .A(n657), .B(KEYINPUT59), .ZN(n658) );
  XNOR2_X1 U388 ( .A(n411), .B(n409), .ZN(n497) );
  XNOR2_X1 U389 ( .A(n413), .B(n412), .ZN(n411) );
  XNOR2_X1 U390 ( .A(n410), .B(n414), .ZN(n409) );
  XNOR2_X1 U391 ( .A(G113), .B(G119), .ZN(n413) );
  XNOR2_X1 U392 ( .A(G101), .B(KEYINPUT3), .ZN(n410) );
  NOR2_X1 U393 ( .A1(n655), .A2(n732), .ZN(n656) );
  NOR2_X1 U394 ( .A1(n647), .A2(n732), .ZN(n649) );
  NOR2_X1 U395 ( .A1(n660), .A2(n732), .ZN(n661) );
  XNOR2_X2 U396 ( .A(n562), .B(KEYINPUT104), .ZN(n702) );
  XNOR2_X2 U397 ( .A(n375), .B(n579), .ZN(n735) );
  XNOR2_X2 U398 ( .A(n526), .B(KEYINPUT4), .ZN(n498) );
  XNOR2_X1 U399 ( .A(n377), .B(n376), .ZN(n415) );
  INV_X1 U400 ( .A(KEYINPUT66), .ZN(n376) );
  NAND2_X1 U401 ( .A1(n379), .A2(n378), .ZN(n377) );
  NAND2_X1 U402 ( .A1(n441), .A2(n440), .ZN(n578) );
  XNOR2_X1 U403 ( .A(n387), .B(KEYINPUT90), .ZN(n441) );
  OR2_X1 U404 ( .A1(G237), .A2(G902), .ZN(n502) );
  NOR2_X1 U405 ( .A1(G237), .A2(G953), .ZN(n445) );
  XNOR2_X1 U406 ( .A(G137), .B(G134), .ZN(n443) );
  XNOR2_X1 U407 ( .A(G131), .B(KEYINPUT68), .ZN(n442) );
  XOR2_X1 U408 ( .A(G146), .B(G125), .Z(n487) );
  XOR2_X1 U409 ( .A(KEYINPUT17), .B(KEYINPUT95), .Z(n489) );
  INV_X1 U410 ( .A(G116), .ZN(n414) );
  OR2_X1 U411 ( .A1(n415), .A2(KEYINPUT89), .ZN(n403) );
  INV_X1 U412 ( .A(KEYINPUT67), .ZN(n385) );
  NAND2_X1 U413 ( .A1(n578), .A2(n407), .ZN(n406) );
  NAND2_X1 U414 ( .A1(n588), .A2(KEYINPUT30), .ZN(n369) );
  XNOR2_X1 U415 ( .A(G113), .B(G143), .ZN(n512) );
  XOR2_X1 U416 ( .A(G104), .B(G122), .Z(n513) );
  XNOR2_X1 U417 ( .A(n557), .B(n361), .ZN(n435) );
  AND2_X1 U418 ( .A1(n422), .A2(n421), .ZN(n420) );
  XNOR2_X1 U419 ( .A(n467), .B(n389), .ZN(n388) );
  INV_X1 U420 ( .A(KEYINPUT25), .ZN(n389) );
  OR2_X1 U421 ( .A1(n553), .A2(n552), .ZN(n386) );
  INV_X1 U422 ( .A(KEYINPUT6), .ZN(n398) );
  XNOR2_X1 U423 ( .A(n637), .B(n636), .ZN(n732) );
  NAND2_X1 U424 ( .A1(n373), .A2(KEYINPUT2), .ZN(n629) );
  AND2_X1 U425 ( .A1(n749), .A2(n408), .ZN(n392) );
  NAND2_X1 U426 ( .A1(n395), .A2(n351), .ZN(n394) );
  INV_X1 U427 ( .A(n576), .ZN(n380) );
  NAND2_X1 U428 ( .A1(n543), .A2(n431), .ZN(n429) );
  NAND2_X1 U429 ( .A1(G234), .A2(G237), .ZN(n472) );
  AND2_X1 U430 ( .A1(n544), .A2(n545), .ZN(n423) );
  NAND2_X1 U431 ( .A1(n712), .A2(KEYINPUT30), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n504), .B(n503), .ZN(n505) );
  INV_X1 U433 ( .A(G902), .ZN(n530) );
  XNOR2_X1 U434 ( .A(G472), .B(KEYINPUT72), .ZN(n450) );
  XNOR2_X1 U435 ( .A(G116), .B(G134), .ZN(n519) );
  XOR2_X1 U436 ( .A(G107), .B(G122), .Z(n520) );
  XNOR2_X1 U437 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U438 ( .A(n487), .B(n439), .ZN(n491) );
  XNOR2_X1 U439 ( .A(KEYINPUT80), .B(KEYINPUT18), .ZN(n488) );
  XNOR2_X1 U440 ( .A(n497), .B(n496), .ZN(n739) );
  XNOR2_X1 U441 ( .A(KEYINPUT73), .B(G122), .ZN(n494) );
  XOR2_X1 U442 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n495) );
  XNOR2_X1 U443 ( .A(n463), .B(KEYINPUT15), .ZN(n631) );
  XNOR2_X1 U444 ( .A(G902), .B(KEYINPUT93), .ZN(n463) );
  INV_X1 U445 ( .A(KEYINPUT2), .ZN(n408) );
  NAND2_X1 U446 ( .A1(n359), .A2(n403), .ZN(n404) );
  XNOR2_X1 U447 ( .A(n390), .B(n746), .ZN(n657) );
  XNOR2_X1 U448 ( .A(n516), .B(n352), .ZN(n390) );
  XOR2_X1 U449 ( .A(G101), .B(G140), .Z(n481) );
  INV_X1 U450 ( .A(n580), .ZN(n434) );
  NOR2_X1 U451 ( .A1(n553), .A2(n599), .ZN(n549) );
  INV_X1 U452 ( .A(n386), .ZN(n571) );
  XNOR2_X1 U453 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U454 ( .A(n381), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U455 ( .A1(n383), .A2(n382), .ZN(n381) );
  OR2_X1 U456 ( .A1(n724), .A2(n358), .ZN(n382) );
  XNOR2_X1 U457 ( .A(n688), .B(KEYINPUT84), .ZN(n383) );
  AND2_X1 U458 ( .A1(n688), .A2(n631), .ZN(n346) );
  XOR2_X1 U459 ( .A(n493), .B(n482), .Z(n347) );
  AND2_X1 U460 ( .A1(n554), .A2(n396), .ZN(n348) );
  AND2_X1 U461 ( .A1(n430), .A2(n360), .ZN(n349) );
  AND2_X1 U462 ( .A1(n552), .A2(KEYINPUT88), .ZN(n350) );
  NOR2_X1 U463 ( .A1(n607), .A2(n348), .ZN(n351) );
  XOR2_X1 U464 ( .A(n510), .B(n509), .Z(n352) );
  XOR2_X1 U465 ( .A(G104), .B(G110), .Z(n353) );
  OR2_X1 U466 ( .A1(n712), .A2(KEYINPUT30), .ZN(n354) );
  AND2_X1 U467 ( .A1(n758), .A2(n669), .ZN(n355) );
  AND2_X1 U468 ( .A1(n486), .A2(n590), .ZN(n356) );
  NOR2_X1 U469 ( .A1(n575), .A2(n577), .ZN(n357) );
  NAND2_X1 U470 ( .A1(n750), .A2(n728), .ZN(n358) );
  NAND2_X1 U471 ( .A1(n384), .A2(n355), .ZN(n359) );
  AND2_X1 U472 ( .A1(n429), .A2(KEYINPUT22), .ZN(n360) );
  INV_X1 U473 ( .A(KEYINPUT88), .ZN(n396) );
  XNOR2_X1 U474 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n361) );
  XOR2_X1 U475 ( .A(KEYINPUT87), .B(KEYINPUT35), .Z(n362) );
  XOR2_X1 U476 ( .A(n615), .B(KEYINPUT46), .Z(n363) );
  AND2_X1 U477 ( .A1(n631), .A2(G475), .ZN(n364) );
  AND2_X1 U478 ( .A1(n631), .A2(G472), .ZN(n365) );
  AND2_X1 U479 ( .A1(n631), .A2(G210), .ZN(n366) );
  NAND2_X2 U480 ( .A1(n370), .A2(n367), .ZN(n372) );
  AND2_X2 U481 ( .A1(n371), .A2(n356), .ZN(n370) );
  OR2_X2 U482 ( .A1(n588), .A2(n354), .ZN(n371) );
  XNOR2_X2 U483 ( .A(n372), .B(KEYINPUT79), .ZN(n582) );
  NAND2_X1 U484 ( .A1(n735), .A2(n374), .ZN(n373) );
  INV_X1 U485 ( .A(n628), .ZN(n374) );
  NOR2_X2 U486 ( .A1(n405), .A2(n404), .ZN(n375) );
  NAND2_X1 U487 ( .A1(n380), .A2(n357), .ZN(n379) );
  NAND2_X1 U488 ( .A1(n688), .A2(n365), .ZN(n646) );
  NAND2_X1 U489 ( .A1(n688), .A2(n366), .ZN(n654) );
  NAND2_X1 U490 ( .A1(n688), .A2(n364), .ZN(n659) );
  XNOR2_X1 U491 ( .A(n500), .B(n501), .ZN(n652) );
  XNOR2_X1 U492 ( .A(n560), .B(n385), .ZN(n384) );
  INV_X1 U493 ( .A(n428), .ZN(n427) );
  NOR2_X1 U494 ( .A1(n397), .A2(KEYINPUT88), .ZN(n393) );
  NAND2_X1 U495 ( .A1(n599), .A2(n598), .ZN(n600) );
  BUF_X2 U496 ( .A(n561), .Z(n695) );
  NOR2_X2 U497 ( .A1(n682), .A2(n664), .ZN(n568) );
  XNOR2_X2 U498 ( .A(n563), .B(KEYINPUT31), .ZN(n682) );
  NAND2_X2 U499 ( .A1(n630), .A2(n629), .ZN(n688) );
  XNOR2_X1 U500 ( .A(n547), .B(n546), .ZN(n551) );
  NAND2_X1 U501 ( .A1(n757), .A2(KEYINPUT44), .ZN(n387) );
  NAND2_X1 U502 ( .A1(n428), .A2(n423), .ZN(n422) );
  NAND2_X1 U503 ( .A1(n391), .A2(n617), .ZN(n619) );
  XNOR2_X1 U504 ( .A(n616), .B(n363), .ZN(n391) );
  XNOR2_X2 U505 ( .A(n561), .B(KEYINPUT109), .ZN(n588) );
  OR2_X2 U506 ( .A1(n644), .A2(G902), .ZN(n399) );
  NAND2_X1 U507 ( .A1(n392), .A2(n735), .ZN(n630) );
  XNOR2_X2 U508 ( .A(n628), .B(KEYINPUT85), .ZN(n749) );
  NAND2_X2 U509 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U510 ( .A(n603), .B(KEYINPUT36), .ZN(n397) );
  NOR2_X1 U511 ( .A1(n394), .A2(n393), .ZN(n608) );
  NAND2_X1 U512 ( .A1(n397), .A2(n350), .ZN(n395) );
  AND2_X1 U513 ( .A1(n397), .A2(n552), .ZN(n685) );
  XNOR2_X2 U514 ( .A(n399), .B(n450), .ZN(n561) );
  XNOR2_X2 U515 ( .A(n437), .B(KEYINPUT77), .ZN(n555) );
  NAND2_X1 U516 ( .A1(n400), .A2(n406), .ZN(n405) );
  NAND2_X1 U517 ( .A1(n402), .A2(n401), .ZN(n400) );
  INV_X1 U518 ( .A(n578), .ZN(n402) );
  INV_X1 U519 ( .A(KEYINPUT89), .ZN(n407) );
  OR2_X1 U520 ( .A1(n544), .A2(n545), .ZN(n416) );
  NAND2_X1 U521 ( .A1(n423), .A2(n418), .ZN(n417) );
  INV_X1 U522 ( .A(n424), .ZN(n418) );
  NAND2_X1 U523 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U524 ( .A1(n349), .A2(n424), .ZN(n421) );
  NAND2_X1 U525 ( .A1(n427), .A2(n424), .ZN(n564) );
  NAND2_X1 U526 ( .A1(n420), .A2(n419), .ZN(n553) );
  NOR2_X1 U527 ( .A1(n543), .A2(n431), .ZN(n425) );
  INV_X1 U528 ( .A(n592), .ZN(n426) );
  NAND2_X1 U529 ( .A1(n592), .A2(n431), .ZN(n430) );
  INV_X1 U530 ( .A(KEYINPUT0), .ZN(n431) );
  XNOR2_X2 U531 ( .A(n432), .B(G143), .ZN(n526) );
  XNOR2_X2 U532 ( .A(G128), .B(KEYINPUT65), .ZN(n432) );
  XNOR2_X2 U533 ( .A(n436), .B(KEYINPUT39), .ZN(n533) );
  INV_X1 U534 ( .A(n552), .ZN(n554) );
  NAND2_X1 U535 ( .A1(n551), .A2(n438), .ZN(n437) );
  INV_X1 U536 ( .A(n689), .ZN(n438) );
  XNOR2_X1 U537 ( .A(n556), .B(KEYINPUT33), .ZN(n710) );
  XNOR2_X2 U538 ( .A(n535), .B(n534), .ZN(n614) );
  XNOR2_X1 U539 ( .A(n483), .B(n347), .ZN(n639) );
  AND2_X1 U540 ( .A1(G224), .A2(n750), .ZN(n439) );
  AND2_X1 U541 ( .A1(n574), .A2(n573), .ZN(n440) );
  INV_X1 U542 ( .A(n662), .ZN(n573) );
  INV_X1 U543 ( .A(KEYINPUT24), .ZN(n456) );
  XNOR2_X1 U544 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U545 ( .A(n459), .B(n458), .ZN(n460) );
  INV_X1 U546 ( .A(KEYINPUT19), .ZN(n537) );
  XNOR2_X1 U547 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X2 U548 ( .A(n498), .B(n444), .ZN(n748) );
  XNOR2_X2 U549 ( .A(n748), .B(G146), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n445), .B(KEYINPUT78), .ZN(n511) );
  NAND2_X1 U551 ( .A1(n511), .A2(G210), .ZN(n447) );
  XNOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT5), .ZN(n446) );
  XNOR2_X1 U553 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U554 ( .A(n497), .B(n448), .ZN(n449) );
  XNOR2_X1 U555 ( .A(n483), .B(n449), .ZN(n644) );
  NAND2_X1 U556 ( .A1(n502), .A2(G214), .ZN(n451) );
  XNOR2_X1 U557 ( .A(n451), .B(KEYINPUT98), .ZN(n602) );
  INV_X1 U558 ( .A(n602), .ZN(n712) );
  XNOR2_X1 U559 ( .A(n487), .B(G140), .ZN(n452) );
  XNOR2_X1 U560 ( .A(n452), .B(KEYINPUT10), .ZN(n746) );
  NAND2_X1 U561 ( .A1(G234), .A2(n750), .ZN(n453) );
  XOR2_X1 U562 ( .A(KEYINPUT8), .B(n453), .Z(n525) );
  NAND2_X1 U563 ( .A1(n525), .A2(G221), .ZN(n461) );
  XOR2_X1 U564 ( .A(KEYINPUT83), .B(KEYINPUT23), .Z(n455) );
  XNOR2_X1 U565 ( .A(G128), .B(G110), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n455), .B(n454), .ZN(n459) );
  XNOR2_X1 U567 ( .A(G119), .B(G137), .ZN(n457) );
  XNOR2_X1 U568 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U569 ( .A(n746), .B(n462), .ZN(n729) );
  NOR2_X1 U570 ( .A1(n729), .A2(G902), .ZN(n468) );
  XOR2_X1 U571 ( .A(KEYINPUT20), .B(KEYINPUT101), .Z(n466) );
  INV_X1 U572 ( .A(n631), .ZN(n464) );
  NAND2_X1 U573 ( .A1(G234), .A2(n464), .ZN(n465) );
  XNOR2_X1 U574 ( .A(n466), .B(n465), .ZN(n469) );
  NAND2_X1 U575 ( .A1(G217), .A2(n469), .ZN(n467) );
  NAND2_X1 U576 ( .A1(G221), .A2(n469), .ZN(n471) );
  XOR2_X1 U577 ( .A(KEYINPUT102), .B(KEYINPUT21), .Z(n470) );
  XNOR2_X1 U578 ( .A(n471), .B(n470), .ZN(n691) );
  XNOR2_X1 U579 ( .A(n472), .B(KEYINPUT14), .ZN(n473) );
  XNOR2_X1 U580 ( .A(KEYINPUT76), .B(n473), .ZN(n475) );
  NAND2_X1 U581 ( .A1(n475), .A2(G952), .ZN(n474) );
  XOR2_X1 U582 ( .A(KEYINPUT99), .B(n474), .Z(n722) );
  NOR2_X1 U583 ( .A1(n722), .A2(G953), .ZN(n541) );
  INV_X1 U584 ( .A(n541), .ZN(n478) );
  AND2_X1 U585 ( .A1(n475), .A2(G953), .ZN(n476) );
  NAND2_X1 U586 ( .A1(G902), .A2(n476), .ZN(n539) );
  OR2_X1 U587 ( .A1(n539), .A2(G900), .ZN(n477) );
  NAND2_X1 U588 ( .A1(n478), .A2(n477), .ZN(n587) );
  INV_X1 U589 ( .A(n587), .ZN(n479) );
  NOR2_X1 U590 ( .A1(n689), .A2(n479), .ZN(n486) );
  XNOR2_X1 U591 ( .A(G107), .B(n353), .ZN(n741) );
  XNOR2_X1 U592 ( .A(KEYINPUT70), .B(n741), .ZN(n493) );
  NAND2_X1 U593 ( .A1(G227), .A2(n750), .ZN(n480) );
  XNOR2_X1 U594 ( .A(n481), .B(n480), .ZN(n482) );
  NAND2_X1 U595 ( .A1(n639), .A2(n530), .ZN(n485) );
  INV_X1 U596 ( .A(G469), .ZN(n484) );
  XNOR2_X2 U597 ( .A(n485), .B(n484), .ZN(n547) );
  INV_X1 U598 ( .A(n547), .ZN(n590) );
  XNOR2_X1 U599 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U600 ( .A(n493), .B(n492), .Z(n501) );
  XNOR2_X1 U601 ( .A(n495), .B(n494), .ZN(n496) );
  INV_X1 U602 ( .A(n498), .ZN(n499) );
  XNOR2_X1 U603 ( .A(n739), .B(n499), .ZN(n500) );
  NOR2_X1 U604 ( .A1(n631), .A2(n652), .ZN(n506) );
  NAND2_X1 U605 ( .A1(G210), .A2(n502), .ZN(n504) );
  XOR2_X1 U606 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n503) );
  XNOR2_X1 U607 ( .A(n506), .B(n505), .ZN(n536) );
  INV_X1 U608 ( .A(n536), .ZN(n623) );
  INV_X1 U609 ( .A(KEYINPUT38), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n623), .B(n507), .ZN(n713) );
  INV_X1 U611 ( .A(n713), .ZN(n508) );
  XOR2_X1 U612 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n510) );
  XNOR2_X1 U613 ( .A(G131), .B(KEYINPUT106), .ZN(n509) );
  NAND2_X1 U614 ( .A1(n511), .A2(G214), .ZN(n515) );
  XNOR2_X1 U615 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U616 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U617 ( .A1(n657), .A2(n530), .ZN(n518) );
  XOR2_X1 U618 ( .A(KEYINPUT13), .B(G475), .Z(n517) );
  XNOR2_X1 U619 ( .A(n518), .B(n517), .ZN(n559) );
  XNOR2_X1 U620 ( .A(n520), .B(n519), .ZN(n524) );
  XOR2_X1 U621 ( .A(KEYINPUT7), .B(KEYINPUT107), .Z(n522) );
  XNOR2_X1 U622 ( .A(KEYINPUT9), .B(KEYINPUT108), .ZN(n521) );
  XNOR2_X1 U623 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U624 ( .A(n524), .B(n523), .Z(n529) );
  NAND2_X1 U625 ( .A1(G217), .A2(n525), .ZN(n527) );
  XNOR2_X1 U626 ( .A(n526), .B(n527), .ZN(n528) );
  XNOR2_X1 U627 ( .A(n529), .B(n528), .ZN(n632) );
  NAND2_X1 U628 ( .A1(n632), .A2(n530), .ZN(n531) );
  XNOR2_X1 U629 ( .A(n531), .B(G478), .ZN(n558) );
  INV_X1 U630 ( .A(n558), .ZN(n532) );
  OR2_X1 U631 ( .A1(n559), .A2(n532), .ZN(n670) );
  INV_X1 U632 ( .A(n670), .ZN(n681) );
  AND2_X1 U633 ( .A1(n533), .A2(n681), .ZN(n625) );
  XOR2_X1 U634 ( .A(G134), .B(n625), .Z(G36) );
  AND2_X1 U635 ( .A1(n559), .A2(n532), .ZN(n678) );
  NAND2_X1 U636 ( .A1(n533), .A2(n678), .ZN(n535) );
  INV_X1 U637 ( .A(KEYINPUT40), .ZN(n534) );
  XOR2_X1 U638 ( .A(n614), .B(G131), .Z(G33) );
  NAND2_X1 U639 ( .A1(n536), .A2(n602), .ZN(n538) );
  XNOR2_X2 U640 ( .A(n538), .B(n537), .ZN(n592) );
  NOR2_X1 U641 ( .A1(G898), .A2(n539), .ZN(n540) );
  NOR2_X1 U642 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U643 ( .A(n542), .B(KEYINPUT100), .ZN(n543) );
  NOR2_X1 U644 ( .A1(n559), .A2(n558), .ZN(n709) );
  AND2_X1 U645 ( .A1(n691), .A2(n709), .ZN(n544) );
  INV_X1 U646 ( .A(KEYINPUT22), .ZN(n545) );
  INV_X1 U647 ( .A(KEYINPUT1), .ZN(n546) );
  NOR2_X1 U648 ( .A1(n692), .A2(n554), .ZN(n548) );
  NAND2_X1 U649 ( .A1(n549), .A2(n548), .ZN(n550) );
  BUF_X1 U650 ( .A(n551), .Z(n552) );
  NAND2_X1 U651 ( .A1(n588), .A2(n585), .ZN(n575) );
  OR2_X1 U652 ( .A1(n576), .A2(n575), .ZN(n669) );
  NAND2_X1 U653 ( .A1(n710), .A2(n564), .ZN(n557) );
  NAND2_X1 U654 ( .A1(n559), .A2(n558), .ZN(n580) );
  NOR2_X1 U655 ( .A1(n757), .A2(KEYINPUT44), .ZN(n560) );
  NAND2_X1 U656 ( .A1(n702), .A2(n564), .ZN(n563) );
  INV_X1 U657 ( .A(n564), .ZN(n567) );
  NOR2_X1 U658 ( .A1(n689), .A2(n695), .ZN(n565) );
  NAND2_X1 U659 ( .A1(n565), .A2(n590), .ZN(n566) );
  NOR2_X1 U660 ( .A1(n567), .A2(n566), .ZN(n664) );
  XNOR2_X1 U661 ( .A(KEYINPUT105), .B(n568), .ZN(n569) );
  NOR2_X1 U662 ( .A1(n678), .A2(n681), .ZN(n604) );
  INV_X1 U663 ( .A(n604), .ZN(n707) );
  NAND2_X1 U664 ( .A1(n569), .A2(n707), .ZN(n574) );
  INV_X1 U665 ( .A(n599), .ZN(n570) );
  NAND2_X1 U666 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U667 ( .A1(n585), .A2(n572), .ZN(n662) );
  INV_X1 U668 ( .A(KEYINPUT44), .ZN(n577) );
  XOR2_X1 U669 ( .A(KEYINPUT86), .B(KEYINPUT45), .Z(n579) );
  NAND2_X1 U670 ( .A1(KEYINPUT47), .A2(n604), .ZN(n583) );
  NOR2_X1 U671 ( .A1(n623), .A2(n580), .ZN(n581) );
  NAND2_X1 U672 ( .A1(n582), .A2(n581), .ZN(n673) );
  NAND2_X1 U673 ( .A1(n583), .A2(n673), .ZN(n584) );
  XNOR2_X1 U674 ( .A(n584), .B(KEYINPUT81), .ZN(n594) );
  AND2_X1 U675 ( .A1(n585), .A2(n691), .ZN(n586) );
  NAND2_X1 U676 ( .A1(n587), .A2(n586), .ZN(n597) );
  OR2_X1 U677 ( .A1(n588), .A2(n597), .ZN(n589) );
  XNOR2_X1 U678 ( .A(n589), .B(KEYINPUT28), .ZN(n591) );
  OR2_X1 U679 ( .A1(n591), .A2(n547), .ZN(n612) );
  OR2_X1 U680 ( .A1(n612), .A2(n592), .ZN(n675) );
  NAND2_X1 U681 ( .A1(KEYINPUT47), .A2(n675), .ZN(n593) );
  NAND2_X1 U682 ( .A1(n594), .A2(n593), .ZN(n596) );
  INV_X1 U683 ( .A(KEYINPUT82), .ZN(n595) );
  XNOR2_X1 U684 ( .A(n596), .B(n595), .ZN(n609) );
  INV_X1 U685 ( .A(n678), .ZN(n676) );
  INV_X1 U686 ( .A(n597), .ZN(n598) );
  NOR2_X1 U687 ( .A1(n676), .A2(n600), .ZN(n601) );
  NAND2_X1 U688 ( .A1(n602), .A2(n601), .ZN(n620) );
  NOR2_X1 U689 ( .A1(KEYINPUT47), .A2(n604), .ZN(n605) );
  XNOR2_X1 U690 ( .A(n605), .B(KEYINPUT75), .ZN(n606) );
  NOR2_X1 U691 ( .A1(n675), .A2(n606), .ZN(n607) );
  AND2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n617) );
  NOR2_X1 U693 ( .A1(n713), .A2(n712), .ZN(n706) );
  NAND2_X1 U694 ( .A1(n706), .A2(n709), .ZN(n611) );
  XNOR2_X1 U695 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n610) );
  XNOR2_X1 U696 ( .A(n611), .B(n610), .ZN(n725) );
  NOR2_X1 U697 ( .A1(n725), .A2(n612), .ZN(n613) );
  XNOR2_X1 U698 ( .A(n613), .B(KEYINPUT42), .ZN(n759) );
  NOR2_X2 U699 ( .A1(n614), .A2(n759), .ZN(n616) );
  INV_X1 U700 ( .A(KEYINPUT64), .ZN(n615) );
  INV_X1 U701 ( .A(KEYINPUT48), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n619), .B(n618), .ZN(n627) );
  NOR2_X1 U703 ( .A1(n552), .A2(n620), .ZN(n622) );
  INV_X1 U704 ( .A(KEYINPUT43), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n622), .B(n621), .ZN(n624) );
  AND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n687) );
  NOR2_X1 U707 ( .A1(n687), .A2(n625), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n346), .A2(G478), .ZN(n634) );
  XOR2_X1 U709 ( .A(n632), .B(KEYINPUT124), .Z(n633) );
  XNOR2_X1 U710 ( .A(n634), .B(n633), .ZN(n638) );
  INV_X1 U711 ( .A(G952), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n635), .A2(G953), .ZN(n637) );
  INV_X1 U713 ( .A(KEYINPUT92), .ZN(n636) );
  NOR2_X1 U714 ( .A1(n638), .A2(n732), .ZN(G63) );
  NAND2_X1 U715 ( .A1(n346), .A2(G469), .ZN(n642) );
  XNOR2_X1 U716 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n639), .B(n640), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n642), .B(n641), .ZN(n643) );
  NOR2_X1 U719 ( .A1(n643), .A2(n732), .ZN(G54) );
  XNOR2_X1 U720 ( .A(n644), .B(KEYINPUT62), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U722 ( .A(KEYINPUT112), .B(KEYINPUT63), .Z(n648) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(G57) );
  XNOR2_X1 U724 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(KEYINPUT55), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U730 ( .A(G101), .B(n662), .Z(G3) );
  NAND2_X1 U731 ( .A1(n664), .A2(n678), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n663), .B(G104), .ZN(G6) );
  XOR2_X1 U733 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n666) );
  NAND2_X1 U734 ( .A1(n664), .A2(n681), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n666), .B(n665), .ZN(n668) );
  XOR2_X1 U736 ( .A(G107), .B(KEYINPUT27), .Z(n667) );
  XNOR2_X1 U737 ( .A(n668), .B(n667), .ZN(G9) );
  XNOR2_X1 U738 ( .A(G110), .B(n669), .ZN(G12) );
  NOR2_X1 U739 ( .A1(n670), .A2(n675), .ZN(n672) );
  XNOR2_X1 U740 ( .A(G128), .B(KEYINPUT29), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n672), .B(n671), .ZN(G30) );
  XNOR2_X1 U742 ( .A(G143), .B(KEYINPUT114), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(G45) );
  NOR2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U745 ( .A(G146), .B(n677), .Z(G48) );
  XOR2_X1 U746 ( .A(G113), .B(KEYINPUT115), .Z(n680) );
  NAND2_X1 U747 ( .A1(n682), .A2(n678), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n680), .B(n679), .ZN(G15) );
  NAND2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U750 ( .A(n683), .B(KEYINPUT116), .ZN(n684) );
  XNOR2_X1 U751 ( .A(G116), .B(n684), .ZN(G18) );
  XNOR2_X1 U752 ( .A(G125), .B(n685), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n686), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U754 ( .A(G140), .B(n687), .Z(G42) );
  NAND2_X1 U755 ( .A1(n554), .A2(n689), .ZN(n690) );
  XOR2_X1 U756 ( .A(KEYINPUT50), .B(n690), .Z(n699) );
  XOR2_X1 U757 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n694) );
  OR2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n694), .B(n693), .ZN(n696) );
  NOR2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U761 ( .A(KEYINPUT118), .B(n697), .Z(n698) );
  NOR2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U763 ( .A(KEYINPUT119), .B(n700), .Z(n701) );
  NOR2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U765 ( .A(KEYINPUT51), .B(n703), .Z(n704) );
  XNOR2_X1 U766 ( .A(n704), .B(KEYINPUT120), .ZN(n705) );
  NOR2_X1 U767 ( .A1(n725), .A2(n705), .ZN(n719) );
  AND2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U769 ( .A1(n709), .A2(n708), .ZN(n716) );
  BUF_X1 U770 ( .A(n710), .Z(n711) );
  NAND2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U772 ( .A1(n711), .A2(n714), .ZN(n715) );
  NOR2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U774 ( .A(KEYINPUT121), .B(n717), .Z(n718) );
  NOR2_X1 U775 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U776 ( .A(n720), .B(KEYINPUT52), .ZN(n721) );
  NOR2_X1 U777 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U778 ( .A(KEYINPUT122), .B(n723), .ZN(n724) );
  INV_X1 U779 ( .A(n711), .ZN(n726) );
  NOR2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U781 ( .A(n727), .B(KEYINPUT123), .ZN(n728) );
  NAND2_X1 U782 ( .A1(n346), .A2(G217), .ZN(n730) );
  XNOR2_X1 U783 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(G66) );
  NAND2_X1 U785 ( .A1(G953), .A2(G224), .ZN(n733) );
  XNOR2_X1 U786 ( .A(KEYINPUT61), .B(n733), .ZN(n734) );
  NAND2_X1 U787 ( .A1(n734), .A2(G898), .ZN(n738) );
  NAND2_X1 U788 ( .A1(n750), .A2(n735), .ZN(n736) );
  XOR2_X1 U789 ( .A(KEYINPUT125), .B(n736), .Z(n737) );
  NAND2_X1 U790 ( .A1(n738), .A2(n737), .ZN(n745) );
  XOR2_X1 U791 ( .A(n739), .B(KEYINPUT126), .Z(n740) );
  XNOR2_X1 U792 ( .A(n741), .B(n740), .ZN(n743) );
  NOR2_X1 U793 ( .A1(G898), .A2(n750), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U795 ( .A(n745), .B(n744), .ZN(G69) );
  XNOR2_X1 U796 ( .A(n746), .B(KEYINPUT127), .ZN(n747) );
  XOR2_X1 U797 ( .A(n748), .B(n747), .Z(n752) );
  XNOR2_X1 U798 ( .A(n749), .B(n752), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n751), .A2(n750), .ZN(n756) );
  XOR2_X1 U800 ( .A(G227), .B(n752), .Z(n753) );
  NAND2_X1 U801 ( .A1(n753), .A2(G900), .ZN(n754) );
  NAND2_X1 U802 ( .A1(G953), .A2(n754), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U804 ( .A(n757), .B(G122), .Z(G24) );
  XNOR2_X1 U805 ( .A(n758), .B(G119), .ZN(G21) );
  XOR2_X1 U806 ( .A(G137), .B(n759), .Z(G39) );
endmodule

