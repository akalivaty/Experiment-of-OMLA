//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT65), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT68), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT67), .B(G2105), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT69), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  AOI211_X1 g051(.A(new_n476), .B(new_n472), .C1(new_n469), .C2(new_n470), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n464), .A2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(new_n467), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(new_n472), .A3(G137), .ZN(new_n483));
  AND4_X1   g058(.A1(new_n475), .A2(new_n478), .A3(new_n481), .A4(new_n483), .ZN(G160));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n472), .C2(G112), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT71), .ZN(new_n486));
  INV_X1    g061(.A(new_n482), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(new_n472), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(G2105), .ZN(new_n489));
  AOI22_X1  g064(.A1(G124), .A2(new_n488), .B1(new_n489), .B2(G136), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(new_n482), .A2(G126), .A3(G2105), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(KEYINPUT67), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n499), .A2(new_n501), .A3(G138), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n502), .A2(new_n503), .A3(new_n462), .A4(new_n468), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n482), .A2(new_n472), .A3(G138), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n504), .A2(new_n505), .B1(KEYINPUT4), .B2(new_n506), .ZN(new_n507));
  AND4_X1   g082(.A1(new_n503), .A2(new_n499), .A3(new_n501), .A4(G138), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n508), .A2(KEYINPUT73), .A3(new_n462), .A4(new_n468), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n498), .B1(new_n507), .B2(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(KEYINPUT75), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT74), .A2(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(G62), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT76), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n520), .A2(new_n521), .B1(G75), .B2(G543), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n522), .B1(new_n521), .B2(new_n520), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n519), .B1(new_n523), .B2(G651), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n517), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(new_n515), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT78), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n518), .A2(KEYINPUT77), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT77), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n533), .A2(new_n535), .A3(G543), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n536), .A2(G51), .B1(new_n515), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n532), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n536), .A2(G52), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n529), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G90), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n541), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(new_n536), .A2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n515), .A2(G56), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n543), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(G81), .B2(new_n545), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND4_X1  g135(.A1(new_n533), .A2(new_n535), .A3(G53), .A4(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n563), .A2(KEYINPUT79), .A3(new_n543), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT79), .B1(new_n563), .B2(new_n543), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(new_n565), .B1(G91), .B2(new_n545), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G299));
  XNOR2_X1  g142(.A(new_n547), .B(KEYINPUT80), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G301));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n536), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n545), .A2(G87), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  AND2_X1   g149(.A1(new_n515), .A2(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(G48), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n528), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n515), .A2(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT81), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n536), .A2(G47), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n545), .A2(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n584), .B(new_n585), .C1(new_n543), .C2(new_n586), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n536), .B2(G54), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT82), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n545), .A2(G92), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT10), .Z(new_n595));
  AND2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n589), .B1(new_n588), .B2(new_n596), .ZN(G284));
  AOI21_X1  g172(.A(new_n589), .B1(new_n588), .B2(new_n596), .ZN(G321));
  NAND2_X1  g173(.A1(G299), .A2(new_n588), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n588), .B2(G168), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(new_n588), .B2(G168), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n596), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n596), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g182(.A1(new_n480), .A2(new_n462), .A3(new_n468), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT83), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n489), .A2(G135), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n472), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n488), .A2(new_n617), .A3(G123), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n488), .B2(G123), .ZN(new_n619));
  OAI221_X1 g194(.A(new_n614), .B1(new_n615), .B2(new_n616), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2096), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n610), .B2(new_n611), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n613), .A2(new_n622), .ZN(G156));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(new_n626), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT85), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT86), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n639), .A2(new_n640), .A3(G14), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT18), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(KEYINPUT17), .ZN(new_n649));
  INV_X1    g224(.A(new_n643), .ZN(new_n650));
  INV_X1    g225(.A(new_n644), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n646), .A3(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(new_n645), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n648), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2096), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n666), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT91), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  OAI221_X1 g247(.A(new_n667), .B1(new_n666), .B2(new_n662), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(G229));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n682), .A2(G24), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G290), .B2(G16), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(G1986), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G25), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n488), .A2(G119), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n489), .A2(G131), .ZN(new_n690));
  OAI221_X1 g265(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n472), .C2(G107), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n688), .B1(new_n693), .B2(new_n687), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT35), .B(G1991), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n684), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n682), .A2(G23), .ZN(new_n699));
  AND3_X1   g274(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n682), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT33), .ZN(new_n702));
  INV_X1    g277(.A(G1976), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G6), .B(G305), .S(G16), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT92), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G22), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G166), .B2(G16), .ZN(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n702), .A2(new_n703), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n704), .A2(new_n708), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  AOI211_X1 g289(.A(new_n686), .B(new_n698), .C1(new_n714), .C2(KEYINPUT34), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(KEYINPUT34), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT36), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n687), .A2(G32), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n489), .A2(G141), .B1(new_n480), .B2(G105), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n488), .A2(G129), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT26), .Z(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT96), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(new_n687), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT27), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1996), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n687), .A2(G35), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT99), .Z(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G162), .B2(new_n687), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT29), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(G2090), .ZN(new_n733));
  NOR2_X1   g308(.A1(G168), .A2(new_n682), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n682), .B2(G21), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT97), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n682), .A2(G4), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n596), .B2(new_n682), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G1348), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n728), .A2(new_n733), .A3(new_n738), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n620), .A2(new_n687), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT98), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT30), .B(G28), .Z(new_n746));
  NOR2_X1   g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  AND2_X1   g322(.A1(KEYINPUT31), .A2(G11), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n745), .B1(G29), .B2(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n687), .A2(G26), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n488), .A2(G128), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n489), .A2(G140), .ZN(new_n754));
  OAI221_X1 g329(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n472), .C2(G116), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n752), .B1(new_n756), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n744), .A2(KEYINPUT98), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n749), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n687), .B1(KEYINPUT24), .B2(G34), .ZN(new_n763));
  OAI22_X1  g338(.A1(G160), .A2(new_n687), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G2084), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(G2084), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n682), .A2(G5), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G171), .B2(new_n682), .ZN(new_n768));
  INV_X1    g343(.A(G1961), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n761), .A2(new_n765), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n740), .A2(G1348), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n735), .A2(new_n736), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n682), .A2(G19), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n555), .B2(new_n682), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G1341), .Z(new_n776));
  NOR2_X1   g351(.A1(G27), .A2(G29), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G164), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G2078), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n773), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n742), .A2(new_n771), .A3(new_n772), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n682), .A2(G20), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT23), .Z(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G299), .B2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G1956), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n732), .B2(G2090), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT100), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n687), .A2(G33), .ZN(new_n790));
  NAND2_X1  g365(.A1(G115), .A2(G2104), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n462), .A2(new_n468), .ZN(new_n792));
  INV_X1    g367(.A(G127), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n472), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT25), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G139), .B2(new_n489), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT95), .Z(new_n802));
  OAI21_X1  g377(.A(new_n790), .B1(new_n802), .B2(new_n687), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(G2072), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n788), .A2(KEYINPUT100), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n782), .A2(new_n789), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n717), .A2(new_n806), .ZN(G311));
  INV_X1    g382(.A(G311), .ZN(G150));
  NAND2_X1  g383(.A1(new_n596), .A2(G559), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT38), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n536), .A2(G55), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n545), .A2(G93), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n811), .B(new_n812), .C1(new_n543), .C2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(new_n554), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n810), .B(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n817), .A2(new_n818), .A3(G860), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n814), .A2(G860), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT37), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n819), .A2(new_n821), .ZN(G145));
  XNOR2_X1  g397(.A(G160), .B(new_n620), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n492), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n499), .A2(new_n501), .A3(new_n503), .A4(G138), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n505), .B1(new_n792), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n827), .A2(new_n509), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n498), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n802), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n756), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n802), .A2(new_n832), .A3(new_n756), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n724), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n724), .B1(new_n835), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n831), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(G164), .A3(new_n837), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n692), .B(KEYINPUT102), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n609), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n489), .A2(G142), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n488), .A2(G130), .ZN(new_n846));
  OAI221_X1 g421(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n472), .C2(G118), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n844), .B(new_n848), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT103), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n840), .A2(new_n842), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n840), .B2(new_n842), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n825), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n840), .A2(new_n842), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n849), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n851), .A3(new_n824), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n596), .B(G299), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n604), .B(new_n815), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n862), .B2(new_n866), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n700), .B(KEYINPUT104), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G305), .ZN(new_n870));
  XNOR2_X1  g445(.A(G290), .B(G166), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT42), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n868), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G868), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n814), .A2(new_n588), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n861), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  AOI211_X1 g453(.A(KEYINPUT105), .B(new_n878), .C1(new_n874), .C2(G868), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n877), .A2(new_n879), .ZN(G295));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n876), .ZN(G331));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n882));
  NAND2_X1  g457(.A1(G286), .A2(new_n547), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(G301), .B2(G286), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n815), .ZN(new_n885));
  INV_X1    g460(.A(new_n862), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n863), .A2(new_n885), .A3(new_n864), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n872), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(G37), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n872), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT43), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n888), .ZN(new_n894));
  INV_X1    g469(.A(new_n872), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n858), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT106), .B1(new_n889), .B2(G37), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n882), .B1(new_n893), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n891), .A3(new_n901), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n904), .A2(KEYINPUT43), .B1(new_n890), .B2(new_n900), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n882), .B2(new_n905), .ZN(G397));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(G164), .B2(G1384), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n481), .A2(G40), .A3(new_n483), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n475), .A2(new_n478), .A3(new_n910), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n908), .A2(KEYINPUT107), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT107), .B1(new_n908), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n756), .B(new_n758), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT108), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n915), .B1(new_n724), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(G1996), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n914), .A2(G1996), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n922), .A2(new_n724), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n692), .B(new_n695), .Z(new_n924));
  NAND2_X1  g499(.A1(new_n915), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(G290), .B(new_n697), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n914), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT61), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT50), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT109), .B1(G164), .B2(G1384), .ZN(new_n932));
  AOI21_X1  g507(.A(G1384), .B1(new_n829), .B2(new_n830), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n931), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n474), .A2(new_n477), .A3(new_n909), .ZN(new_n937));
  INV_X1    g512(.A(new_n933), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n937), .B1(new_n938), .B2(KEYINPUT50), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n786), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n911), .B1(KEYINPUT45), .B2(new_n933), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n942));
  XNOR2_X1  g517(.A(KEYINPUT56), .B(G2072), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n908), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n933), .A2(KEYINPUT45), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n908), .A2(new_n945), .A3(new_n937), .A4(new_n943), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT113), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n940), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(G299), .A2(KEYINPUT57), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT57), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n562), .B2(new_n566), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n930), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n934), .B1(new_n831), .B2(new_n955), .ZN(new_n956));
  AOI211_X1 g531(.A(KEYINPUT109), .B(G1384), .C1(new_n829), .C2(new_n830), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT50), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n911), .B1(new_n931), .B2(new_n933), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n960), .A2(new_n786), .B1(KEYINPUT113), .B2(new_n946), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(KEYINPUT117), .A3(new_n952), .A4(new_n944), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n940), .A2(new_n952), .A3(new_n944), .A4(new_n947), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT117), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n954), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n952), .B1(new_n961), .B2(new_n944), .ZN(new_n967));
  AND4_X1   g542(.A1(new_n952), .A2(new_n940), .A3(new_n944), .A4(new_n947), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n930), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n932), .A2(new_n937), .A3(new_n935), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT58), .B(G1341), .Z(new_n971));
  AND2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n908), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n945), .A2(new_n937), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(new_n974), .A3(G1996), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n555), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT59), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT59), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n555), .C1(new_n972), .C2(new_n975), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n966), .A2(new_n969), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT118), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n966), .A2(new_n969), .A3(KEYINPUT118), .A4(new_n980), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n932), .A2(new_n935), .A3(new_n758), .A4(new_n937), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT114), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n956), .A2(new_n957), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n758), .A4(new_n937), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n937), .B1(new_n931), .B2(new_n933), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n987), .B2(new_n931), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n986), .B(new_n989), .C1(new_n991), .C2(G1348), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT60), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n995), .A2(new_n596), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n596), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n983), .A2(new_n984), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n992), .A2(new_n596), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n1000), .A2(new_n1001), .B1(new_n953), .B2(new_n948), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n992), .A2(KEYINPUT115), .A3(new_n596), .ZN(new_n1003));
  AOI211_X1 g578(.A(KEYINPUT116), .B(new_n968), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n948), .A2(new_n953), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n1003), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1005), .B1(new_n1008), .B2(new_n963), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n999), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n990), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n932), .A2(new_n935), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n769), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n907), .B1(new_n956), .B2(new_n957), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1016), .A2(KEYINPUT53), .A3(new_n779), .A4(new_n941), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n908), .A2(new_n945), .A3(new_n779), .A4(new_n937), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1015), .B(new_n1017), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(KEYINPUT122), .A3(new_n568), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT122), .B1(new_n1023), .B2(new_n568), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n471), .A2(new_n473), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n909), .A2(new_n1020), .A3(G2078), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n908), .A2(new_n945), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1015), .B(new_n1030), .C1(new_n1022), .C2(new_n1021), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1031), .A2(new_n568), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT54), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1035));
  NAND3_X1  g610(.A1(G303), .A2(G8), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1035), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(G166), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G2090), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n958), .A2(new_n1042), .A3(new_n959), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n711), .B1(new_n973), .B2(new_n974), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1034), .B(new_n1041), .C1(new_n1045), .C2(new_n1038), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1038), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT112), .B1(new_n1047), .B2(new_n1040), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1012), .B(new_n1042), .C1(new_n1013), .C2(KEYINPUT50), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1038), .B1(new_n1049), .B2(new_n1044), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1040), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n700), .A2(G1976), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n970), .A2(G8), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT52), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT52), .B1(G288), .B2(new_n703), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n970), .A2(G8), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G305), .A2(G1981), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n578), .A2(new_n582), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT111), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(KEYINPUT111), .A3(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1062), .A2(new_n970), .A3(G8), .A4(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1054), .A2(new_n1056), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1046), .A2(new_n1048), .A3(new_n1051), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1966), .B1(new_n1016), .B2(new_n941), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G2084), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1012), .B(new_n1073), .C1(new_n1013), .C2(KEYINPUT50), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1038), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1070), .B1(new_n1075), .B2(G286), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G286), .A2(G8), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT120), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AOI211_X1 g654(.A(G2084), .B(new_n990), .C1(new_n987), .C2(new_n931), .ZN(new_n1080));
  OAI21_X1  g655(.A(G8), .B1(new_n1080), .B2(new_n1071), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1081), .B2(KEYINPUT119), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1075), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1076), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1031), .A2(G171), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1086), .B(KEYINPUT54), .C1(new_n568), .C2(new_n1023), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1081), .A2(new_n1070), .A3(new_n1077), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1069), .A2(new_n1085), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1033), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1011), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  OAI211_X1 g667(.A(G8), .B(G286), .C1(new_n1080), .C2(new_n1071), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT51), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1078), .B1(new_n1075), .B2(new_n1083), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1081), .A2(KEYINPUT119), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1088), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1092), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1026), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1068), .B1(new_n1100), .B2(new_n1024), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1085), .A2(KEYINPUT62), .A3(new_n1088), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n970), .A2(G8), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1059), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G288), .A2(G1976), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1065), .B2(new_n1106), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1051), .A2(new_n1066), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1075), .A2(G168), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1050), .A2(new_n1040), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n1051), .A3(new_n1067), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1068), .B2(new_n1109), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1108), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1103), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n929), .B1(new_n1091), .B2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n922), .A2(KEYINPUT46), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n922), .A2(KEYINPUT46), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n919), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT47), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n921), .A2(new_n923), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n693), .A2(new_n695), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1127), .A2(new_n1128), .B1(G2067), .B2(new_n756), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n915), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1122), .A2(new_n1123), .A3(KEYINPUT123), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n927), .A2(KEYINPUT124), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n926), .A2(new_n1133), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n914), .A2(G1986), .A3(G290), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT48), .Z(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1126), .A2(new_n1130), .A3(new_n1131), .A4(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT125), .B1(new_n1117), .B2(new_n1138), .ZN(new_n1139));
  AND4_X1   g714(.A1(new_n1126), .A2(new_n1130), .A3(new_n1131), .A4(new_n1137), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1103), .A2(new_n1115), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1011), .B2(new_n1090), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1140), .B(new_n1141), .C1(new_n1143), .C2(new_n929), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1139), .A2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g720(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n1147));
  NAND2_X1  g721(.A1(new_n900), .A2(new_n890), .ZN(new_n1148));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g723(.A(G319), .ZN(new_n1150));
  NOR3_X1   g724(.A1(new_n641), .A2(new_n1150), .A3(G227), .ZN(new_n1151));
  OAI21_X1  g725(.A(new_n1151), .B1(new_n679), .B2(new_n680), .ZN(new_n1152));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g728(.A(KEYINPUT126), .B(new_n1151), .C1(new_n679), .C2(new_n680), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AND3_X1   g730(.A1(new_n1149), .A2(new_n859), .A3(new_n1156), .ZN(G308));
  NAND3_X1  g731(.A1(new_n1149), .A2(new_n859), .A3(new_n1156), .ZN(G225));
endmodule


