

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  AND2_X2 U324 ( .A1(n496), .A2(n483), .ZN(n484) );
  XNOR2_X1 U325 ( .A(n377), .B(n301), .ZN(n302) );
  XNOR2_X1 U326 ( .A(n402), .B(KEYINPUT98), .ZN(n403) );
  XNOR2_X1 U327 ( .A(n308), .B(n307), .ZN(n313) );
  XNOR2_X1 U328 ( .A(KEYINPUT25), .B(n407), .ZN(n292) );
  XOR2_X1 U329 ( .A(G218GAT), .B(G99GAT), .Z(n293) );
  AND2_X1 U330 ( .A1(n408), .A2(n292), .ZN(n294) );
  XOR2_X1 U331 ( .A(n305), .B(n304), .Z(n295) );
  XNOR2_X1 U332 ( .A(KEYINPUT119), .B(KEYINPUT45), .ZN(n465) );
  XNOR2_X1 U333 ( .A(n466), .B(n465), .ZN(n467) );
  INV_X1 U334 ( .A(KEYINPUT69), .ZN(n299) );
  INV_X1 U335 ( .A(n377), .ZN(n378) );
  XNOR2_X1 U336 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U337 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U338 ( .A(n447), .B(n293), .ZN(n448) );
  XNOR2_X1 U339 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U340 ( .A(n306), .B(n295), .ZN(n307) );
  XNOR2_X1 U341 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U342 ( .A(KEYINPUT36), .B(n565), .Z(n585) );
  INV_X1 U343 ( .A(KEYINPUT58), .ZN(n480) );
  XOR2_X1 U344 ( .A(n453), .B(n452), .Z(n565) );
  XOR2_X1 U345 ( .A(KEYINPUT116), .B(n457), .Z(n534) );
  XNOR2_X1 U346 ( .A(n485), .B(n484), .ZN(n515) );
  XNOR2_X1 U347 ( .A(n480), .B(G190GAT), .ZN(n481) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n458) );
  XNOR2_X1 U349 ( .A(n486), .B(G43GAT), .ZN(n487) );
  XNOR2_X1 U350 ( .A(n482), .B(n481), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n488), .B(n487), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT33), .B(KEYINPUT68), .Z(n297) );
  XNOR2_X1 U353 ( .A(KEYINPUT67), .B(KEYINPUT73), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n303) );
  XNOR2_X1 U355 ( .A(G148GAT), .B(G106GAT), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n298), .B(G78GAT), .ZN(n377) );
  NAND2_X1 U357 ( .A1(G230GAT), .A2(G233GAT), .ZN(n300) );
  XOR2_X1 U358 ( .A(n303), .B(n302), .Z(n308) );
  XNOR2_X1 U359 ( .A(G85GAT), .B(G92GAT), .ZN(n452) );
  XOR2_X1 U360 ( .A(G57GAT), .B(KEYINPUT13), .Z(n421) );
  XOR2_X1 U361 ( .A(n452), .B(n421), .Z(n306) );
  XOR2_X1 U362 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n305) );
  XNOR2_X1 U363 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n304) );
  XOR2_X1 U364 ( .A(KEYINPUT70), .B(G176GAT), .Z(n310) );
  XNOR2_X1 U365 ( .A(G64GAT), .B(G204GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n366) );
  XNOR2_X1 U367 ( .A(G120GAT), .B(G99GAT), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n311), .B(G71GAT), .ZN(n386) );
  XNOR2_X1 U369 ( .A(n366), .B(n386), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n580) );
  XNOR2_X1 U371 ( .A(n580), .B(KEYINPUT41), .ZN(n557) );
  INV_X1 U372 ( .A(n557), .ZN(n543) );
  XNOR2_X1 U373 ( .A(G1GAT), .B(G8GAT), .ZN(n417) );
  XOR2_X1 U374 ( .A(G50GAT), .B(G43GAT), .Z(n315) );
  XNOR2_X1 U375 ( .A(G141GAT), .B(G36GAT), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n417), .B(n316), .ZN(n318) );
  NAND2_X1 U378 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U380 ( .A(n319), .B(KEYINPUT66), .Z(n322) );
  XNOR2_X1 U381 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n320), .B(KEYINPUT7), .ZN(n443) );
  XNOR2_X1 U383 ( .A(n443), .B(KEYINPUT29), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n330) );
  XOR2_X1 U385 ( .A(G169GAT), .B(G197GAT), .Z(n324) );
  XNOR2_X1 U386 ( .A(G22GAT), .B(G15GAT), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U388 ( .A(KEYINPUT64), .B(KEYINPUT30), .Z(n326) );
  XNOR2_X1 U389 ( .A(G113GAT), .B(KEYINPUT65), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U391 ( .A(n328), .B(n327), .Z(n329) );
  XOR2_X1 U392 ( .A(n330), .B(n329), .Z(n577) );
  INV_X1 U393 ( .A(n577), .ZN(n568) );
  NAND2_X1 U394 ( .A1(n543), .A2(n568), .ZN(n331) );
  XOR2_X1 U395 ( .A(KEYINPUT112), .B(n331), .Z(n518) );
  XOR2_X1 U396 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n333) );
  XNOR2_X1 U397 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n339) );
  XOR2_X1 U399 ( .A(G141GAT), .B(KEYINPUT3), .Z(n335) );
  XNOR2_X1 U400 ( .A(KEYINPUT91), .B(KEYINPUT2), .ZN(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n374) );
  XOR2_X1 U402 ( .A(n374), .B(KEYINPUT5), .Z(n337) );
  NAND2_X1 U403 ( .A1(G225GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n354) );
  XOR2_X1 U406 ( .A(G120GAT), .B(G127GAT), .Z(n341) );
  XNOR2_X1 U407 ( .A(G155GAT), .B(G148GAT), .ZN(n340) );
  XNOR2_X1 U408 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U409 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n343) );
  XNOR2_X1 U410 ( .A(G57GAT), .B(G1GAT), .ZN(n342) );
  XNOR2_X1 U411 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U412 ( .A(n345), .B(n344), .Z(n352) );
  XOR2_X1 U413 ( .A(G134GAT), .B(G85GAT), .Z(n349) );
  XOR2_X1 U414 ( .A(G113GAT), .B(KEYINPUT80), .Z(n347) );
  XNOR2_X1 U415 ( .A(KEYINPUT0), .B(KEYINPUT79), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n347), .B(n346), .ZN(n397) );
  XNOR2_X1 U417 ( .A(G162GAT), .B(n397), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(n350), .ZN(n351) );
  XNOR2_X1 U420 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U421 ( .A(n354), .B(n353), .Z(n529) );
  XOR2_X1 U422 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n356) );
  XNOR2_X1 U423 ( .A(G211GAT), .B(G197GAT), .ZN(n355) );
  XNOR2_X1 U424 ( .A(n356), .B(n355), .ZN(n358) );
  XOR2_X1 U425 ( .A(G218GAT), .B(KEYINPUT21), .Z(n357) );
  XOR2_X1 U426 ( .A(n358), .B(n357), .Z(n384) );
  XNOR2_X1 U427 ( .A(KEYINPUT18), .B(KEYINPUT83), .ZN(n359) );
  XNOR2_X1 U428 ( .A(n359), .B(G169GAT), .ZN(n360) );
  XOR2_X1 U429 ( .A(n360), .B(KEYINPUT17), .Z(n362) );
  XNOR2_X1 U430 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n362), .B(n361), .ZN(n390) );
  XOR2_X1 U432 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n364) );
  XNOR2_X1 U433 ( .A(G92GAT), .B(G8GAT), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n390), .B(n365), .ZN(n370) );
  XOR2_X1 U436 ( .A(G190GAT), .B(G36GAT), .Z(n447) );
  XOR2_X1 U437 ( .A(n447), .B(n366), .Z(n368) );
  NAND2_X1 U438 ( .A1(G226GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U439 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U441 ( .A(n384), .B(n371), .Z(n531) );
  INV_X1 U442 ( .A(n531), .ZN(n510) );
  XOR2_X1 U443 ( .A(n510), .B(KEYINPUT27), .Z(n411) );
  XOR2_X1 U444 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n373) );
  XNOR2_X1 U445 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n372) );
  XNOR2_X1 U446 ( .A(n373), .B(n372), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n374), .B(KEYINPUT88), .ZN(n376) );
  AND2_X1 U448 ( .A1(G228GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U449 ( .A(n376), .B(n375), .ZN(n381) );
  XOR2_X1 U450 ( .A(G162GAT), .B(G50GAT), .Z(n438) );
  XOR2_X1 U451 ( .A(G155GAT), .B(G22GAT), .Z(n424) );
  XNOR2_X1 U452 ( .A(n438), .B(n424), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U454 ( .A(n385), .B(n384), .Z(n474) );
  XOR2_X1 U455 ( .A(G134GAT), .B(G43GAT), .Z(n437) );
  XOR2_X1 U456 ( .A(n437), .B(n386), .Z(n388) );
  NAND2_X1 U457 ( .A1(G227GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n401) );
  XOR2_X1 U460 ( .A(KEYINPUT86), .B(KEYINPUT82), .Z(n392) );
  XNOR2_X1 U461 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n391) );
  XNOR2_X1 U462 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U463 ( .A(n393), .B(KEYINPUT84), .Z(n395) );
  XOR2_X1 U464 ( .A(G127GAT), .B(G15GAT), .Z(n420) );
  XNOR2_X1 U465 ( .A(G190GAT), .B(n420), .ZN(n394) );
  XNOR2_X1 U466 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U467 ( .A(n396), .B(KEYINPUT81), .Z(n399) );
  XNOR2_X1 U468 ( .A(n397), .B(KEYINPUT85), .ZN(n398) );
  XNOR2_X1 U469 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X2 U470 ( .A(n401), .B(n400), .Z(n538) );
  INV_X1 U471 ( .A(n538), .ZN(n500) );
  NAND2_X1 U472 ( .A1(n474), .A2(n500), .ZN(n404) );
  INV_X1 U473 ( .A(KEYINPUT26), .ZN(n402) );
  XNOR2_X1 U474 ( .A(n404), .B(n403), .ZN(n554) );
  AND2_X1 U475 ( .A1(n411), .A2(n554), .ZN(n405) );
  XNOR2_X1 U476 ( .A(n405), .B(KEYINPUT99), .ZN(n408) );
  NOR2_X1 U477 ( .A1(n500), .A2(n510), .ZN(n406) );
  NOR2_X1 U478 ( .A1(n474), .A2(n406), .ZN(n407) );
  XNOR2_X1 U479 ( .A(n294), .B(KEYINPUT100), .ZN(n409) );
  NOR2_X1 U480 ( .A1(n529), .A2(n409), .ZN(n410) );
  XNOR2_X1 U481 ( .A(n410), .B(KEYINPUT101), .ZN(n416) );
  XOR2_X1 U482 ( .A(KEYINPUT28), .B(n474), .Z(n514) );
  INV_X1 U483 ( .A(n514), .ZN(n540) );
  NAND2_X1 U484 ( .A1(n529), .A2(n411), .ZN(n537) );
  NOR2_X1 U485 ( .A1(n540), .A2(n537), .ZN(n412) );
  XOR2_X1 U486 ( .A(KEYINPUT97), .B(n412), .Z(n414) );
  XOR2_X1 U487 ( .A(n500), .B(KEYINPUT87), .Z(n413) );
  NAND2_X1 U488 ( .A1(n414), .A2(n413), .ZN(n415) );
  NAND2_X1 U489 ( .A1(n416), .A2(n415), .ZN(n491) );
  XNOR2_X1 U490 ( .A(G211GAT), .B(G78GAT), .ZN(n419) );
  INV_X1 U491 ( .A(n417), .ZN(n418) );
  XOR2_X1 U492 ( .A(n419), .B(n418), .Z(n435) );
  XOR2_X1 U493 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U494 ( .A1(G231GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U495 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U496 ( .A(n425), .B(n424), .Z(n433) );
  XOR2_X1 U497 ( .A(KEYINPUT14), .B(G64GAT), .Z(n427) );
  XNOR2_X1 U498 ( .A(G183GAT), .B(G71GAT), .ZN(n426) );
  XNOR2_X1 U499 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U500 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n429) );
  XNOR2_X1 U501 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n428) );
  XNOR2_X1 U502 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U503 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U504 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U505 ( .A(n435), .B(n434), .Z(n583) );
  INV_X1 U506 ( .A(n583), .ZN(n571) );
  NAND2_X1 U507 ( .A1(n491), .A2(n571), .ZN(n436) );
  XNOR2_X1 U508 ( .A(n436), .B(KEYINPUT107), .ZN(n454) );
  XOR2_X1 U509 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U510 ( .A1(G232GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U511 ( .A(n440), .B(n439), .ZN(n451) );
  XOR2_X1 U512 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n446) );
  XOR2_X1 U513 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n442) );
  XNOR2_X1 U514 ( .A(KEYINPUT10), .B(G106GAT), .ZN(n441) );
  XNOR2_X1 U515 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U516 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U517 ( .A(n446), .B(n445), .ZN(n449) );
  XNOR2_X1 U518 ( .A(n451), .B(n450), .ZN(n453) );
  NAND2_X1 U519 ( .A1(n454), .A2(n585), .ZN(n456) );
  XNOR2_X1 U520 ( .A(KEYINPUT108), .B(KEYINPUT37), .ZN(n455) );
  XNOR2_X1 U521 ( .A(n456), .B(n455), .ZN(n483) );
  NAND2_X1 U522 ( .A1(n518), .A2(n483), .ZN(n457) );
  NAND2_X1 U523 ( .A1(n534), .A2(n540), .ZN(n459) );
  XNOR2_X1 U524 ( .A(n459), .B(n458), .ZN(G1339GAT) );
  XOR2_X1 U525 ( .A(KEYINPUT46), .B(KEYINPUT118), .Z(n461) );
  NAND2_X1 U526 ( .A1(n543), .A2(n577), .ZN(n460) );
  XNOR2_X1 U527 ( .A(n461), .B(n460), .ZN(n462) );
  INV_X1 U528 ( .A(n565), .ZN(n550) );
  NOR2_X1 U529 ( .A1(n462), .A2(n550), .ZN(n463) );
  NAND2_X1 U530 ( .A1(n463), .A2(n571), .ZN(n464) );
  XNOR2_X1 U531 ( .A(n464), .B(KEYINPUT47), .ZN(n470) );
  NAND2_X1 U532 ( .A1(n583), .A2(n585), .ZN(n466) );
  NAND2_X1 U533 ( .A1(n467), .A2(n568), .ZN(n468) );
  NOR2_X1 U534 ( .A1(n468), .A2(n580), .ZN(n469) );
  NOR2_X1 U535 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U536 ( .A(KEYINPUT48), .B(n471), .ZN(n536) );
  NOR2_X1 U537 ( .A1(n510), .A2(n536), .ZN(n472) );
  XNOR2_X1 U538 ( .A(KEYINPUT54), .B(n472), .ZN(n473) );
  INV_X1 U539 ( .A(n529), .ZN(n507) );
  NAND2_X1 U540 ( .A1(n473), .A2(n507), .ZN(n575) );
  NOR2_X1 U541 ( .A1(n474), .A2(n575), .ZN(n475) );
  XOR2_X1 U542 ( .A(KEYINPUT55), .B(n475), .Z(n476) );
  NAND2_X1 U543 ( .A1(n476), .A2(n538), .ZN(n570) );
  NOR2_X1 U544 ( .A1(n557), .A2(n570), .ZN(n479) );
  XNOR2_X1 U545 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n477) );
  XNOR2_X1 U546 ( .A(n477), .B(G176GAT), .ZN(n478) );
  XNOR2_X1 U547 ( .A(n479), .B(n478), .ZN(G1349GAT) );
  NOR2_X1 U548 ( .A1(n565), .A2(n570), .ZN(n482) );
  INV_X1 U549 ( .A(KEYINPUT38), .ZN(n485) );
  NOR2_X1 U550 ( .A1(n580), .A2(n568), .ZN(n496) );
  NOR2_X1 U551 ( .A1(n500), .A2(n515), .ZN(n488) );
  XNOR2_X1 U552 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n486) );
  XOR2_X1 U553 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n490) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n490), .B(n489), .ZN(n498) );
  NOR2_X1 U556 ( .A1(n571), .A2(n550), .ZN(n493) );
  XNOR2_X1 U557 ( .A(KEYINPUT78), .B(KEYINPUT16), .ZN(n492) );
  XNOR2_X1 U558 ( .A(n493), .B(n492), .ZN(n494) );
  NAND2_X1 U559 ( .A1(n491), .A2(n494), .ZN(n495) );
  XOR2_X1 U560 ( .A(KEYINPUT102), .B(n495), .Z(n517) );
  NAND2_X1 U561 ( .A1(n496), .A2(n517), .ZN(n504) );
  NOR2_X1 U562 ( .A1(n507), .A2(n504), .ZN(n497) );
  XOR2_X1 U563 ( .A(n498), .B(n497), .Z(G1324GAT) );
  NOR2_X1 U564 ( .A1(n510), .A2(n504), .ZN(n499) );
  XOR2_X1 U565 ( .A(G8GAT), .B(n499), .Z(G1325GAT) );
  NOR2_X1 U566 ( .A1(n500), .A2(n504), .ZN(n502) );
  XNOR2_X1 U567 ( .A(KEYINPUT105), .B(KEYINPUT35), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U569 ( .A(G15GAT), .B(n503), .Z(G1326GAT) );
  NOR2_X1 U570 ( .A1(n514), .A2(n504), .ZN(n505) );
  XOR2_X1 U571 ( .A(KEYINPUT106), .B(n505), .Z(n506) );
  XNOR2_X1 U572 ( .A(G22GAT), .B(n506), .ZN(G1327GAT) );
  NOR2_X1 U573 ( .A1(n507), .A2(n515), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(KEYINPUT39), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G29GAT), .B(n509), .ZN(G1328GAT) );
  NOR2_X1 U576 ( .A1(n515), .A2(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G36GAT), .B(n513), .ZN(G1329GAT) );
  NOR2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U581 ( .A(G50GAT), .B(n516), .Z(G1331GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(KEYINPUT113), .B(n519), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n529), .A2(n526), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(KEYINPUT42), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(n521), .ZN(G1332GAT) );
  NAND2_X1 U587 ( .A1(n526), .A2(n531), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(KEYINPUT114), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G64GAT), .B(n523), .ZN(G1333GAT) );
  XOR2_X1 U590 ( .A(G71GAT), .B(KEYINPUT115), .Z(n525) );
  NAND2_X1 U591 ( .A1(n526), .A2(n538), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT43), .Z(n528) );
  NAND2_X1 U594 ( .A1(n526), .A2(n540), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  NAND2_X1 U596 ( .A1(n529), .A2(n534), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G85GAT), .B(n530), .ZN(G1336GAT) );
  XOR2_X1 U598 ( .A(G92GAT), .B(KEYINPUT117), .Z(n533) );
  NAND2_X1 U599 ( .A1(n531), .A2(n534), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(G1337GAT) );
  NAND2_X1 U601 ( .A1(n534), .A2(n538), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(G99GAT), .ZN(G1338GAT) );
  NOR2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n555) );
  NAND2_X1 U604 ( .A1(n555), .A2(n538), .ZN(n539) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n577), .A2(n551), .ZN(n541) );
  XNOR2_X1 U607 ( .A(KEYINPUT120), .B(n541), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT49), .B(KEYINPUT121), .Z(n545) );
  NAND2_X1 U610 ( .A1(n551), .A2(n543), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G120GAT), .B(n546), .Z(G1341GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT50), .B(KEYINPUT122), .Z(n548) );
  NAND2_X1 U614 ( .A1(n551), .A2(n583), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U616 ( .A(G127GAT), .B(n549), .Z(G1342GAT) );
  XOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NAND2_X1 U620 ( .A1(n554), .A2(n555), .ZN(n564) );
  NOR2_X1 U621 ( .A1(n568), .A2(n564), .ZN(n556) );
  XOR2_X1 U622 ( .A(G141GAT), .B(n556), .Z(G1344GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n564), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n571), .A2(n564), .ZN(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n563), .ZN(G1346GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(KEYINPUT125), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1347GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n570), .ZN(n569) );
  XOR2_X1 U635 ( .A(G169GAT), .B(n569), .Z(G1348GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G183GAT), .B(n572), .Z(G1350GAT) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT126), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(n574), .Z(n579) );
  INV_X1 U641 ( .A(n554), .ZN(n576) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n586) );
  NAND2_X1 U643 ( .A1(n586), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U646 ( .A1(n586), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n586), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n588) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

