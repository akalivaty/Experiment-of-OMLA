//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n201), .A2(new_n202), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n203), .A2(new_n204), .A3(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n210), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT65), .Z(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n216), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G97), .B(G107), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G41), .ZN(new_n244));
  INV_X1    g0044(.A(G45), .ZN(new_n245));
  AOI21_X1  g0045(.A(G1), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n246), .A2(new_n248), .A3(G274), .ZN(new_n249));
  INV_X1    g0049(.A(G226), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n249), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G222), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(G223), .A3(G1698), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G77), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n257), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n248), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G169), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT8), .B(G58), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n212), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G150), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n212), .A2(new_n272), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n269), .A2(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(G20), .B1(new_n203), .B2(new_n204), .ZN(new_n277));
  OAI221_X1 g0077(.A(KEYINPUT68), .B1(new_n271), .B2(new_n273), .C1(new_n269), .C2(new_n270), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n282), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(new_n211), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n281), .A2(new_n283), .A3(new_n211), .A4(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n212), .A2(G1), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n287), .A2(new_n290), .B1(G50), .B2(new_n286), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n268), .B(new_n293), .C1(G179), .C2(new_n266), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT69), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n255), .A2(G232), .A3(new_n256), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n255), .A2(G238), .A3(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G107), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n255), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n264), .ZN(new_n300));
  INV_X1    g0100(.A(new_n253), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  AND2_X1   g0102(.A1(G1), .A2(G13), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n247), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n301), .A2(G244), .B1(new_n304), .B2(new_n246), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n267), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n281), .A2(new_n211), .A3(new_n283), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n269), .B(KEYINPUT70), .Z(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n312), .A2(new_n313), .B1(G20), .B2(G77), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT71), .ZN(new_n315));
  INV_X1    g0115(.A(G87), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n316), .A2(KEYINPUT15), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(KEYINPUT15), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT71), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n272), .A2(G20), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n311), .B1(new_n314), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n288), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n329), .A2(new_n287), .B1(G77), .B2(new_n286), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n309), .B(new_n310), .C1(new_n326), .C2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n326), .A2(new_n330), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n306), .A2(G200), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n307), .A2(G190), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n295), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  INV_X1    g0139(.A(G68), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n255), .B2(G20), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G58), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n340), .ZN(new_n346));
  NOR2_X1   g0146(.A1(G58), .A2(G68), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n313), .A2(G159), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n339), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT7), .B1(new_n261), .B2(new_n212), .ZN(new_n352));
  NOR4_X1   g0152(.A1(new_n259), .A2(new_n260), .A3(new_n341), .A4(G20), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n350), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(KEYINPUT16), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(new_n356), .A3(new_n284), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n269), .A2(new_n288), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n287), .ZN(new_n361));
  INV_X1    g0161(.A(new_n286), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n360), .A2(new_n361), .B1(new_n362), .B2(new_n269), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT18), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n248), .A2(G232), .A3(new_n252), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n249), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(G226), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n368));
  OAI211_X1 g0168(.A(G223), .B(new_n256), .C1(new_n259), .C2(new_n260), .ZN(new_n369));
  AND3_X1   g0169(.A1(KEYINPUT75), .A2(G33), .A3(G87), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT75), .B1(G33), .B2(G87), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n367), .B1(new_n264), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n374), .A2(new_n308), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(G169), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n364), .A2(new_n365), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n365), .B1(new_n364), .B2(new_n377), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n264), .ZN(new_n381));
  INV_X1    g0181(.A(G190), .ZN(new_n382));
  INV_X1    g0182(.A(new_n367), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(G200), .B2(new_n374), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n357), .A2(new_n385), .A3(new_n363), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n357), .A2(new_n385), .A3(KEYINPUT17), .A4(new_n363), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n212), .A2(G33), .A3(G77), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n340), .A2(G20), .ZN(new_n392));
  INV_X1    g0192(.A(G50), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n391), .B(new_n392), .C1(new_n273), .C2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n284), .A2(new_n394), .A3(KEYINPUT11), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n289), .A2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n287), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT11), .B1(new_n284), .B2(new_n394), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n286), .A2(G68), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT12), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n250), .A2(new_n256), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n229), .A2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n259), .C2(new_n260), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n264), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n248), .A2(G238), .A3(new_n252), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n249), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT13), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n248), .B1(new_n404), .B2(new_n405), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n249), .A2(new_n408), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT13), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(G190), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n401), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G200), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n411), .B2(new_n414), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n410), .B1(new_n407), .B2(new_n409), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT13), .ZN(new_n421));
  OAI21_X1  g0221(.A(G169), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT14), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n411), .A2(G179), .A3(new_n414), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n425), .B(G169), .C1(new_n420), .C2(new_n421), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n401), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n419), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n338), .A2(new_n380), .A3(new_n390), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n265), .A2(G190), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n417), .B2(new_n265), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n291), .B1(new_n279), .B2(new_n284), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT9), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n432), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT10), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT73), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n265), .A2(new_n417), .ZN(new_n440));
  AOI211_X1 g0240(.A(new_n382), .B(new_n254), .C1(new_n264), .C2(new_n263), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n434), .A2(new_n435), .ZN(new_n443));
  AOI211_X1 g0243(.A(KEYINPUT9), .B(new_n291), .C1(new_n279), .C2(new_n284), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT73), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT10), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n437), .A2(KEYINPUT72), .A3(new_n438), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n442), .B(new_n438), .C1(new_n443), .C2(new_n444), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT72), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n439), .A2(new_n447), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n430), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n272), .A2(G1), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n311), .A2(G116), .A3(new_n286), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n362), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(G20), .B1(G33), .B2(G283), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n272), .A2(G97), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n459), .A2(new_n460), .B1(G20), .B2(new_n457), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n284), .A2(KEYINPUT20), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT20), .B1(new_n284), .B2(new_n461), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n456), .B(new_n458), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n256), .A2(G264), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G257), .A2(G1698), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n465), .A2(new_n466), .B1(new_n259), .B2(new_n260), .ZN(new_n467));
  INV_X1    g0267(.A(new_n260), .ZN(new_n468));
  INV_X1    g0268(.A(G303), .ZN(new_n469));
  NAND2_X1  g0269(.A1(KEYINPUT3), .A2(G33), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n471), .A3(new_n264), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n245), .A2(G1), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n304), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(G270), .A3(new_n248), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n472), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT82), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n472), .A2(new_n479), .A3(KEYINPUT82), .A4(new_n475), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n464), .A2(new_n482), .A3(G169), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n480), .A2(new_n308), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n464), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n484), .B2(new_n485), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n482), .A2(new_n483), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n464), .B1(new_n492), .B2(G190), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n417), .B2(new_n492), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n298), .A2(KEYINPUT23), .A3(G20), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT23), .B1(new_n298), .B2(G20), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G116), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n496), .A2(new_n497), .B1(G20), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n212), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n255), .A2(new_n502), .A3(new_n212), .A4(G87), .ZN(new_n503));
  AOI211_X1 g0303(.A(KEYINPUT24), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(new_n503), .ZN(new_n506));
  INV_X1    g0306(.A(new_n499), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n284), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n362), .A2(new_n298), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT25), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n287), .A2(new_n454), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(G107), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n478), .A2(G264), .A3(new_n248), .ZN(new_n515));
  NOR2_X1   g0315(.A1(G250), .A2(G1698), .ZN(new_n516));
  INV_X1    g0316(.A(G257), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(G1698), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(new_n255), .B1(G33), .B2(G294), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n475), .B(new_n515), .C1(new_n519), .C2(new_n248), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G169), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(G1698), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(G250), .B2(G1698), .ZN(new_n523));
  INV_X1    g0323(.A(G294), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n523), .A2(new_n261), .B1(new_n272), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n264), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n526), .A2(G179), .A3(new_n475), .A4(new_n515), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT83), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n521), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n514), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT84), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT84), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n514), .A2(new_n529), .A3(new_n534), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n520), .A2(G200), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n382), .B2(new_n520), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n514), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n533), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n313), .A2(KEYINPUT76), .A3(G77), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT76), .B1(new_n313), .B2(G77), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT6), .ZN(new_n544));
  INV_X1    g0344(.A(G97), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n544), .A2(new_n545), .A3(G107), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n543), .B1(new_n548), .B2(new_n212), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n298), .B1(new_n342), .B2(new_n343), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n284), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n512), .A2(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n362), .A2(new_n545), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT78), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G244), .B(new_n256), .C1(new_n259), .C2(new_n260), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT4), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(G283), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n272), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G250), .A2(G1698), .ZN(new_n562));
  NAND2_X1  g0362(.A1(KEYINPUT4), .A2(G244), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(G1698), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n255), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n248), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n478), .A2(G257), .A3(new_n248), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n475), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n267), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n568), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n566), .A2(KEYINPUT77), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT77), .ZN(new_n572));
  AOI211_X1 g0372(.A(new_n572), .B(new_n248), .C1(new_n559), .C2(new_n565), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n308), .B(new_n570), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n551), .A2(KEYINPUT78), .A3(new_n552), .A4(new_n553), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n556), .A2(new_n569), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n566), .A2(new_n568), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n559), .A2(new_n565), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n572), .B1(new_n580), .B2(new_n248), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n566), .A2(KEYINPUT77), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n568), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n577), .B(new_n579), .C1(new_n417), .C2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G250), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n251), .B2(G45), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n304), .A2(new_n473), .B1(new_n248), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n498), .ZN(new_n588));
  NOR2_X1   g0388(.A1(G238), .A2(G1698), .ZN(new_n589));
  INV_X1    g0389(.A(G244), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(G1698), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n588), .B1(new_n591), .B2(new_n255), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n587), .B1(new_n592), .B2(new_n248), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(G179), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n267), .B2(new_n593), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT81), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n286), .B1(new_n319), .B2(new_n321), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n212), .B(G68), .C1(new_n259), .C2(new_n260), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT80), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT80), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n255), .A2(new_n600), .A3(new_n212), .A4(G68), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT19), .B1(new_n324), .B2(G97), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n316), .A2(KEYINPUT79), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT79), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G87), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(new_n606), .A3(new_n545), .A4(new_n298), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n405), .B2(new_n212), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n603), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n597), .B1(new_n611), .B2(new_n284), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n322), .A2(new_n287), .A3(new_n454), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n596), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n311), .B1(new_n602), .B2(new_n610), .ZN(new_n616));
  NOR4_X1   g0416(.A1(new_n616), .A2(new_n613), .A3(KEYINPUT81), .A4(new_n597), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n595), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n512), .A2(G87), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n593), .A2(G200), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n382), .B2(new_n593), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n576), .A2(new_n584), .A3(new_n618), .A4(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n453), .A2(new_n495), .A3(new_n540), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT85), .ZN(G372));
  INV_X1    g0427(.A(new_n295), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n364), .A2(new_n377), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT18), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n364), .A2(new_n377), .A3(new_n365), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n426), .A2(new_n424), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n411), .A2(new_n414), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n425), .B1(new_n634), .B2(G169), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n428), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n331), .B2(new_n419), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n632), .B1(new_n637), .B2(new_n390), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n628), .B1(new_n452), .B2(new_n638), .ZN(new_n639));
  XOR2_X1   g0439(.A(new_n639), .B(KEYINPUT86), .Z(new_n640));
  AOI22_X1  g0440(.A1(new_n509), .A2(new_n513), .B1(new_n521), .B2(new_n527), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n487), .A2(new_n490), .A3(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n624), .A2(new_n642), .A3(new_n538), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n618), .A2(new_n623), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT26), .B1(new_n644), .B2(new_n576), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n574), .A2(new_n569), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n577), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n647), .A2(new_n618), .A3(new_n648), .A4(new_n623), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n645), .A2(new_n618), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n453), .B1(new_n643), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n640), .A2(new_n651), .ZN(G369));
  NAND3_X1  g0452(.A1(new_n251), .A2(new_n212), .A3(G13), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n464), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n495), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n491), .B2(new_n659), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n514), .ZN(new_n664));
  INV_X1    g0464(.A(new_n658), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n540), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n532), .B2(new_n665), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n484), .A2(new_n485), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n486), .A3(new_n489), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n665), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n540), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n641), .A2(new_n665), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT87), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n673), .A2(KEYINPUT87), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n668), .A2(new_n679), .ZN(G399));
  NOR2_X1   g0480(.A1(new_n607), .A2(G116), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n208), .A2(new_n244), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n214), .B2(new_n682), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n620), .A2(new_n622), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n611), .A2(new_n284), .ZN(new_n687));
  INV_X1    g0487(.A(new_n597), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n614), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT81), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n612), .A2(new_n596), .A3(new_n614), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n686), .B1(new_n692), .B2(new_n595), .ZN(new_n693));
  INV_X1    g0493(.A(new_n576), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n648), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n647), .A2(new_n618), .A3(new_n623), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT26), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n695), .A2(new_n697), .A3(new_n618), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n533), .A2(new_n535), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n625), .B(new_n539), .C1(new_n670), .C2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .A3(new_n665), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n650), .A2(new_n643), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n658), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n704), .B2(KEYINPUT29), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT90), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n515), .B1(new_n519), .B2(new_n248), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT88), .B1(new_n707), .B2(new_n593), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n474), .A2(new_n473), .B1(new_n303), .B2(new_n247), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n525), .A2(new_n264), .B1(new_n709), .B2(G264), .ZN(new_n710));
  OR2_X1    g0510(.A1(G238), .A2(G1698), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n590), .A2(G1698), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n711), .B(new_n712), .C1(new_n259), .C2(new_n260), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n248), .B1(new_n713), .B2(new_n498), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n248), .A2(G274), .A3(new_n473), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n586), .A2(new_n248), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT88), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n710), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n708), .A2(new_n720), .A3(new_n488), .A4(new_n578), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n566), .A2(new_n568), .A3(new_n722), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n708), .A2(new_n720), .A3(new_n724), .A4(new_n488), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n570), .B1(new_n571), .B2(new_n573), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n520), .A2(new_n308), .A3(new_n593), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n482), .A4(new_n483), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n723), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n665), .B1(new_n729), .B2(KEYINPUT89), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT89), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n723), .A2(new_n728), .A3(new_n731), .A4(new_n725), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT31), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n706), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n721), .A2(new_n722), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n718), .A2(G179), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(new_n482), .A3(new_n483), .A4(new_n520), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n725), .B1(new_n738), .B2(new_n583), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT89), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n658), .A3(new_n732), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n734), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(KEYINPUT90), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n540), .A2(new_n625), .A3(new_n495), .A4(new_n665), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n735), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n705), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n685), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(G13), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n251), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n682), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n661), .A2(G330), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n663), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT91), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n661), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n211), .B1(G20), .B2(new_n267), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n212), .A2(G179), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n604), .B2(new_n606), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n382), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n212), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n769), .B1(G97), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n212), .A2(new_n308), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n382), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n767), .A2(new_n382), .A3(G200), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n773), .B1(new_n393), .B2(new_n777), .C1(new_n298), .C2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT92), .B(G159), .Z(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n767), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT32), .ZN(new_n783));
  OAI21_X1  g0583(.A(KEYINPUT32), .B1(new_n780), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n775), .A2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n784), .B1(new_n786), .B2(new_n340), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n774), .A2(new_n781), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n774), .A2(G190), .A3(new_n417), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n255), .B1(new_n788), .B2(new_n327), .C1(new_n345), .C2(new_n789), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n779), .A2(new_n783), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G317), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n785), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G326), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n469), .B2(new_n768), .C1(new_n796), .C2(new_n777), .ZN(new_n797));
  INV_X1    g0597(.A(new_n789), .ZN(new_n798));
  INV_X1    g0598(.A(new_n782), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n798), .A2(G322), .B1(new_n799), .B2(G329), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n800), .B(new_n261), .C1(new_n801), .C2(new_n788), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n771), .A2(new_n524), .B1(new_n778), .B2(new_n560), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n797), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n766), .B1(new_n791), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n763), .A2(new_n766), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n255), .A2(new_n208), .ZN(new_n808));
  INV_X1    g0608(.A(G355), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n808), .A2(new_n809), .B1(G116), .B2(new_n208), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n239), .A2(new_n245), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n261), .A2(new_n208), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n245), .B2(new_n215), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n810), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n805), .B(new_n757), .C1(new_n807), .C2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n760), .B1(new_n765), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  NOR2_X1   g0618(.A1(new_n331), .A2(new_n658), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n336), .B1(new_n333), .B2(new_n665), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n820), .B2(new_n331), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n704), .B(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n757), .B1(new_n822), .B2(new_n748), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n748), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n778), .A2(new_n340), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n261), .B(new_n825), .C1(G132), .C2(new_n799), .ZN(new_n826));
  INV_X1    g0626(.A(new_n768), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n772), .A2(G58), .B1(new_n827), .B2(G50), .ZN(new_n828));
  INV_X1    g0628(.A(new_n780), .ZN(new_n829));
  INV_X1    g0629(.A(new_n788), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G143), .A2(new_n798), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n832), .B2(new_n777), .C1(new_n271), .C2(new_n786), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n826), .B(new_n828), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n560), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n772), .A2(G97), .B1(new_n827), .B2(G107), .ZN(new_n841));
  INV_X1    g0641(.A(new_n778), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n776), .A2(G303), .B1(new_n842), .B2(G87), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n255), .B1(new_n798), .B2(G294), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G116), .A2(new_n830), .B1(new_n799), .B2(G311), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n841), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n835), .A2(new_n836), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n766), .ZN(new_n848));
  INV_X1    g0648(.A(new_n757), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n766), .A2(new_n761), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n327), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(new_n821), .C2(new_n762), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n824), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  NAND2_X1  g0654(.A1(new_n213), .A2(G116), .ZN(new_n855));
  INV_X1    g0655(.A(new_n548), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(KEYINPUT35), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(KEYINPUT35), .B2(new_n856), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT36), .ZN(new_n859));
  OAI21_X1  g0659(.A(G77), .B1(new_n345), .B2(new_n340), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n860), .A2(new_n214), .B1(G50), .B2(new_n340), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(G1), .A3(new_n752), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT96), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n656), .B1(new_n357), .B2(new_n363), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n388), .A2(new_n389), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n865), .B1(new_n632), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n357), .A2(new_n385), .A3(new_n363), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(new_n865), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT100), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n869), .B(new_n629), .C1(new_n870), .C2(KEYINPUT37), .ZN(new_n871));
  INV_X1    g0671(.A(new_n656), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n364), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n629), .A2(new_n873), .A3(new_n386), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n870), .A3(new_n386), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n871), .A4(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT101), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n871), .A2(new_n877), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n881), .A2(KEYINPUT101), .A3(KEYINPUT38), .A4(new_n867), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n871), .A2(new_n877), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n873), .B1(new_n380), .B2(new_n390), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n866), .A2(KEYINPUT102), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n388), .A2(new_n891), .A3(new_n389), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n380), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n884), .B1(new_n865), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n889), .B(new_n878), .C1(new_n894), .C2(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n427), .A2(new_n428), .A3(new_n665), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n665), .B(new_n821), .C1(new_n650), .C2(new_n643), .ZN(new_n900));
  INV_X1    g0700(.A(new_n819), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n427), .A2(new_n419), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n428), .A2(new_n658), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT97), .B1(new_n429), .B2(new_n904), .ZN(new_n906));
  INV_X1    g0706(.A(new_n419), .ZN(new_n907));
  AND4_X1   g0707(.A1(KEYINPUT97), .A2(new_n636), .A3(new_n907), .A4(new_n904), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n905), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT98), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n636), .A2(new_n907), .A3(new_n904), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT97), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n429), .A2(KEYINPUT97), .A3(new_n904), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT98), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(new_n905), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n902), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT99), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n901), .A2(new_n900), .B1(new_n910), .B2(new_n917), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT99), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(new_n923), .A3(new_n887), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n632), .A2(new_n656), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n899), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n702), .B(new_n453), .C1(KEYINPUT29), .C2(new_n704), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n927), .A2(new_n640), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(G330), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n732), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n746), .A2(new_n743), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n903), .A2(new_n904), .ZN(new_n933));
  AOI211_X1 g0733(.A(KEYINPUT98), .B(new_n933), .C1(new_n913), .C2(new_n914), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n916), .B1(new_n915), .B2(new_n905), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n932), .B(new_n821), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n893), .A2(new_n865), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n937), .B2(new_n881), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n884), .A2(new_n885), .A3(new_n883), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT40), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n821), .ZN(new_n942));
  AND4_X1   g0742(.A1(KEYINPUT31), .A2(new_n740), .A3(new_n658), .A4(new_n732), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n733), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n942), .B1(new_n944), .B2(new_n746), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n887), .A2(new_n945), .A3(new_n946), .A4(new_n918), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n453), .A2(new_n932), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n930), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n929), .A2(new_n951), .B1(new_n251), .B2(new_n753), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT103), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n929), .A2(new_n951), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n952), .A2(KEYINPUT103), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n864), .B1(new_n955), .B2(new_n956), .ZN(G367));
  NAND2_X1  g0757(.A1(new_n554), .A2(new_n658), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n576), .A2(new_n584), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n646), .A2(new_n958), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n540), .A2(new_n672), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT42), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT105), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT106), .ZN(new_n965));
  INV_X1    g0765(.A(new_n961), .ZN(new_n966));
  INV_X1    g0766(.A(new_n699), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n576), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n968), .A2(new_n665), .B1(KEYINPUT42), .B2(new_n962), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n964), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n965), .B1(new_n964), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n620), .A2(new_n658), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n693), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(KEYINPUT104), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(KEYINPUT104), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n618), .C2(new_n972), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT43), .Z(new_n977));
  OR3_X1    g0777(.A1(new_n970), .A2(new_n971), .A3(new_n977), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n970), .A2(new_n971), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n663), .A2(new_n667), .A3(new_n961), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n682), .B(KEYINPUT41), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n679), .A2(new_n961), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n677), .A2(new_n678), .A3(new_n966), .ZN(new_n987));
  NOR2_X1   g0787(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND2_X1  g0790(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n668), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n673), .B1(new_n667), .B2(new_n672), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n663), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n986), .A2(new_n668), .A3(new_n992), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n750), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n983), .B1(new_n998), .B2(new_n750), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n982), .B1(new_n999), .B2(new_n755), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n806), .B1(new_n208), .B2(new_n322), .C1(new_n235), .C2(new_n812), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1001), .A2(new_n757), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n766), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n261), .B1(new_n789), .B2(new_n469), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G317), .B2(new_n799), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n776), .A2(G311), .B1(new_n842), .B2(G97), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(new_n839), .C2(new_n524), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n771), .A2(new_n298), .B1(new_n788), .B2(new_n560), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT108), .Z(new_n1009));
  NAND2_X1  g0809(.A1(new_n827), .A2(G116), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT46), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n839), .A2(new_n780), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n771), .A2(new_n340), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G58), .B2(new_n827), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n261), .B1(new_n798), .B2(G150), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G50), .A2(new_n830), .B1(new_n799), .B2(G137), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n776), .A2(G143), .B1(new_n842), .B2(G77), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1007), .A2(new_n1012), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  OAI221_X1 g0821(.A(new_n1002), .B1(new_n1003), .B2(new_n1021), .C1(new_n976), .C2(new_n764), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1000), .A2(new_n1022), .ZN(G387));
  OAI22_X1  g0823(.A1(new_n681), .A2(new_n808), .B1(G107), .B2(new_n208), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n232), .A2(new_n245), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT109), .Z(new_n1026));
  NAND2_X1  g0826(.A1(new_n312), .A2(new_n393), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT50), .Z(new_n1028));
  INV_X1    g0828(.A(new_n681), .ZN(new_n1029));
  AOI211_X1 g0829(.A(G45), .B(new_n1029), .C1(G68), .C2(G77), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n812), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1024), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT110), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n806), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n757), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n789), .A2(new_n393), .B1(new_n782), .B2(new_n271), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n261), .B(new_n1037), .C1(G68), .C2(new_n830), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n768), .A2(new_n327), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G97), .B2(new_n842), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n269), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G159), .A2(new_n776), .B1(new_n785), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n323), .A2(new_n772), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n839), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1046), .A2(G311), .B1(G322), .B2(new_n776), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1047), .A2(KEYINPUT112), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(KEYINPUT112), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n798), .A2(G317), .B1(new_n830), .B2(G303), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n772), .A2(G283), .B1(new_n827), .B2(G294), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT49), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n261), .B1(new_n782), .B2(new_n796), .C1(new_n457), .C2(new_n778), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1045), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1036), .B1(new_n1062), .B2(new_n766), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n667), .A2(new_n764), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1063), .A2(new_n1064), .B1(new_n755), .B2(new_n996), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n750), .A2(new_n996), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n756), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n750), .A2(new_n996), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(G393));
  INV_X1    g0869(.A(new_n997), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1066), .B1(new_n1070), .B2(new_n993), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n998), .A2(new_n1071), .A3(new_n756), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n261), .B1(new_n799), .B2(G143), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n340), .B2(new_n768), .C1(new_n316), .C2(new_n778), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT114), .Z(new_n1075));
  NAND2_X1  g0875(.A1(new_n1046), .A2(G50), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n312), .A2(new_n830), .B1(G77), .B2(new_n772), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G150), .A2(new_n776), .B1(new_n798), .B2(G159), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT51), .Z(new_n1079));
  NAND4_X1  g0879(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1046), .A2(G303), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n777), .A2(new_n792), .B1(new_n801), .B2(new_n789), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT52), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n788), .A2(new_n524), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n255), .B(new_n1084), .C1(G322), .C2(new_n799), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n298), .A2(new_n778), .B1(new_n768), .B2(new_n560), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G116), .B2(new_n772), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1081), .A2(new_n1083), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1003), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n806), .B1(new_n545), .B2(new_n208), .C1(new_n242), .C2(new_n812), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n757), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT113), .Z(new_n1092));
  AOI211_X1 g0892(.A(new_n1089), .B(new_n1092), .C1(new_n966), .C2(new_n763), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1070), .A2(new_n993), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n755), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1072), .A2(new_n1095), .ZN(G390));
  NOR3_X1   g0896(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT39), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(KEYINPUT39), .B2(new_n887), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT115), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n922), .B2(new_n898), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n919), .A2(KEYINPUT115), .A3(new_n897), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n747), .A2(new_n918), .A3(G330), .A4(new_n821), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n878), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n658), .B1(new_n698), .B2(new_n700), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n820), .A2(new_n331), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n819), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n934), .A2(new_n935), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n897), .B(new_n1104), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1102), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n945), .A2(G330), .A3(new_n918), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1102), .B2(new_n1109), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1098), .A2(new_n761), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n839), .A2(new_n298), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n261), .B1(new_n788), .B2(new_n545), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n789), .A2(new_n457), .B1(new_n782), .B2(new_n524), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n825), .B1(G77), .B2(new_n772), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n316), .B2(new_n768), .C1(new_n560), .C2(new_n777), .ZN(new_n1119));
  NOR4_X1   g0919(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G159), .A2(new_n772), .B1(new_n776), .B2(G128), .ZN(new_n1121));
  XOR2_X1   g0921(.A(KEYINPUT54), .B(G143), .Z(new_n1122));
  AOI21_X1  g0922(.A(new_n261), .B1(new_n830), .B2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n798), .A2(G132), .B1(new_n799), .B2(G125), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n842), .A2(G50), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n768), .A2(new_n271), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT53), .Z(new_n1128));
  AOI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(new_n1046), .C2(G137), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1120), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n1003), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n849), .B(new_n1131), .C1(new_n269), .C2(new_n850), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1113), .A2(new_n755), .B1(new_n1114), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n453), .A2(G330), .A3(new_n932), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n927), .A2(new_n640), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n902), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n734), .B1(new_n741), .B2(new_n742), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n746), .B1(new_n1137), .B2(KEYINPUT90), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n733), .A2(new_n706), .A3(new_n734), .ZN(new_n1139));
  OAI211_X1 g0939(.A(G330), .B(new_n821), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1108), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1136), .B1(new_n1141), .B2(new_n1111), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n932), .A2(G330), .A3(new_n821), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1108), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1103), .A2(new_n1107), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1135), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT116), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1135), .B(KEYINPUT116), .C1(new_n1142), .C2(new_n1145), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n756), .B1(new_n1150), .B2(new_n1113), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1102), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1109), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT115), .B1(new_n919), .B2(new_n897), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(new_n896), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n1155), .B2(new_n1101), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1152), .B1(new_n1156), .B2(new_n1111), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1133), .B1(new_n1151), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT117), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(KEYINPUT117), .B(new_n1133), .C1(new_n1151), .C2(new_n1158), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(G378));
  NOR2_X1   g0964(.A1(new_n434), .A2(new_n656), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n294), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n452), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1165), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n447), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n446), .B1(new_n445), .B2(KEYINPUT10), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n449), .B(KEYINPUT72), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n294), .B(new_n1168), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1167), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n945), .A2(new_n946), .A3(new_n918), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1104), .A2(new_n945), .A3(new_n918), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1178), .A2(new_n887), .B1(new_n1179), .B2(KEYINPUT40), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1177), .B1(new_n1180), .B2(new_n930), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1177), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n948), .A2(G330), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n926), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n899), .A2(new_n924), .A3(new_n925), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1182), .B1(new_n948), .B2(G330), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n930), .B(new_n1177), .C1(new_n941), .C2(new_n947), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n755), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n849), .B1(new_n393), .B2(new_n850), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n780), .B2(new_n778), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n827), .A2(new_n1122), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT118), .Z(new_n1195));
  NAND2_X1  g0995(.A1(new_n776), .A2(G125), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n798), .A2(G128), .B1(new_n830), .B2(G137), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G150), .A2(new_n772), .B1(new_n785), .B2(G132), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT119), .Z(new_n1200));
  AOI21_X1  g1000(.A(new_n1193), .B1(new_n1200), .B2(KEYINPUT59), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(KEYINPUT59), .B2(new_n1200), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n777), .A2(new_n457), .B1(new_n778), .B2(new_n345), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G97), .B2(new_n785), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n255), .A2(G41), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n560), .B2(new_n782), .C1(new_n298), .C2(new_n789), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1206), .A2(new_n1014), .A3(new_n1039), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1204), .B(new_n1207), .C1(new_n322), .C2(new_n788), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT58), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1205), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(new_n393), .C1(G33), .C2(G41), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1213));
  AND4_X1   g1013(.A1(new_n1202), .A2(new_n1210), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1191), .B1(new_n1003), .B2(new_n1214), .C1(new_n1182), .C2(new_n762), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT120), .Z(new_n1216));
  AND2_X1   g1016(.A1(new_n1190), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT121), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1184), .B2(new_n1188), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT121), .B1(new_n1220), .B2(new_n1185), .ZN(new_n1221));
  OAI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1135), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1150), .B2(new_n1113), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n756), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1150), .A2(new_n1113), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1135), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1189), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1217), .B1(new_n1225), .B2(new_n1228), .ZN(G375));
  OR3_X1    g1029(.A1(new_n1135), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1148), .A2(new_n1230), .A3(new_n1149), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(new_n983), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT122), .Z(new_n1233));
  OAI21_X1  g1033(.A(new_n755), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n849), .B1(new_n340), .B2(new_n850), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1046), .A2(new_n1122), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n789), .A2(new_n832), .B1(new_n788), .B2(new_n271), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n261), .B(new_n1237), .C1(G128), .C2(new_n799), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n776), .A2(G132), .B1(new_n842), .B2(G58), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n772), .A2(G50), .B1(new_n827), .B2(G159), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1046), .A2(G116), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n777), .A2(new_n524), .B1(new_n778), .B2(new_n327), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G97), .B2(new_n827), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n788), .A2(new_n298), .B1(new_n782), .B2(new_n469), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n255), .B(new_n1245), .C1(G283), .C2(new_n798), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1242), .A2(new_n1043), .A3(new_n1244), .A4(new_n1246), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1241), .A2(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1235), .B1(new_n1003), .B2(new_n1248), .C1(new_n918), .C2(new_n762), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1234), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1233), .A2(new_n1250), .ZN(G381));
  OR2_X1    g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(G387), .A2(G384), .A3(G390), .A4(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n1250), .A3(new_n1233), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(KEYINPUT123), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1159), .ZN(new_n1256));
  INV_X1    g1056(.A(G375), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(KEYINPUT123), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(G407));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n657), .A3(new_n1256), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(G407), .A2(G213), .A3(new_n1260), .ZN(G409));
  AND3_X1   g1061(.A1(new_n1000), .A2(new_n1022), .A3(G390), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G390), .B1(new_n1000), .B2(new_n1022), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT124), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(G393), .B(G396), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(KEYINPUT124), .B(new_n1265), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1189), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1224), .A2(new_n1270), .A3(new_n983), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n755), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1216), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1256), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(G375), .B2(new_n1163), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n657), .A2(G213), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT60), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n682), .B1(new_n1230), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1231), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1278), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1250), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n853), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(G384), .A3(new_n1250), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1276), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(G2897), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1277), .B2(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1275), .A2(new_n1291), .A3(new_n1276), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT57), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1224), .B2(new_n1270), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1296), .B(new_n756), .C1(new_n1224), .C2(new_n1222), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1297), .A2(new_n1161), .A3(new_n1162), .A4(new_n1217), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1285), .B1(new_n1298), .B2(new_n1274), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1269), .A2(new_n1290), .A3(new_n1294), .A4(new_n1300), .ZN(new_n1301));
  AND4_X1   g1101(.A1(KEYINPUT62), .A2(new_n1275), .A3(new_n1291), .A4(new_n1276), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT62), .B1(new_n1299), .B2(new_n1291), .ZN(new_n1303));
  OAI211_X1 g1103(.A(KEYINPUT125), .B(new_n1290), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT126), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1267), .A2(new_n1305), .A3(new_n1268), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1292), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1299), .A2(KEYINPUT62), .A3(new_n1291), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT125), .B1(new_n1313), .B2(new_n1290), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1301), .B1(new_n1309), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT127), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1317), .B(new_n1301), .C1(new_n1309), .C2(new_n1314), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(G405));
  OAI21_X1  g1119(.A(new_n1298), .B1(new_n1257), .B2(new_n1159), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(new_n1291), .ZN(new_n1321));
  XOR2_X1   g1121(.A(new_n1321), .B(new_n1269), .Z(G402));
endmodule


