//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n205), .A2(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(KEYINPUT15), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n210));
  XOR2_X1   g009(.A(new_n209), .B(new_n210), .Z(new_n211));
  INV_X1    g010(.A(KEYINPUT17), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(G1gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT16), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n209), .B(new_n210), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n213), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT84), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n218), .B(G8gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n211), .B2(new_n226), .ZN(new_n227));
  NOR3_X1   g026(.A1(new_n221), .A2(new_n220), .A3(KEYINPUT84), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n223), .B(new_n224), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n227), .A2(new_n228), .ZN(new_n232));
  INV_X1    g031(.A(new_n230), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n232), .A2(new_n224), .A3(new_n223), .A4(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT11), .B(G169gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XOR2_X1   g036(.A(G113gat), .B(G141gat), .Z(new_n238));
  XOR2_X1   g037(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  OAI22_X1  g039(.A1(new_n227), .A2(new_n228), .B1(new_n211), .B2(new_n226), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n224), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n235), .A2(KEYINPUT86), .A3(new_n240), .A4(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n231), .A2(new_n234), .A3(new_n243), .A4(new_n240), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT86), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n235), .A2(new_n243), .ZN(new_n248));
  INV_X1    g047(.A(new_n240), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n244), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G15gat), .B(G43gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(G71gat), .B(G99gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT27), .B(G183gat), .ZN(new_n254));
  INV_X1    g053(.A(G190gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT28), .ZN(new_n257));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n254), .A2(new_n259), .A3(new_n255), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT26), .ZN(new_n264));
  OR3_X1    g063(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n257), .A2(new_n258), .A3(new_n260), .A4(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n258), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT24), .ZN(new_n270));
  OR2_X1    g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n258), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT65), .B(G176gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT23), .A3(new_n261), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n274), .A2(new_n276), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n266), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n268), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n266), .B1(new_n263), .B2(new_n278), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n271), .A2(new_n285), .A3(new_n258), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n269), .A2(KEYINPUT67), .A3(new_n272), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n286), .A2(new_n287), .A3(new_n279), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n277), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(G127gat), .A2(G134gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G127gat), .A2(G134gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G113gat), .B(G120gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(KEYINPUT1), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G113gat), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G120gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT1), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT68), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n305), .A3(new_n302), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n296), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n282), .A2(new_n289), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n301), .A2(new_n305), .A3(new_n302), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n305), .B1(new_n301), .B2(new_n302), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n295), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT64), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n308), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT33), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n253), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(KEYINPUT32), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n317), .B(KEYINPUT32), .C1(new_n318), .C2(new_n253), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n313), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n314), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT34), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT34), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n327), .A3(new_n315), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n321), .A2(new_n326), .A3(new_n328), .A4(new_n322), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT69), .B(KEYINPUT36), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n330), .A2(new_n331), .B1(KEYINPUT69), .B2(KEYINPUT36), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(G92gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT72), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(G64gat), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G226gat), .ZN(new_n342));
  INV_X1    g141(.A(G233gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n309), .B2(KEYINPUT29), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n290), .A2(new_n344), .ZN(new_n347));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G197gat), .B(G204gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351));
  INV_X1    g150(.A(G211gat), .ZN(new_n352));
  INV_X1    g151(.A(G218gat), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT70), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n349), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n350), .A2(new_n354), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(KEYINPUT70), .A3(new_n348), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n347), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n360), .B(KEYINPUT71), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n346), .B2(new_n347), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n341), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n344), .B1(new_n290), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n309), .A2(new_n345), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n364), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n340), .A3(new_n362), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(KEYINPUT30), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n363), .A2(new_n366), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n375), .A3(new_n340), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n379));
  XOR2_X1   g178(.A(G155gat), .B(G162gat), .Z(new_n380));
  OR2_X1    g179(.A1(KEYINPUT73), .A2(KEYINPUT2), .ZN(new_n381));
  NAND2_X1  g180(.A1(KEYINPUT73), .A2(KEYINPUT2), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G141gat), .B(G148gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386));
  INV_X1    g185(.A(G155gat), .ZN(new_n387));
  INV_X1    g186(.A(G162gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n389), .B2(KEYINPUT2), .ZN(new_n390));
  XOR2_X1   g189(.A(G141gat), .B(G148gat), .Z(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n385), .A2(new_n392), .A3(new_n295), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n393), .B1(new_n304), .B2(new_n306), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n379), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n393), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n304), .A2(new_n306), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT77), .B(new_n395), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n400));
  INV_X1    g199(.A(G141gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(G148gat), .ZN(new_n402));
  INV_X1    g201(.A(G148gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(G141gat), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n381), .B(new_n382), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n405), .A2(new_n380), .B1(new_n391), .B2(new_n390), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n406), .B(new_n295), .C1(new_n311), .C2(new_n310), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n400), .B1(new_n407), .B2(KEYINPUT4), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n396), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n310), .A2(new_n311), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT4), .B1(new_n410), .B2(new_n393), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT77), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT76), .B1(new_n407), .B2(KEYINPUT4), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n400), .A3(KEYINPUT4), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT75), .B(KEYINPUT5), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n385), .A2(new_n392), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT3), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT3), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n312), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n416), .A2(new_n417), .A3(new_n419), .A4(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT0), .B(G57gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(G85gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  AOI21_X1  g228(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n410), .A2(KEYINPUT4), .A3(new_n393), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n417), .B(new_n424), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n307), .B2(new_n406), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n312), .A2(KEYINPUT74), .A3(new_n420), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n394), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n432), .B(new_n418), .C1(new_n436), .C2(new_n417), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n425), .A2(new_n429), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n437), .ZN(new_n441));
  INV_X1    g240(.A(new_n429), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n442), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n378), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G22gat), .B(G50gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G228gat), .A2(G233gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n423), .A2(new_n368), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n364), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n357), .A2(new_n368), .A3(new_n359), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n453), .A2(KEYINPUT78), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n422), .B1(new_n453), .B2(KEYINPUT78), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n420), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n450), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n451), .A2(new_n360), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n450), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n355), .A2(new_n349), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n368), .B1(new_n358), .B2(new_n348), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n422), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n459), .B1(new_n420), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT31), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n457), .A2(new_n463), .A3(KEYINPUT31), .ZN(new_n466));
  XOR2_X1   g265(.A(G78gat), .B(G106gat), .Z(new_n467));
  NOR3_X1   g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  INV_X1    g268(.A(new_n466), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(new_n464), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n449), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n465), .B2(new_n466), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n464), .A3(new_n469), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n448), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n336), .B1(new_n447), .B2(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT81), .B(KEYINPUT38), .Z(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT82), .B(KEYINPUT37), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n340), .B1(new_n374), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT37), .B1(new_n363), .B2(new_n366), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n441), .B2(new_n442), .ZN(new_n487));
  AOI211_X1 g286(.A(KEYINPUT79), .B(new_n429), .C1(new_n425), .C2(new_n437), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n440), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n361), .B1(new_n369), .B2(new_n370), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n346), .A2(new_n347), .A3(new_n364), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT37), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n492), .A2(new_n480), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n483), .A2(new_n493), .B1(new_n374), .B2(new_n340), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(new_n494), .A3(new_n445), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT83), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n489), .A2(new_n494), .A3(new_n497), .A4(new_n445), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n485), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n436), .A2(new_n417), .ZN(new_n500));
  INV_X1    g299(.A(new_n424), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(new_n409), .B2(new_n415), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT39), .B(new_n500), .C1(new_n502), .C2(new_n417), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n413), .B1(new_n412), .B2(new_n414), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n424), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT39), .ZN(new_n507));
  INV_X1    g306(.A(new_n417), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n503), .A2(new_n509), .A3(new_n429), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT40), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n487), .B2(new_n488), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n503), .A2(new_n509), .A3(KEYINPUT40), .A4(new_n429), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n373), .A2(new_n514), .A3(new_n376), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT80), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n437), .ZN(new_n518));
  AOI211_X1 g317(.A(new_n508), .B(new_n501), .C1(new_n409), .C2(new_n415), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(new_n419), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT79), .B1(new_n520), .B2(new_n429), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n441), .A2(new_n486), .A3(new_n442), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n521), .A2(new_n522), .B1(new_n511), .B2(new_n510), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n373), .A2(new_n514), .A3(new_n376), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT80), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n476), .B1(new_n517), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n478), .B1(new_n499), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n330), .A2(new_n331), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n472), .B2(new_n475), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n446), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT35), .ZN(new_n531));
  INV_X1    g330(.A(new_n445), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n521), .A2(new_n522), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(new_n440), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n534), .A2(KEYINPUT35), .A3(new_n378), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n529), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n250), .B1(new_n527), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT21), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT9), .ZN(new_n540));
  INV_X1    g339(.A(G71gat), .ZN(new_n541));
  INV_X1    g340(.A(G78gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n543), .A2(KEYINPUT87), .ZN(new_n544));
  XOR2_X1   g343(.A(G71gat), .B(G78gat), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G57gat), .B(G64gat), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(KEYINPUT87), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n544), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n547), .A2(KEYINPUT9), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n220), .B1(new_n539), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n552), .A2(G183gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(G183gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G231gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(new_n343), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n553), .A2(G231gat), .A3(G233gat), .A4(new_n554), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G127gat), .B(G155gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT20), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n551), .A2(new_n539), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(new_n352), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(new_n561), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n562), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n566), .B1(new_n562), .B2(new_n567), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n574), .A2(G85gat), .A3(G92gat), .A4(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n573), .A2(new_n578), .B1(new_n579), .B2(KEYINPUT8), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n579), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n576), .A2(new_n580), .A3(new_n584), .A4(new_n577), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n572), .B1(new_n221), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT91), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n213), .A2(new_n222), .A3(new_n586), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G190gat), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n587), .A2(KEYINPUT91), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n587), .A2(KEYINPUT91), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n255), .B(new_n589), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(G218gat), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n255), .B1(new_n588), .B2(new_n589), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n353), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT89), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT92), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n595), .A2(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n601), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n595), .A2(new_n598), .A3(new_n607), .A4(new_n602), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n604), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G230gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(new_n343), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n586), .A2(new_n551), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n586), .A2(new_n551), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OR3_X1    g414(.A1(new_n586), .A2(new_n551), .A3(new_n613), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n611), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n614), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n611), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT93), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G120gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n403), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  INV_X1    g425(.A(new_n620), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(new_n617), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(KEYINPUT94), .B(new_n626), .C1(new_n627), .C2(new_n617), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n571), .A2(new_n609), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n538), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n444), .A2(new_n445), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(new_n215), .ZN(G1324gat));
  NOR2_X1   g436(.A1(new_n634), .A2(new_n377), .ZN(new_n638));
  NAND2_X1  g437(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n639));
  OR2_X1    g438(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n642), .A2(KEYINPUT42), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(KEYINPUT42), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n643), .B(new_n644), .C1(new_n219), .C2(new_n638), .ZN(G1325gat));
  INV_X1    g444(.A(G15gat), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n334), .A2(new_n335), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n634), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n528), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n538), .A2(new_n649), .A3(new_n633), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(new_n646), .B2(new_n650), .ZN(G1326gat));
  NOR2_X1   g450(.A1(new_n634), .A2(new_n476), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT43), .B(G22gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  NOR2_X1   g453(.A1(new_n570), .A2(new_n632), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n609), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(KEYINPUT95), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n538), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(KEYINPUT95), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n660), .A2(G29gat), .A3(new_n635), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT45), .Z(new_n662));
  XOR2_X1   g461(.A(KEYINPUT97), .B(KEYINPUT44), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n647), .B1(new_n446), .B2(new_n476), .ZN(new_n665));
  INV_X1    g464(.A(new_n485), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n497), .B1(new_n534), .B2(new_n494), .ZN(new_n667));
  INV_X1    g466(.A(new_n498), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n525), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT80), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n477), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n665), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n530), .A2(KEYINPUT35), .B1(new_n535), .B2(new_n529), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n609), .B(new_n664), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n609), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n527), .B2(new_n537), .ZN(new_n677));
  NOR2_X1   g476(.A1(KEYINPUT97), .A2(KEYINPUT44), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n248), .A2(new_n249), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n245), .A2(new_n246), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n245), .A2(new_n246), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n655), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT96), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n686), .B2(new_n635), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n662), .A2(new_n687), .ZN(G1328gat));
  NOR3_X1   g487(.A1(new_n660), .A2(G36gat), .A3(new_n377), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT46), .ZN(new_n690));
  OAI21_X1  g489(.A(G36gat), .B1(new_n686), .B2(new_n377), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(G1329gat));
  OR3_X1    g491(.A1(new_n660), .A2(G43gat), .A3(new_n528), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT98), .ZN(new_n695));
  OAI21_X1  g494(.A(G43gat), .B1(new_n686), .B2(new_n647), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n694), .A2(KEYINPUT98), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1330gat));
  OAI21_X1  g498(.A(G50gat), .B1(new_n686), .B2(new_n476), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT48), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n660), .A2(G50gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n703), .B2(new_n476), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n702), .B(new_n704), .ZN(G1331gat));
  AOI21_X1  g504(.A(new_n683), .B1(new_n527), .B2(new_n537), .ZN(new_n706));
  INV_X1    g505(.A(new_n632), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n571), .A2(new_n609), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n635), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g512(.A(new_n377), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT100), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n716), .B(new_n717), .Z(G1333gat));
  NOR3_X1   g517(.A1(new_n709), .A2(new_n541), .A3(new_n647), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT101), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n528), .B(KEYINPUT102), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n541), .B1(new_n709), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n476), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(new_n542), .ZN(G1335gat));
  NAND2_X1  g526(.A1(new_n571), .A2(new_n250), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n676), .B(new_n728), .C1(new_n527), .C2(new_n537), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT104), .B1(new_n729), .B2(KEYINPUT51), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n527), .A2(new_n537), .ZN(new_n731));
  INV_X1    g530(.A(new_n728), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(new_n609), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n731), .A2(KEYINPUT51), .A3(new_n609), .A4(new_n732), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n677), .A2(KEYINPUT103), .A3(KEYINPUT51), .A4(new_n732), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n730), .A2(new_n736), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n711), .A3(new_n632), .ZN(new_n742));
  INV_X1    g541(.A(G85gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n677), .A2(new_n678), .ZN(new_n745));
  AOI211_X1 g544(.A(new_n676), .B(new_n663), .C1(new_n527), .C2(new_n537), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n632), .B(new_n732), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n747), .A2(new_n743), .A3(new_n635), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n744), .A2(KEYINPUT105), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1336gat));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n377), .A2(G92gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n741), .A2(new_n632), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n679), .A2(new_n378), .A3(new_n632), .A4(new_n732), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(new_n757), .B2(G92gat), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(G92gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n733), .A2(new_n735), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n737), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n632), .A3(new_n755), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n754), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n756), .A2(new_n758), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n761), .A2(new_n764), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n767), .B(KEYINPUT106), .C1(new_n768), .C2(new_n760), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1337gat));
  NOR3_X1   g569(.A1(new_n707), .A2(new_n528), .A3(G99gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT107), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n741), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(G99gat), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n747), .A2(new_n647), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT108), .ZN(G1338gat));
  NOR2_X1   g576(.A1(new_n476), .A2(G106gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n741), .A2(new_n632), .A3(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n679), .A2(new_n477), .A3(new_n632), .A4(new_n732), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT53), .B1(new_n780), .B2(G106gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n780), .A2(KEYINPUT109), .A3(G106gat), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT109), .B1(new_n780), .B2(G106gat), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n763), .A2(new_n632), .A3(new_n778), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(G1339gat));
  NAND2_X1  g587(.A1(new_n711), .A2(new_n377), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n615), .A2(new_n616), .A3(new_n611), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n618), .A2(new_n792), .A3(KEYINPUT54), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(KEYINPUT54), .ZN(new_n795));
  AND2_X1   g594(.A1(KEYINPUT110), .A2(KEYINPUT54), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n617), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n797), .A3(new_n626), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n794), .A2(new_n797), .A3(KEYINPUT55), .A4(new_n626), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n800), .A2(new_n625), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n683), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n239), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n232), .A2(new_n223), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n224), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n241), .A2(new_n242), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n804), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n632), .B(new_n809), .C1(new_n681), .C2(new_n682), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n609), .B1(new_n803), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n809), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n244), .B2(new_n247), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n609), .A2(new_n813), .A3(new_n802), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n571), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n676), .A2(new_n250), .A3(new_n570), .A4(new_n707), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n791), .B1(new_n817), .B2(new_n476), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n625), .A3(new_n801), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n810), .B1(new_n250), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n676), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n609), .A2(new_n813), .A3(new_n802), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n570), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n816), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n791), .B(new_n476), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n649), .B(new_n790), .C1(new_n818), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n823), .A2(new_n824), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT111), .B1(new_n829), .B2(new_n477), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n825), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n649), .A4(new_n790), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n683), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G113gat), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n817), .A2(new_n529), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n790), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT113), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n299), .A3(new_n683), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT114), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n835), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1340gat));
  NAND3_X1  g643(.A1(new_n838), .A2(new_n297), .A3(new_n632), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n828), .A2(new_n833), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n632), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n847), .B2(new_n297), .ZN(G1341gat));
  NAND4_X1  g647(.A1(new_n828), .A2(G127gat), .A3(new_n833), .A4(new_n570), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  INV_X1    g651(.A(new_n837), .ZN(new_n853));
  AOI21_X1  g652(.A(G127gat), .B1(new_n853), .B2(new_n570), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(G1342gat));
  NAND2_X1  g654(.A1(new_n846), .A2(new_n609), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G134gat), .ZN(new_n857));
  AOI21_X1  g656(.A(G134gat), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n853), .A2(new_n609), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n861), .ZN(G1343gat));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n829), .B2(new_n476), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n817), .A2(KEYINPUT57), .A3(new_n477), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n789), .A2(new_n336), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n829), .A2(new_n476), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n401), .B1(new_n871), .B2(new_n683), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n868), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(G141gat), .A3(new_n250), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n872), .A2(KEYINPUT58), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT58), .B1(new_n872), .B2(new_n874), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1344gat));
  NAND4_X1  g676(.A1(new_n867), .A2(new_n870), .A3(new_n632), .A4(new_n868), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n879), .A3(G148gat), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT118), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n882), .A3(new_n866), .ZN(new_n883));
  OAI211_X1 g682(.A(KEYINPUT119), .B(new_n863), .C1(new_n829), .C2(new_n476), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n632), .A3(new_n868), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n879), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n632), .A2(new_n403), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n881), .A2(new_n887), .B1(new_n873), .B2(new_n888), .ZN(G1345gat));
  NAND3_X1  g688(.A1(new_n871), .A2(G155gat), .A3(new_n570), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n387), .B1(new_n873), .B2(new_n571), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(G1346gat));
  NAND3_X1  g691(.A1(new_n871), .A2(G162gat), .A3(new_n609), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n388), .B1(new_n873), .B2(new_n676), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n711), .A2(new_n377), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n831), .A2(new_n721), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n250), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n836), .A2(new_n896), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n261), .A3(new_n683), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(G1348gat));
  OAI21_X1  g701(.A(new_n262), .B1(new_n899), .B2(new_n707), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT120), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n897), .A2(new_n275), .A3(new_n707), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT121), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1349gat));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n570), .A2(new_n254), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n900), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n912), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT122), .B1(new_n899), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G183gat), .B1(new_n897), .B2(new_n571), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g718(.A1(new_n831), .A2(new_n609), .A3(new_n721), .A4(new_n896), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G190gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT123), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n923), .A3(G190gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(KEYINPUT124), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n900), .A2(new_n255), .A3(new_n609), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(KEYINPUT124), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n926), .A2(KEYINPUT124), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n922), .A2(new_n929), .A3(new_n930), .A4(new_n924), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(G1351gat));
  NAND2_X1  g731(.A1(new_n896), .A2(new_n647), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n885), .A2(new_n683), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G197gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n869), .A2(new_n934), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT125), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n683), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n936), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1352gat));
  NAND3_X1  g744(.A1(new_n885), .A2(new_n632), .A3(new_n934), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G204gat), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n937), .A2(G204gat), .A3(new_n707), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT62), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n938), .A2(new_n352), .A3(new_n570), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n883), .A2(new_n570), .A3(new_n884), .A4(new_n934), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g756(.A(KEYINPUT127), .B(new_n951), .C1(new_n953), .C2(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n938), .A2(new_n353), .A3(new_n609), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n885), .A2(new_n609), .A3(new_n934), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n353), .ZN(G1355gat));
endmodule


