//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n205), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n204), .A2(new_n216), .A3(new_n212), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n216), .B1(new_n204), .B2(new_n212), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G1gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G1gat), .B2(new_n222), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(G8gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n215), .B(KEYINPUT17), .C1(new_n217), .C2(new_n218), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n230), .B(KEYINPUT88), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n219), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n229), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT90), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n231), .B(KEYINPUT13), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n226), .A2(new_n219), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(new_n232), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(new_n233), .B2(new_n234), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT11), .ZN(new_n245));
  INV_X1    g044(.A(G169gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n240), .B(new_n243), .C1(KEYINPUT89), .C2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n239), .A3(KEYINPUT89), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n239), .A3(new_n243), .ZN(new_n252));
  INV_X1    g051(.A(new_n249), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT96), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT94), .B(G92gat), .ZN(new_n258));
  INV_X1    g057(.A(G85gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G85gat), .A2(G92gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT7), .ZN(new_n262));
  INV_X1    g061(.A(G99gat), .ZN(new_n263));
  INV_X1    g062(.A(G106gat), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT8), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT95), .ZN(new_n267));
  XOR2_X1   g066(.A(G99gat), .B(G106gat), .Z(new_n268));
  INV_X1    g067(.A(KEYINPUT95), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n260), .A2(new_n262), .A3(new_n269), .A4(new_n265), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n268), .B1(new_n267), .B2(new_n270), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n257), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n270), .ZN(new_n274));
  INV_X1    g073(.A(new_n268), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT96), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G71gat), .B(G78gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n273), .A2(new_n278), .A3(KEYINPUT10), .A4(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n283), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n271), .B2(new_n272), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(new_n277), .A3(new_n283), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT10), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G230gat), .A2(G233gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n287), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(G230gat), .A3(G233gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G120gat), .B(G148gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(G176gat), .ZN(new_n296));
  INV_X1    g095(.A(G204gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT98), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n292), .A2(new_n294), .ZN(new_n302));
  INV_X1    g101(.A(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G190gat), .B(G218gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n273), .A2(new_n278), .A3(new_n219), .ZN(new_n307));
  NAND2_X1  g106(.A1(G232gat), .A2(G233gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n308), .B(KEYINPUT93), .Z(new_n309));
  INV_X1    g108(.A(KEYINPUT41), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n221), .A2(new_n228), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(new_n273), .B2(new_n278), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n306), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT97), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n310), .ZN(new_n317));
  XNOR2_X1  g116(.A(G134gat), .B(G162gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n273), .A2(new_n278), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(new_n228), .A3(new_n221), .ZN(new_n321));
  INV_X1    g120(.A(new_n306), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n307), .A4(new_n311), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n316), .A2(new_n319), .B1(new_n315), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT97), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n315), .A2(new_n323), .A3(new_n325), .A4(new_n319), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n226), .B1(KEYINPUT21), .B2(new_n283), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT92), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n331), .B(new_n333), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n283), .A2(KEYINPUT21), .ZN(new_n335));
  NAND2_X1  g134(.A1(G231gat), .A2(G233gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G127gat), .B(G155gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT20), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n340), .ZN(new_n342));
  XNOR2_X1  g141(.A(G183gat), .B(G211gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n341), .B2(new_n342), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n334), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n347), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n331), .B(new_n332), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n345), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n305), .A2(new_n329), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT0), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G57gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(new_n259), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G141gat), .B(G148gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT2), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(G155gat), .B2(G162gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G141gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G148gat), .ZN(new_n367));
  INV_X1    g166(.A(G148gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G141gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G155gat), .B(G162gat), .ZN(new_n371));
  INV_X1    g170(.A(G155gat), .ZN(new_n372));
  INV_X1    g171(.A(G162gat), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT2), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n377));
  INV_X1    g176(.A(G127gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G134gat), .ZN(new_n379));
  INV_X1    g178(.A(G134gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G127gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT1), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(G113gat), .B2(G120gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(G113gat), .A2(G120gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI22_X1  g184(.A1(new_n379), .A2(new_n381), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G113gat), .ZN(new_n387));
  INV_X1    g186(.A(G120gat), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT1), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n380), .A2(G127gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n378), .A2(G134gat), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n389), .A2(new_n384), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n365), .A2(new_n375), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n377), .A2(KEYINPUT76), .A3(new_n393), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT5), .ZN(new_n401));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n376), .A2(new_n393), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n386), .A2(new_n392), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n408), .A2(KEYINPUT77), .A3(new_n365), .A4(new_n375), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT77), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n376), .B2(new_n393), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n406), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n407), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI211_X1 g213(.A(KEYINPUT79), .B(new_n406), .C1(new_n409), .C2(new_n411), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n404), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n365), .A2(new_n375), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT77), .B1(new_n417), .B2(new_n408), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n376), .A2(new_n393), .A3(new_n410), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT4), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT79), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n412), .A2(new_n413), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT80), .A4(new_n407), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n403), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n409), .A2(new_n411), .B1(new_n376), .B2(new_n393), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT5), .B1(new_n425), .B2(new_n402), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT78), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT78), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(KEYINPUT5), .C1(new_n425), .C2(new_n402), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n376), .A2(new_n393), .A3(new_n406), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n411), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n430), .B1(new_n431), .B2(new_n406), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n400), .A2(new_n432), .A3(new_n402), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n427), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n358), .B1(new_n424), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n403), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n420), .A2(KEYINPUT79), .B1(new_n406), .B2(new_n405), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT80), .B1(new_n437), .B2(new_n422), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n414), .A2(new_n404), .A3(new_n415), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n427), .A2(new_n429), .A3(new_n433), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n357), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n435), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n357), .B1(new_n440), .B2(new_n441), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT81), .B1(new_n445), .B2(KEYINPUT6), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT6), .B(new_n358), .C1(new_n424), .C2(new_n434), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n444), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G226gat), .ZN(new_n451));
  INV_X1    g250(.A(G233gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G169gat), .A2(G176gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT26), .ZN(new_n457));
  NOR2_X1   g256(.A1(G169gat), .A2(G176gat), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n459), .A2(new_n460), .B1(G183gat), .B2(G190gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT67), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT27), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G183gat), .ZN(new_n465));
  INV_X1    g264(.A(G183gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT27), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n463), .B1(new_n466), .B2(KEYINPUT27), .ZN(new_n469));
  INV_X1    g268(.A(G190gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n462), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n466), .A2(KEYINPUT27), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n464), .A2(G183gat), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT69), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT69), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(new_n467), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n470), .A2(KEYINPUT28), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n472), .A2(new_n480), .A3(KEYINPUT70), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT70), .B1(new_n472), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n461), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT66), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n458), .A2(KEYINPUT23), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT23), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(G169gat), .B2(G176gat), .ZN(new_n487));
  AND4_X1   g286(.A1(KEYINPUT25), .A2(new_n485), .A3(new_n455), .A4(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT24), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n466), .B2(new_n470), .ZN(new_n490));
  NAND3_X1  g289(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT65), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n466), .A2(new_n470), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n490), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n484), .B1(new_n488), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n488), .A2(new_n484), .A3(new_n496), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n485), .A2(new_n455), .A3(new_n487), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n490), .A2(new_n491), .A3(new_n495), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n498), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n454), .B1(new_n483), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n483), .A2(new_n506), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(new_n510), .B2(new_n454), .ZN(new_n511));
  AND2_X1   g310(.A1(G211gat), .A2(G218gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(G211gat), .A2(G218gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT74), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(G197gat), .ZN(new_n517));
  INV_X1    g316(.A(G197gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(KEYINPUT74), .ZN(new_n519));
  OAI21_X1  g318(.A(G204gat), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(G197gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(new_n297), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n512), .A2(KEYINPUT22), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n515), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AOI211_X1 g326(.A(new_n514), .B(new_n525), .C1(new_n520), .C2(new_n523), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G8gat), .B(G36gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G64gat), .ZN(new_n533));
  INV_X1    g332(.A(G92gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n508), .A2(new_n453), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT75), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n507), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n537), .A2(new_n539), .B1(new_n454), .B2(new_n510), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n531), .B(new_n535), .C1(new_n540), .C2(new_n530), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n535), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n540), .A2(new_n530), .ZN(new_n545));
  INV_X1    g344(.A(new_n531), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n510), .A2(new_n454), .ZN(new_n548));
  INV_X1    g347(.A(new_n539), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n507), .A2(new_n538), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n529), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n552), .A2(KEYINPUT30), .A3(new_n531), .A4(new_n535), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n543), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n450), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT82), .B(G22gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G78gat), .B(G106gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT31), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n509), .B1(new_n527), .B2(new_n528), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n417), .B1(new_n561), .B2(new_n394), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n395), .A2(new_n509), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n521), .A2(new_n522), .A3(new_n297), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n297), .B1(new_n521), .B2(new_n522), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n526), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n514), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n524), .A2(new_n515), .A3(new_n526), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n562), .A2(G50gat), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G50gat), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT29), .B1(new_n567), .B2(new_n568), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n376), .B1(new_n572), .B2(KEYINPUT3), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n529), .A2(new_n563), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n560), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G228gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(new_n452), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(G50gat), .B1(new_n562), .B2(new_n569), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n573), .A2(new_n571), .A3(new_n574), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n559), .A3(new_n581), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n576), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n579), .B1(new_n576), .B2(new_n582), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n557), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n582), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n559), .B1(new_n580), .B2(new_n581), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n578), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n576), .A2(new_n579), .A3(new_n582), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n556), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G15gat), .B(G43gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT71), .ZN(new_n592));
  XNOR2_X1  g391(.A(G71gat), .B(G99gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G227gat), .A2(G233gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n461), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT70), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n465), .A2(new_n467), .A3(new_n476), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n476), .B1(new_n465), .B2(new_n467), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n598), .A2(new_n599), .A3(new_n478), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n601));
  OAI21_X1  g400(.A(KEYINPUT67), .B1(new_n473), .B2(new_n474), .ZN(new_n602));
  AOI21_X1  g401(.A(G190gat), .B1(new_n465), .B2(new_n463), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n597), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n472), .A2(new_n480), .A3(KEYINPUT70), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n596), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n488), .A2(new_n484), .A3(new_n496), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n608), .A2(new_n497), .A3(new_n504), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n393), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n483), .A2(new_n408), .A3(new_n506), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n595), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n594), .B1(new_n612), .B2(KEYINPUT33), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT32), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n611), .ZN(new_n617));
  INV_X1    g416(.A(new_n595), .ZN(new_n618));
  AOI221_X4 g417(.A(new_n614), .B1(KEYINPUT33), .B2(new_n594), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n610), .A2(new_n595), .A3(new_n611), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT34), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT34), .A4(new_n595), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n585), .A2(new_n590), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT72), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n623), .A2(new_n627), .A3(new_n624), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n623), .B2(new_n624), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n607), .A2(new_n609), .A3(new_n393), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n408), .B1(new_n483), .B2(new_n506), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n618), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT32), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n636), .A3(new_n594), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n613), .A2(new_n615), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n630), .A2(new_n639), .A3(KEYINPUT73), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT73), .B1(new_n630), .B2(new_n639), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n626), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT35), .B1(new_n555), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT86), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(KEYINPUT86), .B(KEYINPUT35), .C1(new_n555), .C2(new_n642), .ZN(new_n646));
  INV_X1    g445(.A(new_n625), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n639), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n585), .A2(new_n590), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n648), .A2(new_n650), .A3(KEYINPUT35), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n450), .A3(new_n554), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n645), .A2(new_n646), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n555), .A2(new_n650), .ZN(new_n654));
  OAI221_X1 g453(.A(KEYINPUT36), .B1(new_n647), .B2(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT36), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n442), .A2(new_n443), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n445), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n447), .A2(new_n448), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n435), .A2(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT84), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n551), .B2(new_n529), .ZN(new_n664));
  OR3_X1    g463(.A1(new_n511), .A2(KEYINPUT85), .A3(new_n530), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT85), .B1(new_n511), .B2(new_n530), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n551), .A2(new_n663), .A3(new_n529), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT37), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n544), .A2(KEYINPUT37), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT38), .B1(new_n547), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n552), .A2(new_n531), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n673), .A2(KEYINPUT37), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n544), .B1(new_n673), .B2(KEYINPUT37), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT38), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AND4_X1   g475(.A1(new_n662), .A2(new_n672), .A3(new_n676), .A4(new_n541), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n416), .A2(new_n423), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n402), .B1(new_n678), .B2(new_n400), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT39), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n425), .B2(new_n402), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n681), .B(new_n357), .C1(new_n679), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n543), .A2(new_n547), .A3(new_n553), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n679), .A2(new_n684), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n689), .A2(KEYINPUT40), .A3(new_n357), .A4(new_n681), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n687), .A2(new_n435), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n649), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n654), .B(new_n658), .C1(new_n677), .C2(new_n692), .ZN(new_n693));
  AOI211_X1 g492(.A(new_n256), .B(new_n353), .C1(new_n653), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n662), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g495(.A1(new_n694), .A2(new_n688), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G8gat), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT16), .B(G8gat), .Z(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n702), .A2(KEYINPUT99), .A3(new_n700), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT99), .B1(new_n702), .B2(new_n700), .ZN(new_n704));
  OAI221_X1 g503(.A(new_n699), .B1(new_n700), .B2(new_n702), .C1(new_n703), .C2(new_n704), .ZN(G1325gat));
  INV_X1    g504(.A(new_n648), .ZN(new_n706));
  AOI21_X1  g505(.A(G15gat), .B1(new_n694), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT100), .ZN(new_n708));
  INV_X1    g507(.A(new_n658), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n694), .A2(G15gat), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(G1326gat));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n650), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT101), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n694), .A2(new_n716), .A3(new_n650), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT102), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n718), .A2(KEYINPUT102), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n713), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n721), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n712), .A3(new_n719), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1327gat));
  AOI21_X1  g524(.A(new_n329), .B1(new_n653), .B2(new_n693), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n301), .A2(new_n304), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n256), .A2(new_n728), .A3(new_n352), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n206), .A3(new_n662), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n653), .A2(new_n693), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n328), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n738));
  AOI211_X1 g537(.A(new_n329), .B(new_n738), .C1(new_n653), .C2(new_n693), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n730), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT104), .B1(new_n742), .B2(new_n450), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G29gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n742), .A2(KEYINPUT104), .A3(new_n450), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n733), .B1(new_n744), .B2(new_n745), .ZN(G1328gat));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747));
  AOI21_X1  g546(.A(G36gat), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n688), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n749), .B(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n207), .B1(new_n741), .B2(new_n688), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n747), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n749), .B(new_n750), .ZN(new_n755));
  INV_X1    g554(.A(new_n753), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(KEYINPUT106), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(G1329gat));
  INV_X1    g557(.A(G43gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n741), .B2(new_n709), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  NOR4_X1   g560(.A1(new_n727), .A2(G43gat), .A3(new_n648), .A4(new_n730), .ZN(new_n762));
  OR3_X1    g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1330gat));
  AOI21_X1  g564(.A(new_n571), .B1(new_n741), .B2(new_n650), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n649), .A2(G50gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n731), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OR3_X1    g569(.A1(new_n766), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n767), .B1(new_n766), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1331gat));
  AND2_X1   g572(.A1(new_n348), .A2(new_n351), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n328), .ZN(new_n775));
  AND4_X1   g574(.A1(new_n735), .A2(new_n256), .A3(new_n775), .A4(new_n728), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n662), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT107), .B(G57gat), .Z(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1332gat));
  OR2_X1    g578(.A1(new_n688), .A2(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n688), .A2(KEYINPUT108), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n776), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT49), .B(G64gat), .Z(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(G1333gat));
  NAND3_X1  g586(.A1(new_n776), .A2(G71gat), .A3(new_n709), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT109), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n776), .A2(new_n706), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n790), .A2(G71gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT50), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n789), .A2(new_n794), .A3(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1334gat));
  NAND2_X1  g595(.A1(new_n776), .A2(new_n650), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g597(.A1(new_n352), .A2(new_n255), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n727), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n305), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n259), .A3(new_n662), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n800), .A2(new_n305), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n736), .B2(new_n739), .ZN(new_n807));
  OAI21_X1  g606(.A(G85gat), .B1(new_n807), .B2(new_n450), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(G1336gat));
  XNOR2_X1  g608(.A(new_n801), .B(KEYINPUT51), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n534), .A3(new_n728), .A4(new_n783), .ZN(new_n811));
  INV_X1    g610(.A(new_n258), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n807), .B2(new_n782), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n782), .A2(G92gat), .A3(new_n305), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n802), .A2(KEYINPUT110), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n726), .A2(new_n799), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n726), .B2(new_n799), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT111), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n812), .B1(new_n807), .B2(new_n554), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n820), .A2(KEYINPUT111), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT52), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n815), .A2(new_n825), .ZN(G1337gat));
  NOR3_X1   g625(.A1(new_n807), .A2(new_n263), .A3(new_n658), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n804), .A2(new_n706), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n263), .ZN(G1338gat));
  OAI211_X1 g628(.A(new_n650), .B(new_n806), .C1(new_n736), .C2(new_n739), .ZN(new_n830));
  XOR2_X1   g629(.A(KEYINPUT112), .B(G106gat), .Z(new_n831));
  AND3_X1   g630(.A1(new_n830), .A2(KEYINPUT113), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT113), .B1(new_n830), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n305), .A2(G106gat), .A3(new_n649), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n818), .B2(new_n819), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT114), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n835), .C1(new_n818), .C2(new_n819), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT53), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n810), .B2(new_n835), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n830), .A2(new_n831), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(G1339gat));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n353), .B2(new_n255), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n775), .A2(KEYINPUT115), .A3(new_n256), .A4(new_n305), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n235), .A2(new_n239), .A3(new_n249), .A4(new_n243), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n237), .A2(new_n232), .A3(new_n236), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n237), .A2(new_n232), .A3(KEYINPUT117), .A4(new_n236), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n231), .B1(new_n229), .B2(new_n232), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n248), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n324), .A2(new_n858), .A3(new_n327), .ZN(new_n859));
  INV_X1    g658(.A(new_n291), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n284), .B2(new_n289), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n291), .B2(new_n290), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n862), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT116), .B1(new_n865), .B2(new_n303), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n867), .B(new_n298), .C1(new_n861), .C2(new_n862), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n864), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT55), .B(new_n864), .C1(new_n866), .C2(new_n868), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n859), .A2(new_n871), .A3(new_n301), .A4(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n872), .A2(new_n301), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n876), .A2(KEYINPUT118), .A3(new_n871), .A4(new_n859), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n255), .A2(new_n871), .A3(new_n301), .A4(new_n872), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n728), .A2(new_n850), .A3(new_n857), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n875), .B(new_n877), .C1(new_n880), .C2(new_n328), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n849), .B1(new_n881), .B2(new_n774), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(new_n450), .A3(new_n642), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(new_n782), .ZN(new_n884));
  AOI21_X1  g683(.A(G113gat), .B1(new_n884), .B2(new_n255), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n782), .A2(new_n662), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT119), .B1(new_n882), .B2(new_n650), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n875), .A2(new_n877), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n328), .B1(new_n878), .B2(new_n879), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n774), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n847), .A2(new_n848), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n649), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n648), .B(new_n886), .C1(new_n887), .C2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n256), .A2(new_n387), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n885), .B1(new_n895), .B2(new_n896), .ZN(G1340gat));
  AOI21_X1  g696(.A(G120gat), .B1(new_n884), .B2(new_n728), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n305), .A2(new_n388), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n895), .B2(new_n899), .ZN(G1341gat));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n378), .A3(new_n352), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n895), .A2(new_n352), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n378), .ZN(G1342gat));
  NAND4_X1  g702(.A1(new_n883), .A2(new_n380), .A3(new_n554), .A4(new_n328), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT56), .Z(new_n905));
  AND2_X1   g704(.A1(new_n895), .A2(new_n328), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n380), .ZN(G1343gat));
  NOR2_X1   g706(.A1(new_n886), .A2(new_n709), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT120), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n649), .A2(KEYINPUT57), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT57), .B1(new_n882), .B2(new_n649), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G141gat), .B1(new_n914), .B2(new_n256), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n709), .A2(new_n649), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n892), .A2(new_n662), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n783), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n366), .A3(new_n255), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT58), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT58), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n915), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1344gat));
  NAND3_X1  g723(.A1(new_n918), .A2(new_n368), .A3(new_n728), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n914), .A2(new_n305), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(KEYINPUT59), .A3(new_n368), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n928));
  INV_X1    g727(.A(new_n889), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n352), .B1(new_n929), .B2(new_n873), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n353), .A2(new_n255), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n910), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n913), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n728), .A3(new_n909), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n928), .B1(new_n934), .B2(G148gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n925), .B1(new_n927), .B2(new_n935), .ZN(G1345gat));
  OAI21_X1  g735(.A(G155gat), .B1(new_n914), .B2(new_n774), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n918), .A2(new_n372), .A3(new_n352), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1346gat));
  OAI21_X1  g738(.A(G162gat), .B1(new_n914), .B2(new_n329), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n554), .A2(new_n373), .A3(new_n328), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n917), .B2(new_n941), .ZN(G1347gat));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n882), .B2(new_n662), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n892), .A2(KEYINPUT121), .A3(new_n450), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n782), .A2(new_n642), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n255), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n887), .A2(new_n894), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n662), .A2(new_n554), .A3(new_n648), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n952), .A2(new_n246), .A3(new_n256), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n949), .A2(new_n953), .ZN(G1348gat));
  INV_X1    g753(.A(G176gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n948), .A2(new_n955), .A3(new_n728), .ZN(new_n956));
  OAI21_X1  g755(.A(G176gat), .B1(new_n952), .B2(new_n305), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1349gat));
  AOI21_X1  g757(.A(new_n893), .B1(new_n892), .B2(new_n649), .ZN(new_n959));
  AOI211_X1 g758(.A(KEYINPUT119), .B(new_n650), .C1(new_n890), .C2(new_n891), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n352), .B(new_n951), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n950), .A2(KEYINPUT123), .A3(new_n352), .A4(new_n951), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(G183gat), .A3(new_n964), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n774), .A2(new_n599), .A3(new_n598), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT121), .B1(new_n892), .B2(new_n450), .ZN(new_n967));
  AOI211_X1 g766(.A(new_n943), .B(new_n662), .C1(new_n890), .C2(new_n891), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n947), .B(new_n966), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT122), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n946), .A2(new_n971), .A3(new_n947), .A4(new_n966), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n965), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT60), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT60), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n965), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1350gat));
  NAND3_X1  g777(.A1(new_n948), .A2(new_n470), .A3(new_n328), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n950), .A2(new_n328), .A3(new_n951), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n980), .A2(new_n981), .A3(G190gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n980), .B2(G190gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(G1351gat));
  NAND2_X1  g783(.A1(new_n916), .A2(new_n783), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n985), .B1(new_n944), .B2(new_n945), .ZN(new_n986));
  XOR2_X1   g785(.A(KEYINPUT124), .B(G197gat), .Z(new_n987));
  NAND3_X1  g786(.A1(new_n986), .A2(new_n255), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n658), .A2(new_n450), .A3(new_n688), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT125), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n933), .A2(new_n255), .A3(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n992), .B2(new_n987), .ZN(G1352gat));
  NAND3_X1  g792(.A1(new_n933), .A2(new_n728), .A3(new_n990), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(G204gat), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n305), .A2(G204gat), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n986), .A2(new_n996), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n997), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT126), .B1(new_n997), .B2(KEYINPUT62), .ZN(new_n999));
  OAI221_X1 g798(.A(new_n995), .B1(KEYINPUT62), .B2(new_n997), .C1(new_n998), .C2(new_n999), .ZN(G1353gat));
  INV_X1    g799(.A(G211gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n1001), .A3(new_n352), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n989), .A2(new_n774), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n913), .A2(new_n932), .A3(new_n1003), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n1004), .A2(KEYINPUT127), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1001), .B1(new_n1004), .B2(KEYINPUT127), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n1005), .A2(KEYINPUT63), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT63), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(G1354gat));
  AOI21_X1  g808(.A(G218gat), .B1(new_n986), .B2(new_n328), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n990), .A2(G218gat), .A3(new_n328), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1010), .B1(new_n933), .B2(new_n1011), .ZN(G1355gat));
endmodule


