//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n449, new_n451, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT64), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(G567), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NOR3_X1   g036(.A1(new_n458), .A2(KEYINPUT68), .A3(new_n451), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(new_n457), .B2(G2106), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n458), .B2(new_n451), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n468), .A2(new_n470), .A3(G137), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(G101), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n468), .A2(new_n470), .A3(G125), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT69), .A4(G125), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n474), .B1(new_n480), .B2(G2105), .ZN(G160));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n468), .A2(new_n470), .A3(G2105), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n484), .B(new_n486), .C1(new_n490), .C2(G124), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n485), .A2(G138), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n500), .A3(G2104), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n471), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(new_n492), .A3(new_n493), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n496), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  NAND2_X1  g081(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(new_n511), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n518), .A2(new_n519), .B1(G651), .B2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n525), .B(new_n527), .C1(new_n528), .C2(new_n515), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n511), .A2(G89), .A3(new_n512), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT74), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n533), .A2(G651), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n513), .ZN(new_n536));
  INV_X1    g111(.A(new_n515), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT75), .B(G52), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n536), .A2(G90), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n513), .A2(new_n545), .B1(new_n515), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT76), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n550), .A2(new_n554), .ZN(G188));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n515), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n536), .A2(G91), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n559), .B(new_n560), .C1(new_n543), .C2(new_n561), .ZN(G299));
  OR2_X1    g137(.A1(G168), .A2(KEYINPUT77), .ZN(new_n563));
  NAND2_X1  g138(.A1(G168), .A2(KEYINPUT77), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  OR2_X1    g141(.A1(new_n511), .A2(G74), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n567), .A2(G651), .B1(new_n537), .B2(G49), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n513), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n536), .A2(KEYINPUT78), .A3(G87), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(G288));
  AND3_X1   g148(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n521), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n574), .B1(new_n577), .B2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n536), .A2(G86), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT79), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT80), .B(G85), .ZN(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n513), .A2(new_n585), .B1(new_n515), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n584), .A2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n521), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n537), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT10), .B1(new_n513), .B2(new_n595), .ZN(new_n596));
  OR3_X1    g171(.A1(new_n513), .A2(KEYINPUT10), .A3(new_n595), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G171), .B2(new_n599), .ZN(G284));
  OAI21_X1  g176(.A(new_n600), .B1(G171), .B2(new_n599), .ZN(G321));
  NAND2_X1  g177(.A1(G299), .A2(new_n599), .ZN(new_n603));
  INV_X1    g178(.A(G286), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n599), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n599), .ZN(G280));
  INV_X1    g181(.A(new_n598), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NOR2_X1   g184(.A1(new_n598), .A2(G559), .ZN(new_n610));
  OR3_X1    g185(.A1(new_n610), .A2(KEYINPUT82), .A3(new_n599), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT82), .B1(new_n610), .B2(new_n599), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n611), .B(new_n612), .C1(G868), .C2(new_n548), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g189(.A1(new_n490), .A2(G123), .B1(G135), .B2(new_n485), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n471), .A2(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT15), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2435), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(G2435), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(KEYINPUT14), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2443), .B(G2446), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n634), .A2(new_n636), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n626), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n641), .A2(new_n637), .A3(new_n625), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n640), .A2(new_n642), .A3(G14), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n648), .A2(KEYINPUT83), .ZN(new_n649));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(new_n647), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n646), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT84), .Z(new_n654));
  XOR2_X1   g229(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n647), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n654), .B1(new_n656), .B2(new_n650), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n645), .A3(new_n650), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n646), .A2(new_n648), .A3(new_n650), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n672), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT88), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n671), .B(new_n674), .C1(new_n666), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  INV_X1    g255(.A(G1981), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  MUX2_X1   g260(.A(G24), .B(G290), .S(G16), .Z(new_n686));
  XOR2_X1   g261(.A(KEYINPUT90), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  AOI22_X1  g263(.A1(new_n490), .A2(G119), .B1(G131), .B2(new_n485), .ZN(new_n689));
  OR2_X1    g264(.A1(G95), .A2(G2105), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n690), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT89), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(G25), .B(new_n693), .S(G29), .Z(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT35), .B(G1991), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(G16), .A2(G23), .ZN(new_n698));
  INV_X1    g273(.A(G288), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT33), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n700), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G6), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n580), .B2(new_n705), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(G166), .A2(G16), .ZN(new_n710));
  OR2_X1    g285(.A1(G16), .A2(G22), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G1971), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n710), .A2(G1971), .A3(new_n711), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n704), .A2(new_n709), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT91), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(KEYINPUT91), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n719), .B1(new_n717), .B2(new_n718), .ZN(new_n722));
  OAI211_X1 g297(.A(KEYINPUT95), .B(new_n697), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G21), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G168), .B2(G16), .ZN(new_n728));
  INV_X1    g303(.A(G1966), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G27), .A2(G29), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G164), .B2(G29), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT30), .B(G28), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n732), .A2(G2078), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n548), .A2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G16), .B2(G19), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT96), .B(G1341), .Z(new_n738));
  OAI211_X1 g313(.A(new_n730), .B(new_n735), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G4), .A2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n607), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(G1348), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G2078), .B2(new_n732), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n739), .B(new_n744), .C1(new_n737), .C2(new_n738), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n490), .A2(G129), .B1(G141), .B2(new_n485), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n746), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G29), .B2(G32), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  OR2_X1    g330(.A1(KEYINPUT24), .A2(G34), .ZN(new_n756));
  NAND2_X1  g331(.A1(KEYINPUT24), .A2(G34), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n756), .A2(new_n733), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G160), .B2(new_n733), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n754), .A2(new_n755), .B1(G2084), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n733), .A2(G33), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n468), .A2(new_n470), .A3(G127), .ZN(new_n762));
  INV_X1    g337(.A(G115), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n467), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n764), .A2(G2105), .B1(G139), .B2(new_n485), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n761), .B1(new_n769), .B2(new_n733), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G2072), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n760), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT99), .ZN(new_n773));
  NAND2_X1  g348(.A1(G171), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G5), .B2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G1961), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT100), .Z(new_n778));
  NAND3_X1  g353(.A1(new_n745), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G29), .A2(G35), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G162), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT29), .B(G2090), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT23), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n705), .A2(G20), .ZN(new_n785));
  AOI22_X1  g360(.A1(G299), .A2(G16), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n733), .A2(G26), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n490), .A2(G128), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT97), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n471), .A2(G116), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n485), .A2(G140), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT97), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n490), .A2(new_n796), .A3(G128), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n791), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n789), .B1(new_n799), .B2(new_n733), .ZN(new_n800));
  MUX2_X1   g375(.A(new_n789), .B(new_n800), .S(KEYINPUT28), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2067), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n779), .A2(new_n783), .A3(new_n788), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n723), .A2(new_n724), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n697), .B1(new_n721), .B2(new_n722), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT36), .B1(new_n805), .B2(new_n724), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n726), .B(new_n803), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  OAI22_X1  g382(.A1(new_n754), .A2(new_n755), .B1(G2084), .B2(new_n759), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n776), .B2(new_n775), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT101), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n618), .A2(new_n733), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT31), .B(G11), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n807), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(G311));
  INV_X1    g389(.A(new_n807), .ZN(new_n815));
  INV_X1    g390(.A(new_n810), .ZN(new_n816));
  INV_X1    g391(.A(new_n811), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n812), .ZN(G150));
  AOI22_X1  g393(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n543), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n513), .A2(new_n821), .B1(new_n515), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n607), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n825), .A2(new_n548), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n824), .B1(new_n544), .B2(new_n547), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT39), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n829), .B(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n827), .B1(new_n834), .B2(G860), .ZN(G145));
  INV_X1    g410(.A(G37), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n618), .B(G160), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G162), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n621), .B1(new_n689), .B2(new_n692), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n490), .A2(G130), .B1(G142), .B2(new_n485), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(G118), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(G2105), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n689), .A2(new_n621), .A3(new_n692), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n840), .A2(new_n841), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n841), .A2(new_n845), .ZN(new_n848));
  INV_X1    g423(.A(new_n846), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(new_n839), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT102), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n847), .A2(new_n850), .A3(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n752), .A2(new_n768), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n751), .A2(new_n769), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n798), .A2(G164), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n791), .A2(new_n505), .A3(new_n795), .A4(new_n797), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n855), .A2(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n838), .B1(new_n854), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n847), .A2(new_n850), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n861), .A2(new_n862), .ZN(new_n867));
  INV_X1    g442(.A(new_n853), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n851), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT103), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT104), .B1(new_n854), .B2(new_n863), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n854), .A2(new_n863), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n870), .A2(new_n871), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n876), .A2(new_n877), .A3(new_n838), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n876), .B2(new_n838), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n836), .B(new_n866), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT106), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n838), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT105), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n876), .A2(new_n877), .A3(new_n838), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n836), .A4(new_n866), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n881), .A2(new_n887), .A3(KEYINPUT40), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT40), .B1(new_n881), .B2(new_n887), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(G395));
  NAND2_X1  g465(.A1(G303), .A2(G290), .ZN(new_n891));
  NAND3_X1  g466(.A1(G166), .A2(new_n589), .A3(new_n584), .ZN(new_n892));
  AOI21_X1  g467(.A(G305), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n892), .A3(G305), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n894), .A2(new_n699), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n699), .B1(new_n894), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT42), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n832), .B(KEYINPUT107), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(new_n610), .Z(new_n901));
  OR2_X1    g476(.A1(G299), .A2(new_n598), .ZN(new_n902));
  NAND2_X1  g477(.A1(G299), .A2(new_n598), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n901), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n903), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n909), .B2(new_n901), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n899), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n899), .A2(new_n910), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n599), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n824), .A2(G868), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n913), .A2(KEYINPUT108), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT108), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(G295));
  OR2_X1    g492(.A1(new_n913), .A2(new_n914), .ZN(G331));
  NAND2_X1  g493(.A1(G301), .A2(G168), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n832), .B(new_n919), .C1(new_n604), .C2(G301), .ZN(new_n920));
  AOI21_X1  g495(.A(G301), .B1(new_n563), .B2(new_n564), .ZN(new_n921));
  INV_X1    g496(.A(new_n919), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n830), .B(new_n831), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n908), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n920), .A2(new_n923), .A3(new_n925), .A4(new_n905), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n906), .A2(new_n904), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n923), .A4(new_n920), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n920), .A2(new_n923), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n909), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(KEYINPUT111), .A3(new_n909), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n931), .A2(new_n898), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n935), .A2(new_n936), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n940), .A2(KEYINPUT112), .A3(new_n898), .A4(new_n931), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n898), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(new_n926), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n942), .A2(KEYINPUT113), .A3(new_n836), .A4(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n939), .A2(new_n941), .A3(new_n945), .A4(new_n836), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(KEYINPUT43), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n931), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n935), .A2(new_n936), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n939), .A2(new_n941), .A3(new_n836), .A4(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(KEYINPUT44), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n942), .A2(new_n957), .A3(new_n836), .A4(new_n945), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n505), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(G160), .A2(G40), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(G1996), .A3(new_n751), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT114), .Z(new_n971));
  INV_X1    g546(.A(G2067), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n799), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n798), .A2(G2067), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n973), .B(new_n974), .C1(G1996), .C2(new_n751), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n971), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n693), .A2(new_n695), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n693), .A2(new_n695), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n969), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(G290), .B(G1986), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n969), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n976), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n967), .A2(KEYINPUT115), .ZN(new_n984));
  INV_X1    g559(.A(G40), .ZN(new_n985));
  AOI211_X1 g560(.A(new_n985), .B(new_n474), .C1(new_n480), .C2(G2105), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n965), .A2(new_n990), .A3(new_n966), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n984), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n505), .A2(new_n993), .A3(new_n964), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n505), .B2(new_n964), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n986), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT58), .B(G1341), .Z(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT122), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT122), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n992), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT59), .B1(new_n1003), .B2(new_n548), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n992), .A2(new_n1001), .A3(new_n998), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1001), .B1(new_n992), .B2(new_n998), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT59), .B(new_n548), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n965), .A2(KEYINPUT116), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n505), .A2(new_n993), .A3(new_n964), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n965), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n986), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1956), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT57), .B1(new_n559), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(G299), .B(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT56), .B(G2072), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n984), .A2(new_n988), .A3(new_n991), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT121), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1022), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1019), .A2(KEYINPUT121), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT61), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n984), .A2(new_n988), .A3(new_n991), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1036), .A2(new_n1023), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1033), .B1(new_n1037), .B2(new_n1022), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1012), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n986), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n742), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n972), .B(new_n986), .C1(new_n994), .C2(new_n995), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(KEYINPUT60), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT60), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(new_n598), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(KEYINPUT60), .A3(new_n607), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1030), .A2(new_n1038), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1009), .A2(new_n1034), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT123), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1030), .B1(new_n598), .B2(new_n1046), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1050), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1012), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n994), .B2(new_n995), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n968), .B1(KEYINPUT50), .B2(new_n965), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1059), .A2(G2090), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1035), .A2(new_n713), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1055), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G166), .A2(new_n1055), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT55), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n580), .A2(new_n681), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT118), .B(G86), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n578), .B1(new_n513), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G1981), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT49), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n996), .A2(G8), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1066), .A2(new_n1069), .A3(KEYINPUT49), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n996), .B(G8), .C1(new_n1076), .C2(G288), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT52), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n699), .A2(G1976), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1077), .A2(KEYINPUT52), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1017), .A2(G2090), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1055), .B1(new_n1083), .B2(new_n1061), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1065), .B(new_n1082), .C1(new_n1064), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1035), .A2(G2078), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1087), .A2(new_n1088), .B1(new_n776), .B2(new_n1059), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT45), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n986), .A2(new_n987), .ZN(new_n1091));
  OR4_X1    g666(.A1(new_n1088), .A2(new_n1090), .A3(G2078), .A4(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(G301), .A3(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT124), .B(G2078), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n988), .A2(KEYINPUT53), .A3(new_n967), .A4(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(KEYINPUT54), .B(new_n1093), .C1(new_n1096), .C2(G301), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1089), .A2(G301), .A3(new_n1095), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n729), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1103));
  INV_X1    g678(.A(G2084), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1057), .A2(new_n1058), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(G168), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1102), .B1(new_n1106), .B2(G8), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(G168), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1109));
  OAI211_X1 g684(.A(G8), .B(new_n1106), .C1(new_n1109), .C2(new_n1102), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1086), .A2(new_n1097), .A3(new_n1101), .A4(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1053), .A2(new_n1054), .A3(new_n1112), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1065), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1065), .A2(new_n1082), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1055), .B(G286), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT63), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1075), .A2(new_n1076), .A3(new_n699), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1066), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1073), .B(KEYINPUT119), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1126));
  INV_X1    g701(.A(G168), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1102), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1106), .A2(G8), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT62), .B1(new_n1130), .B2(new_n1107), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1108), .A2(new_n1110), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(new_n1100), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1117), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1115), .B(new_n1125), .C1(new_n1137), .C2(new_n1085), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n983), .B1(new_n1113), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n969), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n976), .A2(new_n978), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(new_n973), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1140), .A2(G1986), .A3(G290), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n1144));
  XOR2_X1   g719(.A(new_n1143), .B(new_n1144), .Z(new_n1145));
  AND3_X1   g720(.A1(new_n1145), .A2(new_n976), .A3(new_n979), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n969), .A2(new_n989), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT46), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n973), .A2(new_n752), .A3(new_n974), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1140), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT47), .Z(new_n1151));
  NOR3_X1   g726(.A1(new_n1142), .A2(new_n1146), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1139), .A2(KEYINPUT126), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT123), .ZN(new_n1156));
  AND4_X1   g731(.A1(new_n1086), .A2(new_n1097), .A3(new_n1101), .A4(new_n1111), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1085), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1160), .A2(new_n1114), .A3(new_n1124), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n982), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1152), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1154), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1153), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g740(.A1(new_n881), .A2(new_n887), .ZN(new_n1167));
  NOR2_X1   g741(.A1(G227), .A2(new_n465), .ZN(new_n1168));
  AND3_X1   g742(.A1(new_n643), .A2(KEYINPUT127), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g743(.A(KEYINPUT127), .B1(new_n643), .B2(new_n1168), .ZN(new_n1170));
  OR2_X1    g744(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AND2_X1   g745(.A1(new_n1171), .A2(new_n684), .ZN(new_n1172));
  AND3_X1   g746(.A1(new_n1167), .A2(new_n1172), .A3(new_n960), .ZN(G308));
  NAND4_X1  g747(.A1(new_n1167), .A2(new_n684), .A3(new_n960), .A4(new_n1171), .ZN(G225));
endmodule


