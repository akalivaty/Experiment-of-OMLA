

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596;

  XNOR2_X1 U326 ( .A(n336), .B(n335), .ZN(n339) );
  XNOR2_X1 U327 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U328 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n474) );
  NOR2_X1 U329 ( .A1(n532), .A2(n531), .ZN(n456) );
  XNOR2_X1 U330 ( .A(n343), .B(n342), .ZN(n346) );
  INV_X1 U331 ( .A(KEYINPUT83), .ZN(n340) );
  XNOR2_X1 U332 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U333 ( .A(n560), .B(KEYINPUT80), .ZN(n571) );
  XNOR2_X1 U334 ( .A(n477), .B(KEYINPUT38), .ZN(n506) );
  XNOR2_X1 U335 ( .A(n326), .B(n294), .ZN(n327) );
  XOR2_X1 U336 ( .A(n325), .B(n324), .Z(n294) );
  XOR2_X1 U337 ( .A(n438), .B(G64GAT), .Z(n295) );
  XOR2_X1 U338 ( .A(n375), .B(n374), .Z(n296) );
  XNOR2_X1 U339 ( .A(n367), .B(KEYINPUT46), .ZN(n368) );
  XNOR2_X1 U340 ( .A(n369), .B(n368), .ZN(n370) );
  INV_X1 U341 ( .A(KEYINPUT15), .ZN(n333) );
  XNOR2_X1 U342 ( .A(n334), .B(n333), .ZN(n335) );
  INV_X1 U343 ( .A(KEYINPUT66), .ZN(n378) );
  XNOR2_X1 U344 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U345 ( .A(n341), .B(n340), .ZN(n342) );
  INV_X1 U346 ( .A(KEYINPUT95), .ZN(n469) );
  XNOR2_X1 U347 ( .A(n360), .B(n359), .ZN(n365) );
  NOR2_X1 U348 ( .A1(n419), .A2(n520), .ZN(n579) );
  XNOR2_X1 U349 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n366) );
  XNOR2_X1 U350 ( .A(n470), .B(n469), .ZN(n484) );
  XNOR2_X1 U351 ( .A(n476), .B(n366), .ZN(n551) );
  XNOR2_X1 U352 ( .A(n475), .B(n474), .ZN(n519) );
  XNOR2_X1 U353 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U354 ( .A(KEYINPUT122), .B(n580), .Z(n593) );
  XNOR2_X1 U355 ( .A(n348), .B(n347), .ZN(n588) );
  INV_X1 U356 ( .A(G43GAT), .ZN(n478) );
  XOR2_X1 U357 ( .A(KEYINPUT90), .B(n465), .Z(n520) );
  XNOR2_X1 U358 ( .A(n453), .B(G169GAT), .ZN(n454) );
  XNOR2_X1 U359 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U360 ( .A(n455), .B(n454), .ZN(G1348GAT) );
  XNOR2_X1 U361 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  XOR2_X1 U362 ( .A(KEYINPUT73), .B(KEYINPUT30), .Z(n298) );
  XNOR2_X1 U363 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n297) );
  XNOR2_X1 U364 ( .A(n298), .B(n297), .ZN(n304) );
  XOR2_X1 U365 ( .A(G15GAT), .B(KEYINPUT71), .Z(n344) );
  XOR2_X1 U366 ( .A(n344), .B(G29GAT), .Z(n302) );
  XOR2_X1 U367 ( .A(KEYINPUT8), .B(G43GAT), .Z(n300) );
  XNOR2_X1 U368 ( .A(KEYINPUT70), .B(KEYINPUT7), .ZN(n299) );
  XNOR2_X1 U369 ( .A(n300), .B(n299), .ZN(n377) );
  XNOR2_X1 U370 ( .A(n377), .B(G50GAT), .ZN(n301) );
  XNOR2_X1 U371 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U372 ( .A(n304), .B(n303), .ZN(n317) );
  XOR2_X1 U373 ( .A(G22GAT), .B(G113GAT), .Z(n306) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(G36GAT), .ZN(n305) );
  XNOR2_X1 U375 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U376 ( .A(G8GAT), .B(G1GAT), .Z(n308) );
  XNOR2_X1 U377 ( .A(G141GAT), .B(G197GAT), .ZN(n307) );
  XNOR2_X1 U378 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U379 ( .A(n310), .B(n309), .Z(n315) );
  XOR2_X1 U380 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n312) );
  NAND2_X1 U381 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U382 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U383 ( .A(KEYINPUT72), .B(n313), .ZN(n314) );
  XNOR2_X1 U384 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U385 ( .A(n317), .B(n316), .ZN(n534) );
  INV_X1 U386 ( .A(KEYINPUT54), .ZN(n399) );
  XOR2_X1 U387 ( .A(G36GAT), .B(G190GAT), .Z(n375) );
  XOR2_X1 U388 ( .A(G176GAT), .B(G204GAT), .Z(n356) );
  XNOR2_X1 U389 ( .A(n375), .B(n356), .ZN(n330) );
  XOR2_X1 U390 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n319) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n318) );
  XNOR2_X1 U392 ( .A(n319), .B(n318), .ZN(n438) );
  NAND2_X1 U393 ( .A1(G226GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U394 ( .A(n295), .B(n320), .ZN(n328) );
  XOR2_X1 U395 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n322) );
  XNOR2_X1 U396 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n321) );
  XNOR2_X1 U397 ( .A(n322), .B(n321), .ZN(n423) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G183GAT), .ZN(n323) );
  XNOR2_X1 U399 ( .A(n323), .B(G211GAT), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n423), .B(n336), .ZN(n326) );
  XOR2_X1 U401 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n325) );
  XNOR2_X1 U402 ( .A(G218GAT), .B(G92GAT), .ZN(n324) );
  XNOR2_X1 U403 ( .A(n330), .B(n329), .ZN(n492) );
  XOR2_X1 U404 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n332) );
  XNOR2_X1 U405 ( .A(KEYINPUT12), .B(KEYINPUT82), .ZN(n331) );
  XNOR2_X1 U406 ( .A(n332), .B(n331), .ZN(n348) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XOR2_X1 U408 ( .A(KEYINPUT13), .B(G64GAT), .Z(n338) );
  XNOR2_X1 U409 ( .A(G71GAT), .B(G78GAT), .ZN(n337) );
  XNOR2_X1 U410 ( .A(n338), .B(n337), .ZN(n353) );
  XOR2_X1 U411 ( .A(n339), .B(n353), .Z(n343) );
  XOR2_X1 U412 ( .A(G22GAT), .B(G155GAT), .Z(n422) );
  XOR2_X1 U413 ( .A(G1GAT), .B(G127GAT), .Z(n410) );
  XNOR2_X1 U414 ( .A(n422), .B(n410), .ZN(n341) );
  XNOR2_X1 U415 ( .A(n344), .B(G57GAT), .ZN(n345) );
  XNOR2_X1 U416 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U417 ( .A(KEYINPUT110), .B(n588), .ZN(n567) );
  XOR2_X1 U418 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n350) );
  NAND2_X1 U419 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U420 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U421 ( .A(n351), .B(KEYINPUT31), .Z(n355) );
  XNOR2_X1 U422 ( .A(G120GAT), .B(G148GAT), .ZN(n352) );
  XNOR2_X1 U423 ( .A(n352), .B(G57GAT), .ZN(n404) );
  XNOR2_X1 U424 ( .A(n404), .B(n353), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n355), .B(n354), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n356), .B(KEYINPUT76), .ZN(n358) );
  INV_X1 U427 ( .A(KEYINPUT74), .ZN(n357) );
  XOR2_X1 U428 ( .A(KEYINPUT75), .B(G92GAT), .Z(n362) );
  XNOR2_X1 U429 ( .A(G99GAT), .B(G106GAT), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U431 ( .A(G85GAT), .B(n363), .Z(n382) );
  INV_X1 U432 ( .A(n382), .ZN(n364) );
  XOR2_X1 U433 ( .A(n365), .B(n364), .Z(n584) );
  INV_X1 U434 ( .A(n584), .ZN(n476) );
  INV_X1 U435 ( .A(n534), .ZN(n581) );
  AND2_X1 U436 ( .A1(n551), .A2(n581), .ZN(n369) );
  INV_X1 U437 ( .A(KEYINPUT111), .ZN(n367) );
  NOR2_X1 U438 ( .A1(n567), .A2(n370), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n371), .B(KEYINPUT112), .ZN(n389) );
  XOR2_X1 U440 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n373) );
  XNOR2_X1 U441 ( .A(KEYINPUT78), .B(KEYINPUT11), .ZN(n372) );
  XNOR2_X1 U442 ( .A(n373), .B(n372), .ZN(n374) );
  NAND2_X1 U443 ( .A1(G232GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n296), .B(n376), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n377), .B(KEYINPUT10), .ZN(n379) );
  XOR2_X1 U446 ( .A(n383), .B(n382), .Z(n388) );
  XOR2_X1 U447 ( .A(G162GAT), .B(KEYINPUT77), .Z(n385) );
  XNOR2_X1 U448 ( .A(G50GAT), .B(G218GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n431) );
  XNOR2_X1 U450 ( .A(G29GAT), .B(G134GAT), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n386), .B(KEYINPUT79), .ZN(n416) );
  XNOR2_X1 U452 ( .A(n431), .B(n416), .ZN(n387) );
  XNOR2_X1 U453 ( .A(n388), .B(n387), .ZN(n560) );
  NAND2_X1 U454 ( .A1(n389), .A2(n560), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n390), .B(KEYINPUT47), .ZN(n396) );
  INV_X1 U456 ( .A(n588), .ZN(n471) );
  XNOR2_X1 U457 ( .A(KEYINPUT36), .B(KEYINPUT100), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n391), .B(n571), .ZN(n591) );
  NOR2_X1 U459 ( .A1(n471), .A2(n591), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n392), .B(KEYINPUT45), .ZN(n393) );
  NAND2_X1 U461 ( .A1(n393), .A2(n476), .ZN(n394) );
  NOR2_X1 U462 ( .A1(n581), .A2(n394), .ZN(n395) );
  NOR2_X1 U463 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n397), .B(KEYINPUT48), .ZN(n548) );
  NOR2_X1 U465 ( .A1(n492), .A2(n548), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n419) );
  XOR2_X1 U467 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n401) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U470 ( .A(n402), .B(KEYINPUT88), .Z(n406) );
  XNOR2_X1 U471 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n403), .B(KEYINPUT3), .ZN(n430) );
  XNOR2_X1 U473 ( .A(n430), .B(n404), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n406), .B(n405), .ZN(n414) );
  XOR2_X1 U475 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n408) );
  XNOR2_X1 U476 ( .A(G155GAT), .B(KEYINPUT89), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U478 ( .A(n409), .B(G85GAT), .Z(n412) );
  XNOR2_X1 U479 ( .A(G162GAT), .B(n410), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U481 ( .A(n414), .B(n413), .Z(n418) );
  XNOR2_X1 U482 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n415) );
  XOR2_X1 U483 ( .A(n415), .B(KEYINPUT85), .Z(n437) );
  XOR2_X1 U484 ( .A(n437), .B(n416), .Z(n417) );
  XNOR2_X1 U485 ( .A(n418), .B(n417), .ZN(n465) );
  XOR2_X1 U486 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n421) );
  XNOR2_X1 U487 ( .A(G106GAT), .B(KEYINPUT23), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n421), .B(n420), .ZN(n435) );
  XOR2_X1 U489 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U492 ( .A(G78GAT), .B(G148GAT), .Z(n427) );
  XNOR2_X1 U493 ( .A(G211GAT), .B(G204GAT), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U495 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U496 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n435), .B(n434), .ZN(n461) );
  NAND2_X1 U499 ( .A1(n579), .A2(n461), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n436), .B(KEYINPUT55), .ZN(n452) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n451) );
  XOR2_X1 U502 ( .A(G120GAT), .B(G71GAT), .Z(n440) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U505 ( .A(G176GAT), .B(G127GAT), .Z(n442) );
  XNOR2_X1 U506 ( .A(KEYINPUT20), .B(G183GAT), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U508 ( .A(n444), .B(n443), .Z(n449) );
  XOR2_X1 U509 ( .A(G190GAT), .B(G134GAT), .Z(n446) );
  XNOR2_X1 U510 ( .A(G43GAT), .B(G99GAT), .ZN(n445) );
  XNOR2_X1 U511 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U512 ( .A(G15GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U513 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U514 ( .A(n451), .B(n450), .ZN(n532) );
  NAND2_X1 U515 ( .A1(n452), .A2(n532), .ZN(n570) );
  NOR2_X1 U516 ( .A1(n534), .A2(n570), .ZN(n455) );
  XNOR2_X1 U517 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n453) );
  XOR2_X1 U518 ( .A(n492), .B(KEYINPUT27), .Z(n459) );
  AND2_X1 U519 ( .A1(n520), .A2(n459), .ZN(n546) );
  XNOR2_X1 U520 ( .A(KEYINPUT28), .B(n461), .ZN(n505) );
  NAND2_X1 U521 ( .A1(n546), .A2(n505), .ZN(n531) );
  XNOR2_X1 U522 ( .A(KEYINPUT93), .B(n456), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n532), .A2(n461), .ZN(n458) );
  XNOR2_X1 U524 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n457) );
  XNOR2_X1 U525 ( .A(n458), .B(n457), .ZN(n578) );
  NAND2_X1 U526 ( .A1(n459), .A2(n578), .ZN(n464) );
  INV_X1 U527 ( .A(n492), .ZN(n522) );
  NAND2_X1 U528 ( .A1(n532), .A2(n522), .ZN(n460) );
  NAND2_X1 U529 ( .A1(n461), .A2(n460), .ZN(n462) );
  XOR2_X1 U530 ( .A(KEYINPUT25), .B(n462), .Z(n463) );
  NAND2_X1 U531 ( .A1(n464), .A2(n463), .ZN(n466) );
  NAND2_X1 U532 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U533 ( .A1(n468), .A2(n467), .ZN(n470) );
  AND2_X1 U534 ( .A1(n484), .A2(n471), .ZN(n472) );
  XNOR2_X1 U535 ( .A(n472), .B(KEYINPUT101), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n591), .A2(n473), .ZN(n475) );
  NAND2_X1 U537 ( .A1(n476), .A2(n581), .ZN(n486) );
  NOR2_X1 U538 ( .A1(n519), .A2(n486), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n506), .A2(n532), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n479) );
  XOR2_X1 U541 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n483) );
  NAND2_X1 U542 ( .A1(n588), .A2(n571), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(n485) );
  NAND2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n508) );
  NOR2_X1 U545 ( .A1(n486), .A2(n508), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT96), .B(n487), .Z(n497) );
  INV_X1 U547 ( .A(n520), .ZN(n488) );
  NOR2_X1 U548 ( .A1(n497), .A2(n488), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NOR2_X1 U552 ( .A1(n492), .A2(n497), .ZN(n493) );
  XOR2_X1 U553 ( .A(G8GAT), .B(n493), .Z(G1325GAT) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n496) );
  INV_X1 U555 ( .A(n532), .ZN(n494) );
  NOR2_X1 U556 ( .A1(n494), .A2(n497), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n505), .A2(n497), .ZN(n498) );
  XOR2_X1 U559 ( .A(KEYINPUT98), .B(n498), .Z(n499) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n499), .ZN(G1327GAT) );
  NAND2_X1 U561 ( .A1(n506), .A2(n520), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT99), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  XOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT103), .Z(n504) );
  NAND2_X1 U566 ( .A1(n506), .A2(n522), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  INV_X1 U568 ( .A(n505), .ZN(n526) );
  NAND2_X1 U569 ( .A1(n506), .A2(n526), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n507), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n510) );
  XOR2_X1 U572 ( .A(n551), .B(KEYINPUT106), .Z(n562) );
  OR2_X1 U573 ( .A1(n581), .A2(n562), .ZN(n518) );
  NOR2_X1 U574 ( .A1(n518), .A2(n508), .ZN(n515) );
  NAND2_X1 U575 ( .A1(n515), .A2(n520), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  XOR2_X1 U578 ( .A(G64GAT), .B(KEYINPUT107), .Z(n513) );
  NAND2_X1 U579 ( .A1(n515), .A2(n522), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n532), .A2(n515), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n514), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U584 ( .A1(n515), .A2(n526), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n527), .A2(n520), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n522), .A2(n527), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n532), .A2(n527), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n524), .B(KEYINPUT108), .ZN(n525) );
  XNOR2_X1 U593 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n529) );
  NAND2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n548), .A2(n531), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n542) );
  NOR2_X1 U600 ( .A1(n534), .A2(n542), .ZN(n535) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n535), .Z(G1340GAT) );
  NOR2_X1 U602 ( .A1(n562), .A2(n542), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U605 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  INV_X1 U606 ( .A(n542), .ZN(n539) );
  NAND2_X1 U607 ( .A1(n539), .A2(n567), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  NOR2_X1 U610 ( .A1(n571), .A2(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(KEYINPUT114), .B(KEYINPUT51), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n545), .ZN(G1343GAT) );
  XOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT115), .Z(n550) );
  NAND2_X1 U615 ( .A1(n578), .A2(n546), .ZN(n547) );
  NOR2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n558), .A2(n581), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n553) );
  NAND2_X1 U621 ( .A1(n558), .A2(n551), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT117), .Z(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n588), .ZN(n556) );
  XNOR2_X1 U626 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  INV_X1 U627 ( .A(n558), .ZN(n559) );
  NOR2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NOR2_X1 U630 ( .A1(n562), .A2(n570), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  INV_X1 U635 ( .A(n570), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT121), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n576) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U645 ( .A(KEYINPUT123), .B(n577), .Z(n583) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n593), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n584), .A2(n593), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(G204GAT), .B(n587), .Z(G1353GAT) );
  NAND2_X1 U653 ( .A1(n593), .A2(n588), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(KEYINPUT126), .ZN(n590) );
  XNOR2_X1 U655 ( .A(G211GAT), .B(n590), .ZN(G1354GAT) );
  INV_X1 U656 ( .A(n591), .ZN(n592) );
  AND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U658 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n596), .B(G218GAT), .ZN(G1355GAT) );
endmodule

