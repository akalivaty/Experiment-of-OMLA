//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n205), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n216));
  AND3_X1   g0016(.A1(new_n215), .A2(G50), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT66), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G20), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT64), .Z(new_n223));
  AOI22_X1  g0023(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G50), .ZN(new_n228));
  INV_X1    g0028(.A(G226), .ZN(new_n229));
  INV_X1    g0029(.A(G77), .ZN(new_n230));
  INV_X1    g0030(.A(G244), .ZN(new_n231));
  OAI22_X1  g0031(.A1(new_n228), .A2(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G87), .ZN(new_n233));
  INV_X1    g0033(.A(G97), .ZN(new_n234));
  OAI22_X1  g0034(.A1(new_n233), .A2(new_n205), .B1(new_n234), .B2(new_n211), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n227), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT67), .B(G68), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G238), .ZN(new_n239));
  AOI21_X1  g0039(.A(new_n208), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(KEYINPUT1), .ZN(new_n241));
  OAI22_X1  g0041(.A1(new_n219), .A2(new_n223), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AOI211_X1 g0042(.A(new_n214), .B(new_n242), .C1(new_n241), .C2(new_n240), .ZN(G361));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT2), .B(G226), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G264), .B(G270), .Z(new_n248));
  XNOR2_X1  g0048(.A(G250), .B(G257), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G358));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G68), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G58), .B(G77), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n254), .B(new_n257), .Z(G351));
  AOI21_X1  g0058(.A(new_n221), .B1(new_n208), .B2(G33), .ZN(new_n259));
  XOR2_X1   g0059(.A(KEYINPUT8), .B(G58), .Z(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n260), .A2(new_n262), .B1(G150), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n209), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n228), .B1(new_n206), .B2(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n270), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n272), .A2(new_n273), .B1(new_n228), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n267), .A2(new_n268), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT9), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n261), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G222), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n283), .B1(new_n230), .B2(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n221), .B1(new_n261), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  AOI21_X1  g0091(.A(G1), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(G274), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n289), .A2(new_n292), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(G226), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G190), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n277), .B(new_n299), .C1(new_n300), .C2(new_n298), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n276), .B(new_n304), .C1(G179), .C2(new_n297), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n206), .A2(G20), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n260), .A2(new_n307), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n271), .A2(new_n308), .B1(new_n270), .B2(new_n260), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT67), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G68), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n314));
  OAI21_X1  g0114(.A(G58), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n207), .B1(new_n315), .B2(new_n202), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n207), .A2(new_n261), .ZN(new_n317));
  INV_X1    g0117(.A(G159), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT71), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n263), .A2(new_n320), .A3(G159), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT72), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n311), .A2(G68), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n225), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(G20), .B1(new_n326), .B2(new_n201), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT72), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n319), .A2(new_n321), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT69), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT69), .A2(G33), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT3), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT70), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT7), .ZN(new_n335));
  AOI21_X1  g0135(.A(G20), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n333), .A2(new_n279), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n338), .A2(G68), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n333), .A2(new_n279), .A3(new_n336), .ZN(new_n340));
  INV_X1    g0140(.A(new_n337), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n323), .A2(new_n330), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n259), .B1(new_n343), .B2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT69), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n261), .ZN(new_n346));
  NAND2_X1  g0146(.A1(KEYINPUT69), .A2(G33), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n278), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n279), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n348), .A2(new_n350), .B1(new_n352), .B2(new_n335), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT73), .B1(new_n353), .B2(new_n237), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n202), .B1(new_n237), .B2(new_n225), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(G20), .B1(new_n319), .B2(new_n321), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n331), .A2(new_n332), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n349), .B1(new_n358), .B2(new_n278), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n279), .B2(new_n351), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n357), .B(new_n238), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n354), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT74), .B1(new_n344), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n342), .A2(G68), .A3(new_n338), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n328), .B1(new_n327), .B2(new_n329), .ZN(new_n368));
  OAI211_X1 g0168(.A(KEYINPUT16), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n259), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n364), .A2(new_n369), .A3(KEYINPUT74), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n310), .B1(new_n365), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT76), .ZN(new_n374));
  INV_X1    g0174(.A(new_n292), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n288), .A2(new_n375), .A3(G232), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n293), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n229), .A2(new_n282), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n278), .B1(new_n346), .B2(new_n347), .ZN(new_n379));
  INV_X1    g0179(.A(new_n279), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n285), .A2(G1698), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  XOR2_X1   g0184(.A(new_n384), .B(KEYINPUT75), .Z(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n377), .B1(new_n386), .B2(new_n289), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n387), .A2(G179), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n303), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n374), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n387), .A2(new_n303), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n387), .A2(G179), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(KEYINPUT76), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n373), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT78), .B1(new_n387), .B2(G200), .ZN(new_n398));
  INV_X1    g0198(.A(G190), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n399), .A2(KEYINPUT77), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(KEYINPUT77), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n387), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n387), .A2(KEYINPUT78), .A3(new_n402), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n310), .B(new_n406), .C1(new_n365), .C2(new_n372), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n364), .A2(new_n369), .A3(new_n370), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT74), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n309), .B1(new_n412), .B2(new_n371), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT18), .B1(new_n413), .B2(new_n394), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(KEYINPUT17), .A3(new_n406), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n397), .A2(new_n409), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n238), .A2(new_n207), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n418), .A2(KEYINPUT12), .A3(new_n269), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT12), .B1(new_n274), .B2(new_n313), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n272), .A2(G68), .A3(new_n307), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT11), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n262), .A2(G77), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n228), .B2(new_n317), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n370), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n421), .B(new_n422), .C1(new_n423), .C2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n423), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n294), .B1(G238), .B2(new_n295), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n281), .A2(G232), .A3(G1698), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n281), .A2(G226), .A3(new_n282), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n289), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n432), .B1(new_n431), .B2(new_n437), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(new_n300), .ZN(new_n442));
  AOI211_X1 g0242(.A(new_n430), .B(new_n442), .C1(G190), .C2(new_n441), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT14), .B1(new_n441), .B2(new_n303), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n439), .A2(new_n440), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(G169), .ZN(new_n447));
  INV_X1    g0247(.A(G179), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n444), .B(new_n447), .C1(new_n448), .C2(new_n445), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n443), .B1(new_n449), .B2(new_n430), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n260), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n451));
  XOR2_X1   g0251(.A(KEYINPUT15), .B(G87), .Z(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n262), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n259), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n307), .A2(G77), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n271), .A2(new_n455), .B1(G77), .B2(new_n270), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n289), .A2(new_n292), .A3(new_n231), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n281), .A2(G232), .A3(new_n282), .ZN(new_n460));
  INV_X1    g0260(.A(G107), .ZN(new_n461));
  INV_X1    g0261(.A(G238), .ZN(new_n462));
  OAI221_X1 g0262(.A(new_n460), .B1(new_n461), .B2(new_n281), .C1(new_n284), .C2(new_n462), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n294), .B(new_n459), .C1(new_n463), .C2(new_n289), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n458), .B1(new_n464), .B2(G190), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n300), .B2(new_n464), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n448), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n467), .B(new_n458), .C1(G169), .C2(new_n464), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n306), .A2(new_n417), .A3(new_n450), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n206), .A2(G45), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n471), .A2(G274), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n205), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n288), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n333), .A2(new_n279), .ZN(new_n476));
  NOR2_X1   g0276(.A1(G238), .A2(G1698), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n231), .B2(G1698), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(G116), .B1(new_n331), .B2(new_n332), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n475), .B1(new_n481), .B2(new_n289), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n448), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n288), .B1(new_n479), .B2(new_n480), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n303), .B1(new_n485), .B2(new_n475), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(new_n482), .B2(new_n448), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT83), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n448), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT82), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(new_n486), .A4(new_n484), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n476), .A2(new_n207), .A3(G68), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT19), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n262), .A2(new_n495), .A3(G97), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G97), .A2(G107), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(new_n233), .B1(new_n435), .B2(new_n207), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n498), .B2(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n452), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n500), .A2(new_n370), .B1(new_n274), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n271), .B1(new_n206), .B2(G33), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n452), .B(KEYINPUT84), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n489), .A2(new_n493), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n482), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(G200), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT85), .B1(new_n482), .B2(G190), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n482), .A2(G190), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n512), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT86), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT86), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n508), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n270), .A2(G116), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n503), .B2(G116), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G283), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(new_n207), .C1(G33), .C2(new_n234), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n370), .B(new_n527), .C1(new_n207), .C2(G116), .ZN(new_n528));
  XNOR2_X1  g0328(.A(new_n528), .B(KEYINPUT20), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n206), .B(G45), .C1(new_n287), .C2(KEYINPUT5), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n534), .A2(G274), .A3(new_n288), .A4(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n535), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n532), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n289), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G270), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n379), .A2(new_n380), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n212), .A2(G1698), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(G257), .B2(G1698), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G303), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n281), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n289), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n531), .A2(KEYINPUT21), .A3(G169), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(G200), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n551), .B(new_n530), .C1(new_n402), .C2(new_n549), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  OAI21_X1  g0353(.A(G169), .B1(new_n525), .B2(new_n529), .ZN(new_n554));
  INV_X1    g0354(.A(new_n549), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n548), .A2(G179), .A3(new_n536), .A4(new_n540), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n530), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n550), .A2(new_n552), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n231), .A2(G1698), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT4), .B1(new_n476), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n281), .A2(G250), .A3(G1698), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n526), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n289), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n539), .A2(G257), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n536), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G190), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(G200), .ZN(new_n570));
  XNOR2_X1  g0370(.A(G97), .B(G107), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT79), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(KEYINPUT6), .ZN(new_n573));
  MUX2_X1   g0373(.A(new_n572), .B(G97), .S(KEYINPUT6), .Z(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT80), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT80), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n573), .B(new_n577), .C1(new_n571), .C2(new_n574), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n207), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n353), .A2(new_n461), .B1(new_n230), .B2(new_n317), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n370), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n270), .A2(G97), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n503), .B2(G97), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n569), .A2(new_n570), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n583), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n568), .A2(new_n448), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n567), .A2(new_n303), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n559), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n476), .A2(new_n207), .A3(G87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT22), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(KEYINPUT87), .A3(KEYINPUT22), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n281), .ZN(new_n598));
  NOR4_X1   g0398(.A1(new_n598), .A2(KEYINPUT22), .A3(G20), .A4(new_n233), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n461), .A2(G20), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT23), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n602), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(G20), .B2(new_n480), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n591), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n599), .B1(new_n595), .B2(new_n596), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n608), .A2(KEYINPUT24), .A3(new_n605), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n370), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT25), .B1(new_n274), .B2(new_n461), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n274), .A2(KEYINPUT25), .A3(new_n461), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n503), .A2(G107), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n211), .A2(G1698), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(G250), .B2(G1698), .ZN(new_n617));
  INV_X1    g0417(.A(G294), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n542), .A2(new_n617), .B1(new_n618), .B2(new_n358), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n289), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n539), .A2(G264), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n536), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(G179), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n303), .B2(new_n622), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n601), .A2(new_n591), .A3(new_n606), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT24), .B1(new_n608), .B2(new_n605), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n259), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n614), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n622), .A2(new_n399), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(G200), .B2(new_n622), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n590), .A2(new_n625), .A3(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n470), .A2(new_n522), .A3(new_n634), .ZN(G372));
  INV_X1    g0435(.A(new_n305), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n449), .A2(new_n430), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n443), .B2(new_n468), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n412), .A2(new_n371), .ZN(new_n639));
  AND4_X1   g0439(.A1(KEYINPUT17), .A2(new_n639), .A3(new_n310), .A4(new_n406), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT17), .B1(new_n413), .B2(new_n406), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n388), .A2(new_n389), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n639), .B2(new_n310), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n636), .B1(new_n647), .B2(new_n302), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n508), .A2(new_n520), .A3(new_n517), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n520), .B1(new_n508), .B2(new_n517), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n588), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n651), .A2(KEYINPUT91), .A3(KEYINPUT26), .A4(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n519), .A2(KEYINPUT26), .A3(new_n521), .A4(new_n652), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n507), .A2(new_n490), .A3(new_n486), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT88), .B1(new_n482), .B2(new_n300), .ZN(new_n657));
  OR3_X1    g0457(.A1(new_n482), .A2(KEYINPUT88), .A3(new_n300), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n657), .B(new_n658), .C1(new_n516), .C2(new_n513), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT89), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n510), .B(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n656), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n655), .B1(new_n662), .B2(new_n588), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT91), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n653), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n656), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n550), .A2(new_n556), .A3(new_n558), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n615), .B2(new_n624), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n669), .B(new_n624), .C1(new_n628), .C2(new_n629), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n668), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n662), .A2(new_n589), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(new_n633), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n667), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n666), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n648), .B1(new_n678), .B2(new_n470), .ZN(G369));
  NAND2_X1  g0479(.A1(new_n269), .A2(new_n207), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n668), .A2(new_n530), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n530), .A2(new_n686), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n559), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n625), .A2(new_n633), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n630), .B2(new_n686), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n615), .A2(new_n624), .A3(new_n685), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  OR3_X1    g0495(.A1(new_n670), .A2(new_n672), .A3(new_n685), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n668), .A2(new_n685), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(G399));
  NOR2_X1   g0499(.A1(new_n210), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n497), .A2(new_n233), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(G1), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n217), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(new_n701), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n651), .A2(new_n655), .A3(new_n652), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n656), .B(KEYINPUT95), .Z(new_n711));
  INV_X1    g0511(.A(new_n662), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n652), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n711), .B1(new_n713), .B2(KEYINPUT26), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n625), .A2(new_n668), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n633), .A3(new_n674), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n710), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n709), .B1(new_n717), .B2(new_n686), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n685), .B1(new_n666), .B2(new_n676), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n709), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT92), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n557), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n482), .A2(new_n621), .A3(new_n620), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n722), .A2(new_n723), .A3(new_n568), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n541), .A2(KEYINPUT92), .A3(G179), .A4(new_n548), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(KEYINPUT93), .A3(KEYINPUT30), .A4(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n722), .A2(new_n725), .A3(new_n723), .A4(new_n568), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n482), .A2(G179), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n567), .A2(new_n549), .A3(new_n622), .A4(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n736), .B2(new_n685), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n738), .B(new_n686), .C1(new_n731), .C2(new_n735), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT94), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n732), .A2(new_n734), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n730), .B2(new_n726), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n738), .B1(new_n742), .B2(new_n686), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT94), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n691), .A2(new_n651), .A3(new_n590), .A4(new_n686), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n740), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G330), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n720), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n708), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR2_X1   g0552(.A1(new_n209), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n206), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n700), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n210), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n281), .ZN(new_n758));
  INV_X1    g0558(.A(G355), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n758), .A2(new_n759), .B1(G116), .B2(new_n757), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n218), .A2(new_n291), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n476), .A2(new_n210), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G45), .B2(new_n257), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n220), .B1(G20), .B2(new_n303), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n756), .B1(new_n765), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n207), .A2(G179), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n598), .B1(new_n774), .B2(new_n546), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n773), .A2(new_n399), .A3(new_n300), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT99), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(KEYINPUT99), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n775), .B1(new_n780), .B2(G329), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n207), .A2(new_n448), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n402), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(G190), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G322), .A2(new_n784), .B1(new_n785), .B2(G311), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n773), .A2(new_n399), .A3(G200), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n781), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n207), .A2(new_n448), .A3(new_n300), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n791));
  INV_X1    g0591(.A(new_n402), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G326), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n399), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n207), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n794), .A2(new_n795), .B1(new_n618), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n789), .B1(KEYINPUT101), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n791), .A2(new_n399), .A3(new_n793), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT100), .Z(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT33), .B(G317), .Z(new_n802));
  OAI221_X1 g0602(.A(new_n799), .B1(KEYINPUT101), .B2(new_n798), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n801), .A2(new_n313), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n784), .B(KEYINPUT96), .Z(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n785), .B(KEYINPUT97), .Z(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G58), .A2(new_n806), .B1(new_n808), .B2(G77), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n788), .A2(new_n461), .ZN(new_n810));
  INV_X1    g0610(.A(new_n797), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(G97), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n812), .B(new_n281), .C1(new_n233), .C2(new_n774), .ZN(new_n813));
  INV_X1    g0613(.A(new_n794), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(G50), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n779), .A2(new_n318), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT32), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n809), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n803), .B1(new_n804), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n772), .B1(new_n819), .B2(new_n769), .ZN(new_n820));
  INV_X1    g0620(.A(new_n768), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n689), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n690), .A2(new_n756), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n689), .A2(G330), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(G396));
  OAI21_X1  g0625(.A(new_n466), .B1(new_n457), .B2(new_n686), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n468), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n468), .A2(new_n685), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n719), .B(new_n831), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(new_n749), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n756), .B1(new_n832), .B2(new_n749), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n769), .A2(new_n766), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n756), .B1(G77), .B2(new_n837), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n807), .A2(new_n702), .B1(new_n546), .B2(new_n794), .ZN(new_n839));
  INV_X1    g0639(.A(new_n784), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n618), .ZN(new_n841));
  INV_X1    g0641(.A(new_n788), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(G87), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n461), .B2(new_n774), .ZN(new_n844));
  INV_X1    g0644(.A(G311), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n598), .B1(new_n234), .B2(new_n797), .C1(new_n779), .C2(new_n845), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n839), .A2(new_n841), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n801), .B(KEYINPUT102), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n787), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n808), .A2(G159), .B1(G137), .B2(new_n814), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  INV_X1    g0651(.A(G143), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n850), .B1(new_n851), .B2(new_n801), .C1(new_n805), .C2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT34), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n476), .B1(new_n313), .B2(new_n788), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n797), .A2(new_n225), .B1(new_n774), .B2(new_n228), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(new_n780), .C2(G132), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n853), .B2(new_n854), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n849), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n838), .B1(new_n860), .B2(new_n769), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n767), .B2(new_n831), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT103), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n835), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  NAND2_X1  g0665(.A1(new_n576), .A2(new_n578), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n702), .B(new_n223), .C1(new_n866), .C2(KEYINPUT35), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(KEYINPUT35), .B2(new_n866), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  NAND3_X1  g0669(.A1(new_n217), .A2(G77), .A3(new_n315), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n313), .A2(G50), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT104), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n206), .B(G13), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n369), .A2(new_n370), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n310), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n683), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n396), .B1(new_n373), .B2(new_n395), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n413), .A2(KEYINPUT18), .A3(new_n394), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n880), .B1(new_n883), .B2(new_n642), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n373), .B1(new_n395), .B2(new_n879), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT37), .B1(new_n413), .B2(new_n406), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n644), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n878), .B1(new_n888), .B2(new_n879), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n407), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n875), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n880), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n416), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n887), .A2(new_n891), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(KEYINPUT105), .A3(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n416), .A2(new_n894), .B1(new_n887), .B2(new_n891), .ZN(new_n899));
  OR3_X1    g0699(.A1(new_n899), .A2(KEYINPUT105), .A3(KEYINPUT38), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT106), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n898), .A2(new_n900), .A3(KEYINPUT106), .A4(KEYINPUT39), .ZN(new_n904));
  INV_X1    g0704(.A(new_n887), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT107), .ZN(new_n906));
  AOI221_X4 g0706(.A(new_n309), .B1(new_n404), .B2(new_n405), .C1(new_n412), .C2(new_n371), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n906), .B1(new_n907), .B2(new_n645), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n373), .A2(new_n879), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n407), .B(KEYINPUT107), .C1(new_n413), .C2(new_n644), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n905), .B1(new_n911), .B2(KEYINPUT37), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n909), .B1(new_n646), .B2(new_n642), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n875), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT108), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n897), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n899), .A2(KEYINPUT108), .A3(KEYINPUT38), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n914), .A2(new_n915), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT109), .ZN(new_n920));
  AND4_X1   g0720(.A1(KEYINPUT108), .A2(new_n895), .A3(KEYINPUT38), .A4(new_n896), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT108), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT109), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n915), .A4(new_n914), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n903), .A2(new_n904), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n449), .A2(new_n430), .A3(new_n686), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n830), .B1(new_n719), .B2(new_n831), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n898), .A2(new_n900), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n430), .A2(new_n685), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n450), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n430), .B(new_n685), .C1(new_n443), .C2(new_n449), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n929), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n646), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n937), .B2(new_n683), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n928), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n648), .B1(new_n720), .B2(new_n470), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(G330), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n747), .A2(new_n743), .A3(new_n744), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT110), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(KEYINPUT40), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n943), .A2(new_n831), .A3(new_n934), .A4(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n943), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n934), .A2(new_n831), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n947), .B1(new_n950), .B2(new_n944), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n930), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT40), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n923), .A2(new_n914), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(new_n950), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n948), .A2(new_n470), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n942), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n957), .B2(new_n956), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n941), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n206), .B2(new_n753), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n941), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n874), .B1(new_n961), .B2(new_n962), .ZN(G367));
  NAND2_X1  g0763(.A1(new_n652), .A2(new_n685), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n585), .A2(new_n685), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n584), .A2(new_n588), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n696), .A2(new_n698), .A3(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT45), .Z(new_n969));
  AOI21_X1  g0769(.A(new_n967), .B1(new_n696), .B2(new_n698), .ZN(new_n970));
  XOR2_X1   g0770(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n969), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n695), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT112), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n698), .B1(new_n694), .B2(new_n697), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(new_n690), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n751), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n978), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT112), .B1(new_n980), .B2(new_n750), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n975), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT113), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n975), .A2(KEYINPUT113), .A3(new_n979), .A4(new_n981), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n750), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n700), .B(KEYINPUT41), .Z(new_n987));
  OAI21_X1  g0787(.A(new_n754), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n691), .A2(new_n697), .A3(new_n967), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(KEYINPUT42), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n588), .B1(new_n625), .B2(new_n966), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n989), .A2(KEYINPUT42), .B1(new_n686), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n661), .A2(new_n685), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n712), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n661), .A2(new_n667), .A3(new_n685), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n990), .A2(new_n992), .B1(KEYINPUT43), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n997), .B(new_n998), .Z(new_n999));
  INV_X1    g0799(.A(new_n967), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n695), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n999), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n988), .A2(new_n1002), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n770), .B1(new_n757), .B2(new_n501), .C1(new_n763), .C2(new_n250), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n756), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n811), .A2(G68), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n225), .B2(new_n774), .C1(new_n840), .C2(new_n851), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n281), .B1(new_n788), .B2(new_n230), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n814), .A2(G143), .B1(KEYINPUT114), .B2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(KEYINPUT114), .B2(new_n1008), .C1(new_n228), .C2(new_n807), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1007), .B(new_n1010), .C1(G137), .C2(new_n780), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n318), .B2(new_n848), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n848), .A2(new_n618), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n806), .A2(G303), .B1(G311), .B2(new_n814), .ZN(new_n1014));
  INV_X1    g0814(.A(G317), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n774), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(G116), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT46), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n779), .A2(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n842), .A2(G97), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n542), .C1(new_n461), .C2(new_n797), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n808), .B2(G283), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1014), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1012), .B1(new_n1013), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1005), .B1(new_n1027), .B2(new_n769), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n994), .A2(new_n768), .A3(new_n995), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1003), .A2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n981), .A2(new_n979), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n700), .C1(new_n751), .C2(new_n978), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1016), .A2(G77), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n785), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n313), .C1(new_n228), .C2(new_n840), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G159), .B2(new_n814), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n780), .A2(G150), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n505), .A2(new_n811), .ZN(new_n1039));
  AND4_X1   g0839(.A1(new_n476), .A2(new_n1038), .A3(new_n1021), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n260), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1037), .B(new_n1040), .C1(new_n1041), .C2(new_n801), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n805), .A2(new_n1015), .B1(new_n807), .B2(new_n546), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G322), .B2(new_n814), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n848), .B2(new_n845), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n797), .A2(new_n787), .B1(new_n774), .B2(new_n618), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n476), .B1(G116), .B2(new_n842), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n795), .C2(new_n779), .ZN(new_n1052));
  AOI21_X1  g0852(.A(KEYINPUT49), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT118), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(KEYINPUT118), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n769), .A3(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n758), .A2(new_n704), .B1(G107), .B2(new_n757), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n247), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT116), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n260), .A2(new_n228), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT50), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n704), .B(new_n291), .C1(new_n313), .C2(new_n230), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n762), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1059), .A2(G45), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1064), .A2(new_n1060), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1058), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n756), .B1(new_n1067), .B2(new_n771), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT117), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1057), .B(new_n1069), .C1(new_n694), .C2(new_n821), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1033), .B(new_n1070), .C1(new_n754), .C2(new_n980), .ZN(G393));
  NAND2_X1  g0871(.A1(new_n975), .A2(new_n755), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n770), .B1(new_n234), .B2(new_n757), .C1(new_n763), .C2(new_n254), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n756), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n848), .A2(new_n228), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n794), .A2(new_n851), .B1(new_n840), .B2(new_n318), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n811), .A2(G77), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1016), .A2(new_n238), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1078), .A2(new_n476), .A3(new_n843), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G143), .B2(new_n780), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1077), .B(new_n1081), .C1(new_n1041), .C2(new_n807), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n848), .A2(new_n546), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n794), .A2(new_n1015), .B1(new_n840), .B2(new_n845), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT52), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1035), .A2(new_n618), .B1(new_n774), .B2(new_n787), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G116), .B2(new_n811), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n281), .B(new_n810), .C1(new_n780), .C2(G322), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1075), .A2(new_n1082), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1074), .B1(new_n1090), .B2(new_n769), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n967), .B2(new_n821), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1072), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n984), .A2(new_n985), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n975), .B1(new_n981), .B2(new_n979), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1095), .A2(new_n701), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(G390));
  NAND2_X1  g0898(.A1(new_n903), .A2(new_n904), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n920), .A2(new_n925), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n927), .B1(new_n929), .B2(new_n935), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n717), .A2(new_n686), .A3(new_n827), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n829), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n934), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n954), .A3(new_n927), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n943), .A2(G330), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1108), .A2(new_n949), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n748), .A2(G330), .A3(new_n831), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1112), .A2(new_n935), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1102), .A2(new_n1106), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1111), .A2(new_n755), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n926), .A2(new_n766), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n756), .B1(new_n260), .B2(new_n837), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT120), .Z(new_n1118));
  INV_X1    g0918(.A(new_n769), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1078), .B1(new_n840), .B2(new_n702), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT121), .Z(new_n1121));
  AOI22_X1  g0921(.A1(new_n808), .A2(G97), .B1(G283), .B2(new_n814), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n598), .B1(new_n788), .B2(new_n313), .C1(new_n233), .C2(new_n774), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n780), .B2(G294), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n848), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(G107), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1128), .A2(KEYINPUT122), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(KEYINPUT122), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT53), .B1(new_n774), .B2(new_n851), .ZN(new_n1131));
  OR3_X1    g0931(.A1(new_n774), .A2(KEYINPUT53), .A3(new_n851), .ZN(new_n1132));
  INV_X1    g0932(.A(G125), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1132), .C1(new_n779), .C2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n797), .A2(new_n318), .B1(new_n788), .B2(new_n228), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n598), .B(new_n1135), .C1(G132), .C2(new_n784), .ZN(new_n1136));
  INV_X1    g0936(.A(G128), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n794), .C1(new_n807), .C2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1134), .B(new_n1139), .C1(new_n1126), .C2(G137), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1129), .A2(new_n1130), .A3(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1116), .B(new_n1118), .C1(new_n1119), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1115), .A2(new_n1142), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1108), .A2(new_n470), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1144), .B(new_n648), .C1(new_n720), .C2(new_n470), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1112), .A2(new_n935), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1109), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n929), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n943), .A2(G330), .A3(new_n831), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1104), .B1(new_n1150), .B2(new_n935), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1113), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1145), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1106), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n926), .B2(new_n1101), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1114), .B(new_n1153), .C1(new_n1155), .C2(new_n1109), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT119), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1111), .A2(KEYINPUT119), .A3(new_n1114), .A4(new_n1153), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1145), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n701), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1143), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(G378));
  NAND2_X1  g0967(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1168));
  OAI21_X1  g0968(.A(G330), .B1(new_n952), .B2(new_n955), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n276), .A2(new_n879), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n306), .B(new_n1170), .Z(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(G330), .C1(new_n952), .C2(new_n955), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(new_n939), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1175), .A2(new_n1176), .B1(new_n928), .B2(new_n938), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT57), .B1(new_n1168), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1145), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT57), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n700), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1174), .A2(new_n766), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n756), .B1(G50), .B2(new_n837), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n542), .A2(new_n287), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n779), .A2(new_n787), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n505), .C2(new_n785), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n788), .A2(new_n225), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n784), .B2(G107), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n1006), .A3(new_n1034), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G116), .B2(new_n814), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1190), .B(new_n1194), .C1(new_n234), .C2(new_n801), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT58), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G50), .B1(new_n261), .B2(new_n287), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1195), .A2(new_n1196), .B1(new_n1188), .B2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n785), .A2(G137), .B1(new_n811), .B2(G150), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n774), .B2(new_n1138), .C1(new_n840), .C2(new_n1137), .ZN(new_n1200));
  INV_X1    g1000(.A(G132), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n801), .A2(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G125), .C2(new_n814), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n780), .A2(G124), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n842), .C2(G159), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT59), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1206), .B(new_n1207), .C1(new_n1203), .C2(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1198), .B1(new_n1196), .B2(new_n1195), .C1(new_n1205), .C2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1187), .B1(new_n1210), .B2(new_n769), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1186), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n754), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1185), .A2(new_n1215), .ZN(G375));
  NAND2_X1  g1016(.A1(new_n935), .A2(new_n766), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n756), .B1(G68), .B2(new_n837), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n848), .A2(new_n1138), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n806), .A2(G137), .B1(G132), .B2(new_n814), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1035), .A2(new_n851), .B1(new_n797), .B2(new_n228), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G159), .B2(new_n1016), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n542), .B(new_n1191), .C1(new_n780), .C2(G128), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1220), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n848), .A2(new_n702), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n808), .A2(G107), .B1(G294), .B2(new_n814), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n840), .A2(new_n787), .B1(new_n234), .B2(new_n774), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n281), .B(new_n1227), .C1(G77), .C2(new_n842), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n780), .A2(G303), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1228), .A3(new_n1039), .A4(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1219), .A2(new_n1224), .B1(new_n1225), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1218), .B1(new_n1231), .B2(new_n769), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1162), .A2(new_n755), .B1(new_n1217), .B2(new_n1232), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1153), .A2(new_n987), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(G381));
  OR2_X1    g1036(.A1(G381), .A2(G384), .ZN(new_n1237));
  OR2_X1    g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(G387), .A2(new_n1237), .A3(G390), .A4(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1239), .A2(new_n1166), .A3(new_n1185), .A4(new_n1215), .ZN(G407));
  NAND2_X1  g1040(.A1(new_n684), .A2(G213), .ZN(new_n1241));
  OR3_X1    g1041(.A1(G375), .A2(G378), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(G407), .A3(G213), .ZN(G409));
  AND3_X1   g1043(.A1(new_n684), .A2(G213), .A3(G2897), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1235), .A2(KEYINPUT60), .A3(new_n1164), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n700), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1235), .B1(KEYINPUT60), .B2(new_n1164), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1233), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(new_n864), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n864), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1244), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1251), .A2(new_n1252), .A3(new_n1244), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G378), .B(new_n1215), .C1(new_n1181), .C2(new_n1184), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1182), .A2(new_n1213), .A3(new_n987), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1166), .B1(new_n1259), .B2(new_n1214), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1258), .A2(new_n1260), .B1(G213), .B2(new_n684), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1251), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT63), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G390), .B1(new_n1003), .B2(new_n1030), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  XOR2_X1   g1066(.A(G393), .B(G396), .Z(new_n1267));
  NAND3_X1  g1067(.A1(new_n1003), .A2(new_n1030), .A3(G390), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1267), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1030), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1271), .B(new_n1097), .C1(new_n988), .C2(new_n1002), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1270), .B1(new_n1265), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  NOR4_X1   g1074(.A1(new_n1262), .A2(new_n1264), .A3(new_n1274), .A4(KEYINPUT61), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1261), .A2(KEYINPUT63), .A3(new_n1263), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT124), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1276), .B(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n1282), .B(KEYINPUT62), .C1(new_n1261), .C2(new_n1263), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(new_n1241), .A3(new_n1263), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT126), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1284), .A2(KEYINPUT62), .A3(new_n1241), .A4(new_n1263), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT127), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1261), .A2(new_n1291), .A3(KEYINPUT62), .A4(new_n1263), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1281), .B1(new_n1288), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1274), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1279), .B1(new_n1294), .B2(new_n1295), .ZN(G405));
  NAND2_X1  g1096(.A1(G375), .A2(new_n1166), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1258), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(new_n1263), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(new_n1274), .ZN(G402));
endmodule


