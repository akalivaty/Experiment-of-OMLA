//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1196, new_n1197,
    new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT65), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n462), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n464), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n460), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n468), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n467), .A2(G136), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT66), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n461), .A2(new_n463), .A3(G2105), .A4(new_n464), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT67), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n480), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT68), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n461), .A2(new_n463), .A3(new_n490), .A4(new_n464), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT4), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n494));
  OR3_X1    g069(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  OAI22_X1  g070(.A1(new_n493), .A2(new_n494), .B1(new_n471), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OR3_X1    g072(.A1(new_n466), .A2(KEYINPUT70), .A3(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT70), .B1(new_n466), .B2(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n465), .A2(KEYINPUT69), .A3(G126), .A4(G2105), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n481), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT72), .A3(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n510), .A2(new_n512), .B1(KEYINPUT5), .B2(new_n509), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n509), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n517), .A2(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT73), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT7), .Z(new_n529));
  NAND3_X1  g104(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(G51), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n530), .B(new_n531), .C1(new_n523), .C2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n529), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n515), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n520), .A2(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n523), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n515), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n522), .A2(G543), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT74), .B(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n523), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT76), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  AND2_X1   g129(.A1(new_n513), .A2(new_n522), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G91), .ZN(new_n556));
  OAI211_X1 g131(.A(G53), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n558), .B2(KEYINPUT77), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(KEYINPUT77), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n515), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT78), .B1(new_n563), .B2(new_n515), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n520), .A2(G49), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n523), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n513), .ZN(new_n574));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n515), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT79), .Z(G288));
  AOI22_X1  g153(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  OR3_X1    g154(.A1(new_n579), .A2(KEYINPUT80), .A3(new_n515), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT80), .B1(new_n579), .B2(new_n515), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n555), .A2(G86), .B1(G48), .B2(new_n520), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n555), .A2(G85), .B1(G47), .B2(new_n520), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT81), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n515), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(G290));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NOR2_X1   g164(.A1(G301), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n574), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n513), .A2(G92), .A3(new_n522), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n590), .B1(new_n600), .B2(new_n589), .ZN(G284));
  AOI21_X1  g176(.A(new_n590), .B1(new_n600), .B2(new_n589), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  XOR2_X1   g180(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g187(.A(new_n471), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n475), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n615), .A2(new_n616), .B1(new_n617), .B2(G2100), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n616), .B2(new_n615), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n617), .A2(G2100), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n467), .A2(G135), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT85), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(G111), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(new_n481), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G123), .ZN(new_n628));
  AND2_X1   g203(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n629), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n621), .A2(new_n631), .A3(new_n633), .ZN(G156));
  INV_X1    g209(.A(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(G401));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT86), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n630), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(KEYINPUT87), .ZN(new_n666));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(KEYINPUT87), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n663), .A2(new_n664), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n668), .B2(new_n665), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(KEYINPUT88), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT89), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(G229));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G24), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n585), .A2(new_n587), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1986), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G25), .ZN(new_n693));
  INV_X1    g268(.A(G119), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n466), .A2(G107), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n696));
  OAI22_X1  g271(.A1(new_n481), .A2(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n467), .B2(G131), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n693), .B1(new_n698), .B2(new_n692), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  NOR2_X1   g277(.A1(new_n691), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(G6), .A2(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G305), .B2(new_n687), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n687), .A2(G22), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n687), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n705), .A2(new_n706), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n687), .A2(G23), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n577), .B2(new_n687), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT33), .B(G1976), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n707), .A2(new_n711), .A3(new_n712), .A4(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n703), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT92), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(KEYINPUT91), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT92), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n703), .A2(new_n725), .A3(new_n720), .A4(new_n718), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n724), .B1(new_n722), .B2(new_n726), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n692), .A2(G35), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G162), .B2(new_n692), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT29), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n736));
  OR3_X1    g311(.A1(new_n735), .A2(G2090), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT97), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(G2090), .B1(new_n735), .B2(new_n736), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n629), .A2(G29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  NAND2_X1  g317(.A1(G164), .A2(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G27), .B2(G29), .ZN(new_n744));
  INV_X1    g319(.A(G2078), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n687), .A2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G168), .B2(new_n687), .ZN(new_n748));
  INV_X1    g323(.A(G1966), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n742), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n687), .A2(G20), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT23), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n604), .B2(new_n687), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT98), .B(G1956), .Z(new_n755));
  OAI22_X1  g330(.A1(new_n754), .A2(new_n755), .B1(new_n745), .B2(new_n744), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G29), .A2(G32), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n467), .A2(G141), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT26), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n762), .A2(new_n763), .B1(G105), .B2(new_n475), .ZN(new_n764));
  INV_X1    g339(.A(G129), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n481), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n758), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n687), .A2(G19), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n547), .B2(new_n687), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G1341), .Z(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n777));
  OR2_X1    g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  NAND2_X1  g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(G29), .B1(new_n781), .B2(KEYINPUT24), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(KEYINPUT24), .B2(new_n781), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n477), .B2(new_n692), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n687), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n687), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1961), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n692), .A2(G26), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT28), .ZN(new_n792));
  OR2_X1    g367(.A1(G104), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n794));
  INV_X1    g369(.A(G128), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n481), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n467), .B2(G140), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n792), .B1(new_n797), .B2(new_n692), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2067), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n790), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n771), .A2(new_n774), .A3(new_n787), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n687), .A2(G4), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n600), .B2(new_n687), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1348), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT25), .Z(new_n806));
  INV_X1    g381(.A(new_n467), .ZN(new_n807));
  INV_X1    g382(.A(G139), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT93), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(KEYINPUT93), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n613), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(new_n466), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT94), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n810), .A2(new_n811), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  MUX2_X1   g392(.A(G33), .B(new_n817), .S(G29), .Z(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(G2072), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n818), .A2(G2072), .B1(new_n755), .B2(new_n754), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n757), .A2(new_n801), .A3(new_n804), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n739), .A2(new_n740), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n737), .A2(new_n738), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n730), .A2(new_n825), .ZN(G311));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n730), .A2(new_n827), .A3(new_n825), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n827), .B1(new_n730), .B2(new_n825), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(G150));
  NAND2_X1  g406(.A1(new_n600), .A2(G559), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT38), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n520), .A2(G55), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n523), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n513), .A2(G67), .ZN(new_n837));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n515), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n547), .A2(new_n840), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n542), .A2(new_n546), .B1(new_n836), .B2(new_n839), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n833), .B(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  INV_X1    g420(.A(G860), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n840), .A2(new_n846), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(G145));
  OR2_X1    g426(.A1(new_n817), .A2(new_n768), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n817), .A2(new_n767), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n797), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n506), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n852), .A2(new_n856), .A3(new_n853), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n698), .B(KEYINPUT100), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n615), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n467), .A2(G142), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n627), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n466), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n862), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n858), .A2(new_n868), .A3(new_n859), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(G162), .A2(new_n477), .ZN(new_n874));
  NAND2_X1  g449(.A1(G162), .A2(new_n477), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n629), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n632), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n876), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n880), .A2(new_n871), .A3(new_n870), .A4(new_n872), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(G395));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n840), .A2(G868), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n843), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n609), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  INV_X1    g466(.A(new_n566), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n558), .A2(KEYINPUT77), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n560), .A3(new_n556), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n892), .A2(new_n894), .A3(new_n598), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n562), .A2(new_n566), .B1(new_n597), .B2(new_n594), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(G299), .A2(new_n598), .ZN(new_n898));
  INV_X1    g473(.A(new_n598), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(new_n562), .A3(new_n566), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n900), .A3(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n890), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n895), .A2(new_n896), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(new_n890), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT42), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n585), .A2(new_n577), .A3(new_n587), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n577), .B1(new_n585), .B2(new_n587), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT103), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n907), .ZN(new_n913));
  XNOR2_X1  g488(.A(G305), .B(G166), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n914), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n916), .A2(new_n912), .A3(new_n911), .A4(new_n907), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n906), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n906), .A2(new_n919), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n886), .B(new_n888), .C1(new_n922), .C2(new_n589), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n589), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT104), .B1(new_n924), .B2(new_n887), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(G295));
  OAI21_X1  g501(.A(new_n888), .B1(new_n922), .B2(new_n589), .ZN(G331));
  AND3_X1   g502(.A1(new_n841), .A2(G301), .A3(new_n842), .ZN(new_n928));
  AOI21_X1  g503(.A(G301), .B1(new_n841), .B2(new_n842), .ZN(new_n929));
  OAI21_X1  g504(.A(G286), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n843), .A2(G171), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n841), .A2(G301), .A3(new_n842), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(G168), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n904), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n897), .A2(new_n901), .A3(new_n933), .A4(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT105), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n919), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n939), .B1(new_n935), .B2(new_n936), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n918), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n941), .A2(new_n944), .A3(new_n945), .A4(new_n882), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n918), .B2(new_n937), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(KEYINPUT44), .B(new_n946), .C1(new_n948), .C2(new_n945), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n941), .A2(new_n944), .A3(new_n882), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n941), .A2(new_n945), .A3(new_n947), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT106), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n956));
  AOI211_X1 g531(.A(new_n956), .B(KEYINPUT44), .C1(new_n951), .C2(new_n952), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n949), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n960), .B(new_n949), .C1(new_n955), .C2(new_n957), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(G397));
  XNOR2_X1  g537(.A(KEYINPUT108), .B(G1384), .ZN(new_n963));
  INV_X1    g538(.A(new_n500), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT69), .B1(new_n627), .B2(G126), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n481), .A2(new_n502), .A3(new_n503), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n495), .A2(new_n471), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT71), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT4), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT45), .B(new_n963), .C1(new_n967), .C2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G40), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n477), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n496), .B2(new_n505), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT56), .B(G2072), .Z(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n967), .B2(new_n972), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n977), .A2(KEYINPUT110), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n975), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT115), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT110), .B1(new_n506), .B2(new_n984), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n986), .B(G1384), .C1(new_n496), .C2(new_n505), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT50), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n975), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n991), .A2(new_n993), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1956), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n982), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n604), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(G299), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n566), .A2(new_n558), .A3(new_n556), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n1004), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT116), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1009), .A3(new_n1004), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1002), .A2(new_n1005), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT118), .B1(new_n1001), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n987), .A2(new_n988), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n990), .B1(new_n1015), .B2(KEYINPUT50), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n992), .B1(new_n1016), .B2(new_n997), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1956), .B1(new_n1017), .B2(new_n991), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1014), .B(new_n1011), .C1(new_n1018), .C2(new_n982), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n987), .A2(new_n983), .A3(new_n988), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT111), .B1(new_n977), .B2(new_n983), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n990), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n987), .A2(new_n988), .A3(KEYINPUT111), .A4(new_n983), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1348), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n987), .A2(new_n988), .A3(new_n975), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G2067), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n899), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1013), .A2(new_n1019), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n998), .A2(new_n993), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n997), .B1(new_n996), .B2(new_n975), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1000), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n982), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1012), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT119), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1028), .A2(new_n1036), .A3(new_n1033), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1001), .A2(new_n1012), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1031), .A2(new_n1012), .A3(new_n1032), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1996), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT58), .B(G1341), .Z(new_n1043));
  AOI22_X1  g618(.A1(new_n1042), .A2(new_n979), .B1(new_n1025), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n547), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(KEYINPUT120), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT59), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1025), .A2(new_n1043), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n976), .A2(new_n978), .A3(G1996), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(new_n1046), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(new_n975), .A3(new_n1023), .ZN(new_n1055));
  INV_X1    g630(.A(G1348), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1026), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n598), .A2(KEYINPUT60), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n598), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1027), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1061), .B1(KEYINPUT60), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1033), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1001), .A2(KEYINPUT122), .A3(new_n1012), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(KEYINPUT61), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1041), .B(new_n1064), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1035), .A2(new_n1037), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G305), .A2(G1981), .ZN(new_n1072));
  INV_X1    g647(.A(G1981), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n580), .A2(new_n1073), .A3(new_n581), .A4(new_n582), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(KEYINPUT49), .A3(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT113), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1025), .ZN(new_n1077));
  INV_X1    g652(.A(G8), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(KEYINPUT49), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1076), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT112), .B(G1976), .Z(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT52), .B1(G288), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  INV_X1    g660(.A(new_n577), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1079), .B(new_n1084), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1025), .B(G8), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1082), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G2090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1022), .A2(new_n1091), .A3(new_n1023), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n980), .A2(new_n710), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1078), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G166), .A2(new_n1078), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT55), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n979), .B2(new_n745), .ZN(new_n1099));
  INV_X1    g674(.A(G1961), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1055), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT45), .B1(new_n987), .B2(new_n988), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT45), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n975), .B1(new_n985), .B2(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n745), .A2(KEYINPUT53), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(G171), .B(KEYINPUT54), .Z(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT45), .B1(new_n506), .B2(new_n963), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n976), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(new_n1108), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1107), .A2(new_n1108), .B1(new_n1101), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1017), .A2(new_n1091), .A3(new_n991), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1078), .B1(new_n1113), .B2(new_n1093), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1097), .B(new_n1112), .C1(new_n1096), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1054), .A2(new_n785), .A3(new_n975), .A4(new_n1023), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n749), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1117), .B(G8), .C1(new_n1120), .C2(G286), .ZN(new_n1121));
  NOR2_X1   g696(.A1(G168), .A2(new_n1078), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g701(.A(KEYINPUT123), .B(new_n1123), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1121), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1117), .B(new_n1122), .C1(new_n1120), .C2(G8), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1116), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1124), .B(new_n1125), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1120), .A2(G8), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(KEYINPUT51), .A3(new_n1123), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1131), .A2(KEYINPUT124), .A3(new_n1133), .A4(new_n1121), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1115), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1071), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1130), .A2(new_n1134), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT62), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1130), .A2(new_n1134), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1097), .B1(new_n1096), .B2(new_n1114), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1107), .A2(G171), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1138), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(G288), .A2(G1976), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1082), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1074), .B(KEYINPUT114), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1079), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1149), .B2(new_n1090), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1120), .A2(G8), .A3(G168), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1141), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1151), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1097), .B(new_n1154), .C1(new_n1096), .C2(new_n1094), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1150), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1136), .A2(new_n1144), .A3(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1109), .A2(new_n975), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n797), .B(G2067), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n767), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1160), .B1(G1996), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n768), .A2(new_n1042), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n698), .B(new_n701), .Z(new_n1166));
  INV_X1    g741(.A(G1986), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1165), .B(new_n1166), .C1(new_n1167), .C2(new_n689), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n689), .A2(new_n1167), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT109), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1158), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1157), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT46), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n767), .B1(new_n1173), .B2(G1996), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1158), .B1(new_n1160), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1158), .A2(new_n1042), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1176), .A2(KEYINPUT126), .A3(new_n1173), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT126), .B1(new_n1176), .B2(new_n1173), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1175), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT47), .Z(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT48), .B1(new_n1170), .B2(new_n1158), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1170), .A2(KEYINPUT48), .A3(new_n1158), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1181), .B(new_n1182), .C1(new_n1158), .C2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n698), .A2(new_n701), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1164), .A2(new_n1185), .B1(G2067), .B2(new_n855), .ZN(new_n1186));
  AOI211_X1 g761(.A(new_n1180), .B(new_n1184), .C1(new_n1158), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1172), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g763(.A1(G401), .A2(new_n457), .A3(G227), .ZN(new_n1190));
  AND4_X1   g764(.A1(new_n684), .A2(new_n883), .A3(new_n685), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n1191), .A2(new_n1192), .A3(new_n953), .ZN(new_n1193));
  AOI21_X1  g767(.A(new_n1192), .B1(new_n1191), .B2(new_n953), .ZN(new_n1194));
  NOR2_X1   g768(.A1(new_n1193), .A2(new_n1194), .ZN(G308));
  NAND2_X1  g769(.A1(new_n1191), .A2(new_n953), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1196), .A2(KEYINPUT127), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n1191), .A2(new_n1192), .A3(new_n953), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n1198), .ZN(G225));
endmodule


