//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR3_X1   g0010(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G68), .A2(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n219), .B(new_n220), .C1(new_n202), .C2(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n218), .B(new_n222), .C1(G97), .C2(G257), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G1), .B2(G20), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n210), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n214), .B(new_n225), .C1(new_n227), .C2(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G257), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT65), .B(G250), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n236), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G238), .A2(G1698), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n256), .B(new_n257), .C1(new_n238), .C2(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n258), .B(new_n261), .C1(G107), .C2(new_n256), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT68), .ZN(new_n266));
  OAI21_X1  g0066(.A(G274), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n266), .B(new_n209), .C1(G41), .C2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n260), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G244), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n260), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n262), .B(new_n271), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT70), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT69), .B(G179), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n275), .B(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G20), .A2(G77), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n253), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT15), .B(G87), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n284), .B1(new_n285), .B2(new_n287), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n226), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n291), .A2(new_n293), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n293), .B1(new_n209), .B2(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G77), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT71), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT71), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n297), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n279), .A2(new_n283), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n288), .A2(G77), .B1(new_n286), .B2(G50), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(new_n210), .B2(G68), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n298), .A2(G68), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n295), .A2(G68), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT12), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT11), .B1(new_n308), .B2(new_n293), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT73), .B1(new_n267), .B2(new_n269), .ZN(new_n318));
  INV_X1    g0118(.A(G274), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n273), .B2(KEYINPUT68), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT73), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n260), .A4(new_n268), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n260), .A2(G238), .A3(new_n273), .ZN(new_n324));
  INV_X1    g0124(.A(G1698), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n221), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n238), .A2(G1698), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n326), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n260), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AND4_X1   g0133(.A1(new_n317), .A2(new_n323), .A3(new_n324), .A4(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n332), .B1(new_n318), .B2(new_n322), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n317), .B1(new_n335), .B2(new_n324), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n316), .B1(new_n337), .B2(G190), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n337), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n303), .B(new_n301), .C1(new_n276), .C2(new_n339), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n281), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n306), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G223), .A2(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n325), .A2(G222), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n256), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n261), .C1(G77), .C2(new_n256), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n271), .B(new_n350), .C1(new_n221), .C2(new_n274), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(new_n277), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n203), .A2(G20), .ZN(new_n353));
  INV_X1    g0153(.A(G150), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n353), .B1(new_n354), .B2(new_n287), .C1(new_n285), .C2(new_n289), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n293), .B1(new_n202), .B2(new_n296), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n298), .A2(G50), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n351), .A2(new_n282), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n351), .A2(new_n343), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT9), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n358), .A2(new_n363), .B1(G200), .B2(new_n351), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n356), .A2(KEYINPUT9), .A3(new_n357), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n365), .A2(KEYINPUT72), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(KEYINPUT72), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n362), .B(new_n364), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n368), .A2(KEYINPUT10), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(KEYINPUT10), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n361), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  INV_X1    g0172(.A(G68), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n254), .A2(new_n210), .A3(new_n255), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n255), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G58), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n373), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n380), .B2(new_n201), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n286), .A2(G159), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n372), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n328), .A2(new_n329), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT7), .B1(new_n385), .B2(new_n210), .ZN(new_n386));
  INV_X1    g0186(.A(new_n377), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n383), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n390), .A3(new_n293), .ZN(new_n391));
  INV_X1    g0191(.A(new_n285), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n295), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n298), .B2(new_n392), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n221), .A2(G1698), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n396), .B1(G223), .B2(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n260), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(new_n270), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n274), .A2(new_n238), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(G169), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n399), .A2(new_n270), .A3(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n278), .ZN(new_n406));
  AND4_X1   g0206(.A1(KEYINPUT18), .A2(new_n395), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n391), .B2(new_n394), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT18), .B1(new_n408), .B2(new_n406), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n395), .ZN(new_n411));
  INV_X1    g0211(.A(new_n399), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n412), .A2(new_n343), .A3(new_n271), .A4(new_n402), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n405), .B2(G200), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n411), .A2(KEYINPUT74), .A3(KEYINPUT17), .A4(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n414), .A2(new_n391), .A3(KEYINPUT74), .A4(new_n394), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT17), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n410), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(G169), .B1(new_n334), .B2(new_n336), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n337), .A2(G179), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n424), .B(G169), .C1(new_n334), .C2(new_n336), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n316), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n346), .A2(new_n371), .A3(new_n420), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT4), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(KEYINPUT78), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  OAI21_X1  g0233(.A(G244), .B1(new_n433), .B2(KEYINPUT4), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n431), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n272), .B1(KEYINPUT78), .B2(new_n429), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n256), .A2(new_n437), .A3(new_n325), .A4(new_n430), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G283), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n435), .A2(new_n436), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n261), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n264), .A2(G1), .ZN(new_n442));
  AND2_X1   g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  NOR2_X1   g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n445), .A2(new_n319), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n260), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G257), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n441), .A2(G190), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT79), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n440), .A2(new_n261), .B1(G257), .B2(new_n447), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT79), .A3(G190), .A4(new_n446), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n339), .B1(new_n452), .B2(new_n446), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n295), .A2(G97), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT76), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n456), .A2(new_n457), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n292), .A2(new_n226), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n209), .A2(G33), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT77), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n209), .A2(KEYINPUT77), .A3(G33), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n295), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n459), .B1(new_n467), .B2(G97), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n206), .B1(new_n376), .B2(new_n377), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n287), .A2(new_n294), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT6), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT75), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n207), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(G97), .A2(G107), .ZN(new_n476));
  NOR2_X1   g0276(.A1(G97), .A2(G107), .ZN(new_n477));
  OAI211_X1 g0277(.A(KEYINPUT75), .B(new_n471), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n210), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n469), .A2(new_n470), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n458), .B(new_n468), .C1(new_n480), .C2(new_n460), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n455), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n454), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n293), .B1(new_n462), .B2(new_n461), .ZN(new_n484));
  INV_X1    g0284(.A(new_n466), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n486), .A2(new_n205), .B1(new_n457), .B2(new_n456), .ZN(new_n487));
  OAI21_X1  g0287(.A(G107), .B1(new_n386), .B2(new_n387), .ZN(new_n488));
  INV_X1    g0288(.A(new_n479), .ZN(new_n489));
  INV_X1    g0289(.A(new_n470), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n487), .B1(new_n491), .B2(new_n293), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n441), .A2(new_n446), .A3(new_n448), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n492), .A2(new_n458), .B1(new_n493), .B2(new_n282), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n452), .A2(new_n278), .A3(new_n446), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n484), .A2(G116), .A3(new_n485), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n296), .A2(new_n216), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n216), .A2(G20), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n293), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n439), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT20), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n293), .A3(new_n499), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT20), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n497), .B(new_n498), .C1(new_n502), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n325), .A2(G257), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G264), .A2(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n256), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n509), .B(new_n261), .C1(G303), .C2(new_n256), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n445), .A2(G270), .A3(new_n260), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n446), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n506), .A2(new_n512), .A3(G169), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G179), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n506), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n506), .A2(new_n512), .A3(KEYINPUT21), .A4(G169), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n510), .A2(G190), .A3(new_n446), .A4(new_n511), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n503), .B(new_n504), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(new_n498), .A4(new_n497), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n446), .A2(new_n511), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n339), .B1(new_n524), .B2(new_n510), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT82), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n512), .A2(G200), .ZN(new_n527));
  INV_X1    g0327(.A(new_n506), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n521), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n483), .A2(new_n496), .A3(new_n520), .A4(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  INV_X1    g0333(.A(new_n290), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n467), .B2(new_n534), .ZN(new_n535));
  NOR4_X1   g0335(.A1(new_n464), .A2(KEYINPUT81), .A3(new_n466), .A4(new_n290), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n534), .A2(new_n295), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n210), .B(G68), .C1(new_n328), .C2(new_n329), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n331), .A2(new_n210), .ZN(new_n544));
  NOR4_X1   g0344(.A1(KEYINPUT80), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT80), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G87), .A2(G97), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n206), .ZN(new_n548));
  OAI211_X1 g0348(.A(KEYINPUT19), .B(new_n544), .C1(new_n545), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n538), .B1(new_n550), .B2(new_n293), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n537), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n272), .A2(G1698), .ZN(new_n553));
  OAI221_X1 g0353(.A(new_n553), .B1(G238), .B2(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n260), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n260), .B(G250), .C1(G1), .C2(new_n264), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n442), .A2(G274), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n278), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n552), .B(new_n561), .C1(G169), .C2(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n467), .A2(G87), .ZN(new_n563));
  INV_X1    g0363(.A(new_n538), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n539), .A2(new_n542), .ZN(new_n565));
  INV_X1    g0365(.A(new_n544), .ZN(new_n566));
  INV_X1    g0366(.A(G87), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n205), .A3(new_n206), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT80), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n547), .A2(new_n546), .A3(new_n206), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n565), .B1(new_n571), .B2(KEYINPUT19), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n563), .B(new_n564), .C1(new_n572), .C2(new_n460), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n560), .A2(G190), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(new_n575), .C1(new_n339), .C2(new_n560), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n562), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT24), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n210), .B(G87), .C1(new_n328), .C2(new_n329), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT22), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n256), .A2(new_n582), .A3(new_n210), .A4(G87), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n288), .A2(G116), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT23), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n586), .A2(new_n210), .A3(G107), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT23), .B1(new_n206), .B2(G20), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AND4_X1   g0390(.A1(new_n579), .A2(new_n584), .A3(new_n585), .A4(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n581), .B2(new_n583), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n579), .B1(new_n592), .B2(new_n585), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n293), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n295), .A2(G107), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT25), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n486), .A2(new_n206), .B1(KEYINPUT25), .B2(new_n596), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n594), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n256), .B1(G257), .B2(new_n325), .ZN(new_n601));
  NOR2_X1   g0401(.A1(G250), .A2(G1698), .ZN(new_n602));
  INV_X1    g0402(.A(G294), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n601), .A2(new_n602), .B1(new_n253), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n261), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n447), .A2(G264), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n446), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n282), .ZN(new_n608));
  INV_X1    g0408(.A(new_n607), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n516), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n600), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(G20), .B1(new_n254), .B2(new_n255), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n582), .B1(new_n612), .B2(G87), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n580), .A2(KEYINPUT22), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n585), .B(new_n590), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT24), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n592), .A2(new_n579), .A3(new_n585), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n598), .B1(new_n618), .B2(new_n293), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n609), .A2(G190), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n607), .A2(G200), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n597), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT83), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n611), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n611), .B2(new_n622), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n532), .B(new_n578), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n428), .A2(new_n626), .ZN(G372));
  INV_X1    g0427(.A(new_n428), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n557), .A2(KEYINPUT84), .A3(new_n558), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT84), .B1(new_n557), .B2(new_n558), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n554), .A2(new_n555), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n629), .A2(new_n630), .B1(new_n631), .B2(new_n260), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n282), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n552), .A2(new_n561), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT86), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n493), .A2(new_n282), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n636), .A2(new_n481), .A3(new_n495), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n578), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n635), .B1(new_n638), .B2(KEYINPUT26), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n621), .A2(new_n594), .A3(new_n597), .A4(new_n599), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n611), .A2(new_n520), .B1(new_n641), .B2(new_n620), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n640), .B(new_n483), .C1(new_n642), .C2(new_n637), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT85), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n573), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n551), .A2(KEYINPUT85), .A3(new_n563), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n632), .A2(G200), .B1(G190), .B2(new_n560), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n537), .A2(new_n551), .B1(new_n278), .B2(new_n560), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n647), .A2(new_n648), .B1(new_n649), .B2(new_n633), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n639), .B1(new_n643), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n628), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n407), .A2(new_n409), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n306), .A2(new_n340), .B1(new_n316), .B2(new_n426), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(new_n419), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n369), .A2(new_n370), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n361), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(G369));
  NOR2_X1   g0459(.A1(new_n624), .A2(new_n625), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n611), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n611), .A2(new_n520), .ZN(new_n662));
  INV_X1    g0462(.A(G13), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n209), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n661), .A2(new_n662), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n526), .B2(new_n530), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT87), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n506), .A2(new_n670), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n673), .B2(new_n676), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n611), .A2(new_n671), .ZN(new_n681));
  INV_X1    g0481(.A(new_n660), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n600), .A2(new_n670), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n672), .B1(new_n680), .B2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n211), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n686), .A2(KEYINPUT88), .A3(G41), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT88), .B1(new_n686), .B2(G41), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G1), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n569), .A2(new_n216), .A3(new_n570), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n690), .A2(new_n691), .B1(new_n229), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT91), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT85), .B1(new_n551), .B2(new_n563), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n460), .B1(new_n543), .B2(new_n549), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n464), .A2(new_n567), .A3(new_n466), .ZN(new_n697));
  NOR4_X1   g0497(.A1(new_n696), .A2(new_n644), .A3(new_n697), .A4(new_n538), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n648), .B1(new_n695), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(KEYINPUT26), .A3(new_n634), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n694), .B1(new_n700), .B2(new_n496), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n640), .B1(new_n577), .B2(new_n496), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n650), .A2(KEYINPUT91), .A3(KEYINPUT26), .A4(new_n637), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n635), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n482), .A2(new_n454), .B1(new_n494), .B2(new_n495), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n662), .A2(new_n706), .A3(new_n622), .A4(new_n650), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n671), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT92), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT92), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n711), .A3(new_n671), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n652), .A2(new_n714), .A3(new_n671), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n609), .A2(new_n517), .A3(new_n452), .A4(new_n560), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n493), .A2(new_n607), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n632), .A2(KEYINPUT89), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT89), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n722), .B1(new_n631), .B2(new_n260), .C1(new_n629), .C2(new_n630), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n277), .B1(new_n524), .B2(new_n510), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT90), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT90), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n721), .A2(new_n723), .A3(new_n727), .A4(new_n724), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n720), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n670), .B1(new_n719), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT31), .B(new_n670), .C1(new_n719), .C2(new_n729), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n732), .B(new_n733), .C1(new_n626), .C2(new_n670), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n716), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n693), .B1(new_n737), .B2(G1), .ZN(G364));
  AOI21_X1  g0538(.A(new_n690), .B1(G45), .B2(new_n664), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n678), .A2(new_n679), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n680), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n678), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n210), .A2(G190), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n277), .A2(new_n339), .A3(new_n747), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT95), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT95), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n277), .A2(G20), .A3(G190), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n339), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n751), .A2(G311), .B1(G326), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n210), .B1(new_n755), .B2(G190), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n754), .B1(new_n603), .B2(new_n756), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n747), .A2(new_n755), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G329), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n747), .A2(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G179), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT97), .ZN(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n210), .A2(new_n343), .A3(new_n339), .A4(G179), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G303), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n278), .A2(new_n762), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  XOR2_X1   g0571(.A(KEYINPUT33), .B(G317), .Z(new_n772));
  OAI221_X1 g0572(.A(new_n385), .B1(new_n768), .B2(new_n769), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n752), .A2(G200), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n774), .A2(KEYINPUT94), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(KEYINPUT94), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n766), .B(new_n773), .C1(new_n778), .C2(G322), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n758), .A2(new_n761), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n751), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n777), .A2(new_n379), .B1(new_n782), .B2(new_n294), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G50), .B2(new_n753), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT96), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n764), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G107), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n759), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n786), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n770), .A2(G68), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n767), .A2(G87), .ZN(new_n794));
  INV_X1    g0594(.A(new_n756), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G97), .ZN(new_n796));
  AND4_X1   g0596(.A1(new_n256), .A2(new_n793), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n784), .B2(new_n785), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n781), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n226), .B1(G20), .B2(new_n282), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n247), .A2(new_n264), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(KEYINPUT93), .B1(new_n264), .B2(new_n230), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n686), .A2(new_n256), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(KEYINPUT93), .C2(new_n801), .ZN(new_n804));
  NAND3_X1  g0604(.A1(G355), .A2(new_n256), .A3(new_n211), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(G116), .C2(new_n211), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n745), .A2(new_n800), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n799), .A2(new_n800), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n746), .A2(new_n739), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n742), .A2(new_n809), .ZN(G396));
  NAND2_X1  g0610(.A1(new_n652), .A2(new_n671), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n305), .A2(new_n670), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n304), .A2(new_n670), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n342), .B2(new_n344), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n305), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n811), .B(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(new_n735), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n740), .ZN(new_n821));
  XNOR2_X1  g0621(.A(KEYINPUT99), .B(G283), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n796), .B1(new_n206), .B2(new_n768), .C1(new_n771), .C2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  INV_X1    g0625(.A(new_n753), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n385), .B1(new_n825), .B2(new_n759), .C1(new_n826), .C2(new_n769), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n824), .B(new_n827), .C1(G116), .C2(new_n751), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n567), .B2(new_n764), .C1(new_n603), .C2(new_n777), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT100), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n764), .A2(new_n373), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n256), .B1(new_n756), .B2(new_n379), .C1(new_n768), .C2(new_n202), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n751), .A2(G159), .B1(G150), .B2(new_n770), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n753), .A2(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G143), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n777), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n831), .B(new_n832), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n837), .B2(new_n836), .C1(new_n839), .C2(new_n759), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n830), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n740), .B1(new_n841), .B2(new_n800), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n800), .A2(new_n743), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n842), .B1(G77), .B2(new_n844), .C1(new_n744), .C2(new_n818), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n821), .A2(new_n845), .ZN(G384));
  INV_X1    g0646(.A(new_n668), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n395), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n410), .B2(new_n419), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n411), .A2(new_n414), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n408), .A2(new_n406), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(new_n853), .A3(new_n848), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT37), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT103), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n856), .B(new_n849), .C1(new_n410), .C2(new_n419), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n851), .A2(KEYINPUT38), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n854), .B(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n415), .A2(new_n418), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n848), .B1(new_n654), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n851), .A2(new_n855), .A3(new_n857), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n859), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(KEYINPUT104), .A3(new_n858), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n851), .A2(new_n857), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT104), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT38), .A4(new_n855), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n866), .B1(new_n873), .B2(KEYINPUT39), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n426), .A2(KEYINPUT102), .A3(new_n316), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT102), .B1(new_n426), .B2(new_n316), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n670), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n410), .A2(new_n668), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n652), .A2(new_n818), .A3(new_n671), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n813), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n316), .A2(new_n670), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n340), .B(new_n884), .C1(new_n875), .C2(new_n876), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n426), .A2(new_n316), .A3(new_n670), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n873), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n880), .A2(new_n881), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n428), .B1(new_n713), .B2(new_n715), .ZN(new_n892));
  INV_X1    g0692(.A(new_n658), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n891), .B(new_n894), .Z(new_n895));
  NAND2_X1  g0695(.A1(new_n858), .A2(new_n864), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n817), .B1(new_n885), .B2(new_n886), .ZN(new_n897));
  AND4_X1   g0697(.A1(KEYINPUT40), .A2(new_n896), .A3(new_n734), .A4(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n734), .A2(new_n887), .A3(new_n818), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n869), .A2(new_n899), .A3(new_n872), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n628), .A2(new_n734), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n895), .A2(new_n905), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(KEYINPUT105), .B2(new_n907), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n908), .B1(KEYINPUT105), .B2(new_n907), .C1(new_n209), .C2(new_n664), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n475), .A2(new_n478), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n216), .B1(new_n910), .B2(KEYINPUT35), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n227), .C1(KEYINPUT35), .C2(new_n910), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT101), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT36), .ZN(new_n914));
  OAI21_X1  g0714(.A(G77), .B1(new_n379), .B2(new_n373), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n229), .A2(new_n915), .B1(G50), .B2(new_n373), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(G1), .A3(new_n663), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n909), .A2(new_n914), .A3(new_n917), .ZN(G367));
  NAND2_X1  g0718(.A1(new_n481), .A2(new_n670), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n706), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT106), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n496), .B2(new_n671), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n520), .A2(new_n670), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n682), .A3(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT42), .Z(new_n925));
  OAI21_X1  g0725(.A(new_n496), .B1(new_n921), .B2(new_n611), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n671), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n647), .A2(new_n671), .ZN(new_n929));
  MUX2_X1   g0729(.A(new_n650), .B(new_n635), .S(new_n929), .Z(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n928), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n928), .B2(new_n933), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT107), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n680), .A2(new_n684), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n922), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n934), .A2(new_n935), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n939), .B1(KEYINPUT107), .B2(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n936), .B(new_n938), .C1(new_n934), .C2(new_n935), .ZN(new_n942));
  INV_X1    g0742(.A(new_n921), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n672), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT44), .Z(new_n945));
  NAND2_X1  g0745(.A1(new_n922), .A2(new_n672), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT45), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n945), .A2(new_n947), .A3(new_n937), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n937), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n680), .B(new_n684), .ZN(new_n951));
  INV_X1    g0751(.A(new_n923), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n737), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n689), .B(KEYINPUT41), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n209), .B1(new_n664), .B2(G45), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n941), .B(new_n942), .C1(new_n957), .C2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n256), .B1(new_n771), .B2(new_n789), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n795), .A2(G68), .ZN(new_n962));
  INV_X1    g0762(.A(new_n763), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n962), .B1(new_n768), .B2(new_n379), .C1(new_n963), .C2(new_n294), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n961), .B(new_n964), .C1(G143), .C2(new_n753), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n778), .A2(G150), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n760), .A2(G137), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n751), .A2(G50), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n777), .A2(new_n769), .B1(new_n825), .B2(new_n826), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT108), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n759), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n256), .B1(new_n770), .B2(G294), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n763), .A2(G97), .B1(new_n795), .B2(G107), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n767), .A2(KEYINPUT46), .A3(G116), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n975), .B(new_n979), .C1(new_n751), .C2(new_n822), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n972), .A2(new_n973), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT46), .B1(new_n767), .B2(G116), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT109), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n969), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n740), .B1(new_n985), .B2(new_n800), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n235), .A2(new_n803), .B1(new_n686), .B2(new_n534), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n807), .ZN(new_n988));
  INV_X1    g0788(.A(new_n745), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n986), .B(new_n988), .C1(new_n989), .C2(new_n930), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n960), .A2(new_n990), .ZN(G387));
  XNOR2_X1  g0791(.A(new_n951), .B(new_n923), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n737), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n953), .A2(new_n736), .ZN(new_n994));
  INV_X1    g0794(.A(new_n689), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n751), .A2(G303), .B1(G311), .B2(new_n770), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n777), .B2(new_n974), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G322), .B2(new_n753), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT48), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n603), .B2(new_n768), .C1(new_n756), .C2(new_n823), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT49), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n760), .A2(G326), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n256), .B1(new_n763), .B2(G116), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n770), .A2(new_n392), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n795), .A2(new_n534), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n294), .B2(new_n768), .C1(new_n354), .C2(new_n759), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n256), .B1(new_n826), .B2(new_n789), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(G97), .C2(new_n787), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n202), .B2(new_n777), .C1(new_n373), .C2(new_n782), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1007), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n800), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n684), .A2(new_n745), .ZN(new_n1018));
  OR3_X1    g0818(.A1(new_n285), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1019));
  OAI21_X1  g0819(.A(KEYINPUT50), .B1(new_n285), .B2(G50), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n264), .A3(new_n1020), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n691), .B(new_n1021), .C1(G68), .C2(G77), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n803), .B1(new_n242), .B2(new_n264), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n691), .A2(new_n211), .A3(new_n256), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n211), .A2(G107), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n807), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1017), .A2(new_n1018), .A3(new_n1027), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n996), .B1(new_n958), .B2(new_n953), .C1(new_n740), .C2(new_n1028), .ZN(G393));
  INV_X1    g0829(.A(new_n803), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n807), .B1(new_n205), .B2(new_n211), .C1(new_n250), .C2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n764), .A2(new_n567), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n767), .A2(G68), .B1(new_n795), .B2(G77), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n256), .C1(new_n771), .C2(new_n202), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n285), .B2(new_n782), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT51), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n777), .A2(new_n789), .B1(new_n354), .B2(new_n826), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n1037), .B2(new_n1038), .C1(new_n835), .C2(new_n759), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n777), .A2(new_n825), .B1(new_n974), .B2(new_n826), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT52), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n782), .A2(new_n603), .B1(new_n216), .B2(new_n756), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n256), .B1(new_n760), .B2(G322), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n788), .B(new_n1044), .C1(new_n768), .C2(new_n823), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1043), .B1(new_n1045), .B2(KEYINPUT111), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1042), .B(new_n1046), .C1(KEYINPUT111), .C2(new_n1045), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n771), .A2(new_n769), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1040), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n740), .B1(new_n1049), .B2(new_n800), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1031), .B(new_n1050), .C1(new_n922), .C2(new_n989), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n950), .B2(new_n958), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n993), .A2(new_n950), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n689), .B1(new_n993), .B2(new_n950), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(G390));
  INV_X1    g0856(.A(KEYINPUT39), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n869), .B2(new_n872), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n743), .B1(new_n1058), .B2(new_n866), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n256), .B1(new_n963), .B2(new_n202), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G159), .B2(new_n795), .ZN(new_n1061));
  INV_X1    g0861(.A(G125), .ZN(new_n1062));
  INV_X1    g0862(.A(G128), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n759), .C1(new_n826), .C2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G132), .B2(new_n778), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT54), .B(G143), .Z(new_n1066));
  AOI22_X1  g0866(.A1(new_n751), .A2(new_n1066), .B1(G137), .B2(new_n770), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT115), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n767), .A2(G150), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT53), .Z(new_n1070));
  NAND3_X1  g0870(.A1(new_n1065), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n385), .B1(new_n603), .B2(new_n759), .C1(new_n826), .C2(new_n765), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n794), .B1(new_n294), .B2(new_n756), .C1(new_n771), .C2(new_n206), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1072), .A2(new_n831), .A3(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n205), .B2(new_n782), .C1(new_n216), .C2(new_n777), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1076), .A2(new_n800), .B1(new_n285), .B2(new_n843), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1059), .A2(new_n739), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n887), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n735), .B2(new_n817), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n734), .A2(new_n887), .A3(G330), .A4(new_n818), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n710), .A2(new_n712), .A3(new_n813), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1084), .A2(KEYINPUT112), .A3(new_n816), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT112), .B1(new_n1084), .B2(new_n816), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1080), .A2(new_n1081), .B1(new_n813), .B2(new_n882), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n903), .A2(new_n679), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n892), .A2(new_n1092), .A3(new_n893), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT113), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT112), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n708), .A2(new_n711), .A3(new_n671), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n711), .B1(new_n708), .B2(new_n671), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n812), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n816), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1082), .B1(new_n1100), .B2(new_n1085), .ZN(new_n1101));
  OAI211_X1 g0901(.A(KEYINPUT113), .B(new_n1093), .C1(new_n1101), .C2(new_n1089), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1094), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT114), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n995), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1100), .A2(new_n887), .A3(new_n1085), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n865), .A2(new_n879), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n888), .B1(new_n670), .B2(new_n878), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n866), .B2(new_n1058), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1109), .A2(new_n1111), .A3(new_n1081), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1081), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1106), .A2(new_n958), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1114), .B1(new_n1117), .B2(new_n995), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1078), .B1(new_n1116), .B2(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(KEYINPUT57), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1093), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT113), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1100), .A2(new_n1085), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1089), .B1(new_n1123), .B2(new_n1083), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(new_n1124), .B2(new_n1121), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1102), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1121), .B1(new_n1114), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n900), .A2(new_n901), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n898), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n358), .A2(new_n847), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT56), .Z(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT55), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n371), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n371), .A2(new_n1133), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1132), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1136), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n1134), .A3(new_n1131), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1137), .A2(new_n1139), .A3(KEYINPUT120), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AND4_X1   g0941(.A1(G330), .A2(new_n1128), .A3(new_n1129), .A4(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT120), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n902), .B2(G330), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n891), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1128), .A2(G330), .A3(new_n1129), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n889), .B1(new_n874), .B2(new_n879), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n902), .A2(G330), .A3(new_n1141), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1149), .A2(new_n881), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1146), .A2(new_n1152), .A3(KEYINPUT121), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT121), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n891), .B(new_n1154), .C1(new_n1142), .C2(new_n1145), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1120), .B1(new_n1127), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT123), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1081), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1109), .A2(new_n1111), .A3(new_n1081), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n1094), .C2(new_n1103), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1164), .A2(new_n1093), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n689), .B1(new_n1165), .B2(KEYINPUT57), .ZN(new_n1166));
  OAI211_X1 g0966(.A(KEYINPUT123), .B(new_n1120), .C1(new_n1127), .C2(new_n1156), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1159), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1153), .A2(new_n959), .A3(new_n1155), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT122), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n202), .B1(new_n328), .B2(G41), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n777), .A2(new_n206), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT116), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n963), .A2(new_n379), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G77), .B2(new_n767), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n962), .C1(new_n205), .C2(new_n771), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n534), .B2(new_n751), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n385), .B1(new_n759), .B2(new_n765), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G41), .B(new_n1178), .C1(new_n753), .C2(G116), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1173), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1171), .B1(new_n1181), .B2(KEYINPUT58), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT117), .Z(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n770), .A2(G132), .B1(new_n767), .B2(new_n1066), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n826), .B2(new_n1062), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G137), .B2(new_n751), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n1063), .B2(new_n777), .C1(new_n354), .C2(new_n756), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT118), .Z(new_n1189));
  INV_X1    g0989(.A(KEYINPUT59), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G33), .B1(new_n760), .B2(G124), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G41), .B1(new_n763), .B2(G159), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1183), .A2(new_n1184), .A3(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT119), .Z(new_n1197));
  AOI21_X1  g0997(.A(new_n740), .B1(new_n1197), .B2(new_n800), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1137), .A2(new_n743), .A3(new_n1139), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(G50), .C2(new_n844), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1169), .A2(new_n1170), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1170), .B1(new_n1169), .B2(new_n1200), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1168), .A2(new_n1203), .ZN(G375));
  NAND2_X1  g1004(.A1(new_n1124), .A2(new_n1121), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1125), .A2(new_n1102), .A3(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1206), .A2(new_n955), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT124), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n777), .A2(new_n765), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n751), .A2(G107), .B1(G116), .B2(new_n770), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT125), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n385), .B1(new_n769), .B2(new_n759), .C1(new_n826), .C2(new_n603), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1009), .B1(new_n205), .B2(new_n768), .C1(new_n764), .C2(new_n294), .ZN(new_n1213));
  OR4_X1    g1013(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT126), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n778), .A2(G137), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n770), .A2(new_n1066), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n751), .A2(G150), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n826), .A2(new_n839), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n768), .A2(new_n789), .B1(new_n756), .B2(new_n202), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n256), .B1(new_n759), .B2(new_n1063), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(new_n1219), .A2(new_n1174), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1215), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n740), .B1(new_n1224), .B2(new_n800), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(G68), .B2(new_n844), .C1(new_n744), .C2(new_n887), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1124), .B2(new_n958), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1208), .A2(new_n1228), .ZN(G381));
  NOR2_X1   g1029(.A1(G375), .A2(G378), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(G381), .A2(G384), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n941), .A2(new_n942), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n959), .B1(new_n954), .B2(new_n956), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n990), .B(new_n1055), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1234), .A2(G396), .A3(G393), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1230), .A2(new_n1231), .A3(new_n1235), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n669), .A2(G213), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT127), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1230), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G407), .A2(G213), .A3(new_n1240), .ZN(G409));
  XOR2_X1   g1041(.A(G393), .B(G396), .Z(new_n1242));
  AOI21_X1  g1042(.A(new_n1055), .B1(new_n960), .B2(new_n990), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1234), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1243), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(G393), .B(G396), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1234), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1168), .A2(G378), .A3(new_n1203), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1078), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1118), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1115), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1127), .A2(new_n1156), .A3(new_n955), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1200), .B1(new_n1255), .B2(new_n958), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1253), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1250), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT60), .B1(new_n1124), .B2(new_n1121), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1206), .B2(KEYINPUT60), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n995), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1228), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n845), .A3(new_n821), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(G384), .A3(new_n1228), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1258), .A2(new_n1237), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1239), .B1(new_n1250), .B2(new_n1257), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1267), .A2(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n669), .A2(G213), .A3(G2897), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1266), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1238), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(G2897), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1272), .B1(new_n1277), .B2(new_n1269), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1249), .B1(new_n1271), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1265), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1249), .B1(new_n1269), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1258), .A2(new_n1237), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1266), .A2(new_n1273), .B1(new_n1275), .B2(G2897), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1280), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1267), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1282), .B(new_n1272), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1279), .A2(new_n1287), .ZN(G405));
  NAND2_X1  g1088(.A1(G375), .A2(new_n1253), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1249), .A2(new_n1250), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1250), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(new_n1245), .A3(new_n1248), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1265), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1290), .A2(new_n1292), .A3(new_n1266), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(G402));
endmodule


