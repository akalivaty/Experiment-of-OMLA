//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n470), .C1(new_n464), .C2(new_n465), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n471), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n472), .B1(new_n471), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n469), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n466), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n466), .A2(new_n470), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n464), .B2(new_n465), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n465), .C2(new_n464), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  NOR2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT68), .B(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n511), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g093(.A(KEYINPUT68), .B(G651), .Z(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n508), .A2(new_n514), .A3(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND2_X1  g097(.A1(new_n513), .A2(G89), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT69), .B(G51), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n507), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n511), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n523), .A2(new_n525), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n513), .A2(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n507), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n503), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n503), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n505), .A2(G81), .A3(new_n511), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n505), .A2(G43), .A3(G543), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND3_X1  g124(.A1(new_n505), .A2(G53), .A3(G543), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT9), .ZN(new_n551));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT70), .Z(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n554), .B2(new_n516), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n513), .A2(G91), .B1(new_n555), .B2(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n551), .A2(new_n556), .ZN(G299));
  OAI21_X1  g132(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n558));
  INV_X1    g133(.A(G49), .ZN(new_n559));
  INV_X1    g134(.A(G87), .ZN(new_n560));
  OAI221_X1 g135(.A(new_n558), .B1(new_n506), .B2(new_n559), .C1(new_n560), .C2(new_n512), .ZN(G288));
  INV_X1    g136(.A(G61), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n509), .B2(new_n510), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT71), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G73), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n566), .B1(new_n563), .B2(KEYINPUT71), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n519), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT72), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n570), .B(new_n519), .C1(new_n565), .C2(new_n567), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n505), .A2(G86), .A3(new_n511), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g149(.A1(G48), .A2(G543), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n572), .A2(new_n573), .B1(new_n505), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n569), .A2(new_n571), .A3(new_n574), .A4(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(new_n507), .A2(G47), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  XOR2_X1   g154(.A(KEYINPUT74), .B(G85), .Z(new_n580));
  OAI221_X1 g155(.A(new_n578), .B1(new_n503), .B2(new_n579), .C1(new_n512), .C2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  INV_X1    g157(.A(G92), .ZN(new_n583));
  XNOR2_X1  g158(.A(KEYINPUT75), .B(KEYINPUT10), .ZN(new_n584));
  OR3_X1    g159(.A1(new_n512), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n512), .B2(new_n583), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G651), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n507), .A2(G54), .ZN(new_n590));
  AND4_X1   g165(.A1(new_n585), .A2(new_n586), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n582), .B1(new_n591), .B2(G868), .ZN(G284));
  OAI21_X1  g167(.A(new_n582), .B1(new_n591), .B2(G868), .ZN(G321));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G286), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g170(.A(G299), .B(KEYINPUT76), .Z(new_n596));
  AOI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n594), .ZN(G297));
  AOI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n594), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n591), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n482), .A2(G123), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT79), .Z(new_n606));
  OAI21_X1  g181(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n607));
  INV_X1    g182(.A(G111), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G2105), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n480), .B2(G135), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G2096), .ZN(new_n613));
  INV_X1    g188(.A(G2096), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT3), .B(G2104), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n474), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT78), .B(G2100), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n611), .A2(new_n614), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n613), .B(new_n621), .C1(new_n620), .C2(new_n619), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2430), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n631), .A2(new_n632), .ZN(new_n637));
  AOI21_X1  g212(.A(KEYINPUT83), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(KEYINPUT83), .A3(new_n637), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n629), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n640), .ZN(new_n642));
  NOR3_X1   g217(.A1(new_n642), .A2(new_n638), .A3(new_n628), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n627), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n628), .B1(new_n642), .B2(new_n638), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n639), .A2(new_n640), .A3(new_n629), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(new_n626), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n644), .A2(new_n649), .A3(new_n647), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2100), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT19), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n669), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(KEYINPUT84), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1981), .B(G1986), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT85), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n681), .B(new_n685), .ZN(G229));
  NAND2_X1  g261(.A1(new_n480), .A2(G139), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT25), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(KEYINPUT90), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n615), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n695));
  OAI22_X1  g270(.A1(new_n691), .A2(new_n694), .B1(new_n470), .B2(new_n695), .ZN(new_n696));
  MUX2_X1   g271(.A(G33), .B(new_n696), .S(G29), .Z(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT91), .Z(new_n698));
  INV_X1    g273(.A(G2072), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G35), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G162), .B2(new_n701), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT29), .Z(new_n704));
  INV_X1    g279(.A(G2090), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT94), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n698), .A2(new_n699), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G20), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT23), .Z(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G299), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1956), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n700), .A2(new_n707), .A3(new_n708), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n701), .A2(G26), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n482), .A2(G128), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT89), .Z(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n719));
  INV_X1    g294(.A(G116), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G2105), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n480), .B2(G140), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2067), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G27), .A2(G29), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G164), .B2(G29), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G2078), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n612), .A2(new_n701), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT31), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(G11), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(G28), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n701), .B1(new_n734), .B2(G28), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n732), .B(new_n733), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NOR4_X1   g312(.A1(new_n726), .A2(new_n729), .A3(new_n730), .A4(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G29), .B2(G32), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n480), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n482), .A2(G129), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT26), .Z(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(new_n701), .ZN(new_n746));
  MUX2_X1   g321(.A(new_n740), .B(new_n739), .S(new_n746), .Z(new_n747));
  XOR2_X1   g322(.A(KEYINPUT27), .B(G1996), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT24), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G34), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n701), .B1(new_n750), .B2(G34), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n753), .B2(new_n752), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G160), .B2(G29), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G2084), .ZN(new_n757));
  NOR2_X1   g332(.A1(G4), .A2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n591), .B2(G16), .ZN(new_n759));
  INV_X1    g334(.A(G1348), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n738), .A2(new_n749), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n709), .A2(G5), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G171), .B2(new_n709), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(G1961), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n705), .B2(new_n704), .ZN(new_n766));
  NAND2_X1  g341(.A1(G286), .A2(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n709), .A2(G21), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G19), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n544), .B2(G16), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n770), .A2(G1966), .B1(G1341), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(G1341), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G2084), .B2(new_n756), .ZN(new_n775));
  INV_X1    g350(.A(G1966), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n769), .A2(new_n776), .B1(new_n764), .B2(G1961), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n766), .A2(new_n773), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n714), .A2(new_n762), .A3(new_n778), .ZN(new_n779));
  MUX2_X1   g354(.A(G6), .B(G305), .S(G16), .Z(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT32), .B(G1981), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n709), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n709), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT87), .B(G1971), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n780), .A2(new_n781), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n709), .A2(G23), .ZN(new_n788));
  INV_X1    g363(.A(G288), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n709), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT33), .B(G1976), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AND4_X1   g367(.A1(new_n782), .A2(new_n786), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT86), .B(KEYINPUT34), .Z(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  MUX2_X1   g371(.A(G24), .B(G290), .S(G16), .Z(new_n797));
  AND2_X1   g372(.A1(new_n797), .A2(G1986), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(G1986), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n480), .A2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n482), .A2(G119), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n470), .A2(G107), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n800), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G25), .B(new_n804), .S(G29), .Z(new_n805));
  XOR2_X1   g380(.A(KEYINPUT35), .B(G1991), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n798), .A2(new_n799), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n795), .A2(new_n796), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n812), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n795), .A2(new_n814), .A3(new_n796), .A4(new_n810), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n779), .A2(new_n813), .A3(new_n815), .ZN(G150));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n817));
  XNOR2_X1  g392(.A(G150), .B(new_n817), .ZN(G311));
  NAND4_X1  g393(.A1(new_n585), .A2(new_n586), .A3(new_n589), .A4(new_n590), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n599), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n511), .A2(G67), .ZN(new_n822));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n822), .A2(KEYINPUT96), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n519), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT96), .B1(new_n822), .B2(new_n823), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n505), .A2(G55), .A3(G543), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n505), .A2(G93), .A3(new_n511), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(new_n544), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n828), .B(new_n829), .C1(new_n825), .C2(new_n826), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(new_n543), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n821), .B(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n837), .A2(new_n838), .A3(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n833), .A2(G860), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT97), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  OR2_X1    g417(.A1(new_n839), .A2(new_n842), .ZN(G145));
  INV_X1    g418(.A(new_n499), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n498), .B1(new_n615), .B2(new_n495), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n488), .B(new_n492), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n723), .B(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(G130), .A2(new_n482), .B1(new_n480), .B2(G142), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  INV_X1    g424(.A(G118), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n849), .A2(KEYINPUT98), .B1(new_n850), .B2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(KEYINPUT98), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n847), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT99), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n804), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n618), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n696), .B(new_n745), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n478), .B(new_n486), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n611), .B(new_n864), .Z(new_n865));
  NAND3_X1  g440(.A1(new_n854), .A2(new_n860), .A3(new_n861), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n863), .A2(new_n866), .ZN(new_n870));
  INV_X1    g445(.A(new_n865), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g449(.A1(new_n833), .A2(new_n594), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n835), .B(new_n601), .ZN(new_n876));
  XNOR2_X1  g451(.A(G299), .B(new_n819), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT100), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n591), .A2(G299), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n819), .A2(new_n551), .A3(new_n556), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(KEYINPUT101), .A3(new_n882), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n591), .A2(G299), .A3(KEYINPUT101), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n877), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n876), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(G290), .B(G305), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n789), .B(G303), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT42), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n890), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n875), .B1(new_n897), .B2(new_n594), .ZN(G295));
  OAI21_X1  g473(.A(new_n875), .B1(new_n897), .B2(new_n594), .ZN(G331));
  AOI21_X1  g474(.A(new_n885), .B1(new_n883), .B2(new_n884), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n835), .A2(G171), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n832), .A2(new_n834), .A3(G301), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(G168), .A3(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n832), .A2(G301), .A3(new_n834), .ZN(new_n904));
  AOI21_X1  g479(.A(G301), .B1(new_n832), .B2(new_n834), .ZN(new_n905));
  OAI21_X1  g480(.A(G286), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n906), .A2(new_n903), .A3(new_n887), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n907), .B1(new_n908), .B2(new_n877), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n909), .B2(new_n893), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n904), .A2(new_n905), .A3(G286), .ZN(new_n912));
  AOI21_X1  g487(.A(G168), .B1(new_n901), .B2(new_n902), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n877), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n886), .A2(new_n906), .A3(new_n903), .A4(new_n888), .ZN(new_n915));
  AOI211_X1 g490(.A(KEYINPUT104), .B(new_n893), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n915), .ZN(new_n918));
  INV_X1    g493(.A(new_n893), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n910), .B(new_n911), .C1(new_n916), .C2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n914), .A2(new_n915), .A3(new_n893), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n868), .B(new_n924), .C1(new_n916), .C2(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n918), .A2(new_n919), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT104), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n918), .A2(new_n917), .A3(new_n919), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(KEYINPUT105), .A3(new_n911), .A4(new_n910), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n923), .A2(new_n926), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n925), .A2(new_n911), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n930), .A2(KEYINPUT43), .A3(new_n910), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(G397));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(G164), .B2(G1384), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n469), .B(G40), .C1(new_n476), .C2(new_n477), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n723), .A2(G2067), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n725), .A3(new_n722), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1996), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n745), .B(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n806), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n804), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n804), .A2(new_n949), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n946), .A2(new_n948), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(G290), .B(G1986), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n943), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1961), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(G164), .B2(G1384), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n844), .A2(new_n845), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT107), .B(new_n959), .C1(new_n960), .C2(new_n493), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n846), .A2(new_n959), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(KEYINPUT50), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n957), .A2(new_n961), .A3(new_n963), .A4(new_n958), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n942), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT118), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT118), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n971), .B(new_n942), .C1(new_n966), .C2(new_n967), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n955), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n957), .B2(new_n961), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n846), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  OR4_X1    g552(.A1(new_n974), .A2(new_n975), .A3(new_n977), .A4(G2078), .ZN(new_n978));
  INV_X1    g553(.A(G2078), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n969), .A2(new_n941), .A3(new_n976), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n974), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT125), .Z(new_n982));
  NAND3_X1  g557(.A1(new_n973), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(G171), .ZN(new_n984));
  INV_X1    g559(.A(new_n941), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n985), .A2(new_n974), .A3(G2078), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n986), .A2(new_n976), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n973), .A2(G301), .A3(new_n982), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT54), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n973), .A2(new_n982), .A3(new_n989), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n994), .B2(G171), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(G171), .B2(new_n983), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n969), .A2(new_n957), .A3(new_n961), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n997), .A2(G8), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n789), .A2(G1976), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT109), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n789), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(G8), .A3(new_n997), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1001), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n505), .A2(new_n575), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n568), .A2(new_n572), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G1981), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT49), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1009), .B(new_n1012), .C1(G305), .C2(G1981), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1013), .A2(new_n998), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1009), .B1(G305), .B2(G1981), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1002), .A2(new_n1006), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G303), .A2(G8), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n1018), .B(KEYINPUT55), .Z(new_n1019));
  AOI211_X1 g594(.A(G2090), .B(new_n942), .C1(new_n966), .C2(new_n967), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n977), .A2(new_n985), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT106), .B(G1971), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1019), .B(G8), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n957), .A2(new_n961), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1026), .B(new_n969), .C1(new_n1027), .C2(new_n958), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n958), .B1(new_n957), .B2(new_n961), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT111), .B1(new_n1029), .B2(new_n942), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G164), .A2(G1384), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n958), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1028), .A2(new_n705), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1023), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1025), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1017), .B(new_n1024), .C1(new_n1019), .C2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n776), .B1(new_n975), .B2(new_n977), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT112), .B(new_n776), .C1(new_n975), .C2(new_n977), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n942), .B1(new_n966), .B2(new_n967), .ZN(new_n1041));
  INV_X1    g616(.A(G2084), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1039), .A2(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G286), .A2(G8), .ZN(new_n1044));
  XOR2_X1   g619(.A(new_n1044), .B(KEYINPUT123), .Z(new_n1045));
  NOR2_X1   g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1043), .B2(new_n1025), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT124), .B(KEYINPUT51), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT51), .B(new_n1045), .C1(new_n1043), .C2(new_n1025), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1036), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n993), .A2(new_n996), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT61), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n969), .A2(new_n941), .A3(new_n976), .A4(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT115), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1058));
  INV_X1    g633(.A(G1956), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g635(.A(G299), .B(KEYINPUT57), .Z(new_n1061));
  AND3_X1   g636(.A1(new_n1060), .A2(KEYINPUT116), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT116), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1054), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n760), .B1(new_n970), .B2(new_n972), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n997), .B(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n725), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n819), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1021), .A2(new_n947), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(G1341), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1069), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n544), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT121), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1075), .A2(new_n819), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1065), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1057), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1061), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT122), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1060), .A2(new_n1091), .A3(new_n1061), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1086), .A2(new_n1090), .A3(KEYINPUT61), .A4(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1066), .A2(new_n1074), .A3(new_n1085), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n819), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(new_n1065), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT119), .B1(new_n1064), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n1098));
  OAI221_X1 g673(.A(new_n1098), .B1(new_n1095), .B2(new_n1065), .C1(new_n1063), .C2(new_n1062), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1053), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1045), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1104), .B2(G8), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1051), .B(new_n1106), .C1(new_n1107), .C2(new_n1048), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT62), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1050), .A2(new_n1110), .A3(new_n1051), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n984), .A2(new_n1036), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI211_X1 g688(.A(G1976), .B(G288), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G305), .A2(G1981), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1024), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1116), .A2(new_n998), .B1(new_n1117), .B2(new_n1017), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1025), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G168), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1119), .B(new_n1120), .C1(new_n1036), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n1124));
  OAI21_X1  g699(.A(G8), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1019), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1127), .A2(KEYINPUT63), .A3(G168), .A4(new_n1121), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1131));
  NOR4_X1   g706(.A1(new_n1043), .A2(new_n1120), .A3(new_n1025), .A4(G286), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(KEYINPUT114), .A3(new_n1132), .A4(new_n1127), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1123), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1035), .A2(new_n1019), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1131), .A2(new_n1135), .A3(G168), .A4(new_n1121), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1119), .B1(new_n1136), .B2(new_n1120), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1113), .B(new_n1118), .C1(new_n1134), .C2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n954), .B1(new_n1101), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G290), .A2(G1986), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT48), .B1(new_n1140), .B2(new_n943), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1140), .A2(KEYINPUT48), .A3(new_n943), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1141), .B(new_n1142), .C1(new_n952), .C2(new_n943), .ZN(new_n1143));
  INV_X1    g718(.A(new_n946), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n943), .B1(new_n1144), .B2(new_n745), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT46), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n943), .B2(new_n947), .ZN(new_n1147));
  NOR4_X1   g722(.A1(new_n941), .A2(new_n942), .A3(KEYINPUT46), .A4(G1996), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1145), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT47), .Z(new_n1150));
  NAND2_X1  g725(.A1(new_n946), .A2(new_n948), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n945), .B1(new_n1151), .B2(new_n950), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n1143), .B(new_n1150), .C1(new_n943), .C2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1139), .A2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g729(.A(G229), .B1(new_n869), .B2(new_n872), .ZN(new_n1156));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n1157));
  NOR2_X1   g731(.A1(G227), .A2(new_n461), .ZN(new_n1158));
  AND3_X1   g732(.A1(new_n653), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n653), .B2(new_n1158), .ZN(new_n1160));
  OAI21_X1  g734(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AND2_X1   g735(.A1(new_n923), .A2(new_n926), .ZN(new_n1162));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n931), .B2(new_n1162), .ZN(G308));
  OAI211_X1 g737(.A(new_n932), .B(new_n1156), .C1(new_n1160), .C2(new_n1159), .ZN(G225));
endmodule


