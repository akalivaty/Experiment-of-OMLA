

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789;

  XNOR2_X1 U381 ( .A(n634), .B(n633), .ZN(n708) );
  AND2_X1 U382 ( .A1(n374), .A2(n373), .ZN(n372) );
  BUF_X1 U383 ( .A(G107), .Z(n358) );
  XNOR2_X1 U384 ( .A(n488), .B(n487), .ZN(n677) );
  XNOR2_X2 U385 ( .A(n357), .B(KEYINPUT64), .ZN(n386) );
  NAND2_X2 U386 ( .A1(n643), .A2(n642), .ZN(n357) );
  NOR2_X1 U387 ( .A1(G953), .A2(G237), .ZN(n532) );
  XNOR2_X1 U388 ( .A(n599), .B(KEYINPUT1), .ZN(n551) );
  OR2_X1 U389 ( .A1(n690), .A2(G902), .ZN(n482) );
  XNOR2_X1 U390 ( .A(n615), .B(n616), .ZN(n788) );
  AND2_X4 U391 ( .A1(n386), .A2(n385), .ZN(n699) );
  XNOR2_X2 U392 ( .A(n485), .B(n484), .ZN(n732) );
  NOR2_X2 U393 ( .A1(n391), .A2(n575), .ZN(n389) );
  XNOR2_X2 U394 ( .A(n777), .B(G146), .ZN(n480) );
  NOR2_X2 U395 ( .A1(n788), .A2(n787), .ZN(n621) );
  NAND2_X1 U396 ( .A1(n422), .A2(n417), .ZN(n682) );
  AND2_X1 U397 ( .A1(n576), .A2(n561), .ZN(n562) );
  XNOR2_X2 U398 ( .A(n476), .B(n675), .ZN(n497) );
  BUF_X1 U399 ( .A(n639), .Z(n359) );
  XNOR2_X1 U400 ( .A(n509), .B(n508), .ZN(n360) );
  XNOR2_X1 U401 ( .A(n509), .B(n508), .ZN(n602) );
  XOR2_X1 U402 ( .A(KEYINPUT62), .B(n690), .Z(n691) );
  XNOR2_X1 U403 ( .A(n558), .B(n557), .ZN(n576) );
  XNOR2_X1 U404 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n552) );
  NAND2_X1 U405 ( .A1(n604), .A2(n375), .ZN(n373) );
  NAND2_X1 U406 ( .A1(n361), .A2(n367), .ZN(n392) );
  XNOR2_X1 U407 ( .A(G902), .B(KEYINPUT15), .ZN(n500) );
  NOR2_X1 U408 ( .A1(n428), .A2(n506), .ZN(n427) );
  AND2_X1 U409 ( .A1(G953), .A2(G902), .ZN(n512) );
  NAND2_X1 U410 ( .A1(G237), .A2(G234), .ZN(n510) );
  XNOR2_X1 U411 ( .A(G131), .B(KEYINPUT4), .ZN(n443) );
  INV_X1 U412 ( .A(n732), .ZN(n396) );
  NOR2_X1 U413 ( .A1(n567), .A2(n364), .ZN(n402) );
  AND2_X1 U414 ( .A1(n401), .A2(n625), .ZN(n400) );
  INV_X1 U415 ( .A(n435), .ZN(n421) );
  NAND2_X1 U416 ( .A1(n549), .A2(n420), .ZN(n419) );
  AND2_X1 U417 ( .A1(n411), .A2(n408), .ZN(n406) );
  AND2_X1 U418 ( .A1(n409), .A2(n413), .ZN(n408) );
  NAND2_X1 U419 ( .A1(n410), .A2(KEYINPUT118), .ZN(n409) );
  NAND2_X1 U420 ( .A1(n371), .A2(n370), .ZN(n369) );
  INV_X1 U421 ( .A(KEYINPUT106), .ZN(n387) );
  INV_X1 U422 ( .A(G237), .ZN(n501) );
  XOR2_X1 U423 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n449) );
  INV_X1 U424 ( .A(G902), .ZN(n445) );
  XOR2_X1 U425 ( .A(G143), .B(G140), .Z(n534) );
  INV_X1 U426 ( .A(KEYINPUT10), .ZN(n462) );
  XOR2_X1 U427 ( .A(G104), .B(G131), .Z(n537) );
  XNOR2_X1 U428 ( .A(KEYINPUT98), .B(KEYINPUT12), .ZN(n530) );
  XOR2_X1 U429 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n531) );
  XOR2_X1 U430 ( .A(G140), .B(G137), .Z(n463) );
  XNOR2_X1 U431 ( .A(G146), .B(G125), .ZN(n495) );
  XNOR2_X1 U432 ( .A(KEYINPUT78), .B(KEYINPUT4), .ZN(n494) );
  NAND2_X1 U433 ( .A1(n504), .A2(n641), .ZN(n432) );
  NAND2_X1 U434 ( .A1(n431), .A2(n500), .ZN(n430) );
  INV_X1 U435 ( .A(n504), .ZN(n431) );
  XNOR2_X1 U436 ( .A(n516), .B(KEYINPUT0), .ZN(n566) );
  XOR2_X1 U437 ( .A(KEYINPUT5), .B(G137), .Z(n472) );
  XNOR2_X1 U438 ( .A(G116), .B(G113), .ZN(n474) );
  XNOR2_X1 U439 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U440 ( .A(G128), .B(G119), .ZN(n456) );
  XOR2_X1 U441 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n521) );
  XNOR2_X1 U442 ( .A(G122), .B(KEYINPUT7), .ZN(n520) );
  INV_X1 U443 ( .A(G134), .ZN(n442) );
  NAND2_X1 U444 ( .A1(n641), .A2(KEYINPUT2), .ZN(n642) );
  NOR2_X1 U445 ( .A1(n646), .A2(n714), .ZN(n717) );
  XNOR2_X1 U446 ( .A(n415), .B(KEYINPUT86), .ZN(n646) );
  XNOR2_X1 U447 ( .A(n438), .B(n437), .ZN(n439) );
  INV_X1 U448 ( .A(KEYINPUT91), .ZN(n437) );
  INV_X1 U449 ( .A(n753), .ZN(n410) );
  XNOR2_X1 U450 ( .A(n384), .B(n388), .ZN(n663) );
  INV_X1 U451 ( .A(KEYINPUT31), .ZN(n388) );
  NOR2_X1 U452 ( .A1(n567), .A2(n728), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n381), .B(KEYINPUT77), .ZN(n628) );
  XNOR2_X1 U454 ( .A(n543), .B(n379), .ZN(n571) );
  XNOR2_X1 U455 ( .A(n544), .B(G475), .ZN(n379) );
  XNOR2_X1 U456 ( .A(n656), .B(KEYINPUT59), .ZN(n657) );
  XNOR2_X1 U457 ( .A(n648), .B(n649), .ZN(n650) );
  NAND2_X1 U458 ( .A1(n652), .A2(G953), .ZN(n697) );
  NAND2_X1 U459 ( .A1(n399), .A2(n398), .ZN(n545) );
  AND2_X1 U460 ( .A1(n397), .A2(n400), .ZN(n399) );
  NAND2_X1 U461 ( .A1(n396), .A2(n402), .ZN(n398) );
  AND2_X1 U462 ( .A1(n425), .A2(n423), .ZN(n422) );
  NOR2_X1 U463 ( .A1(n421), .A2(n419), .ZN(n418) );
  NAND2_X1 U464 ( .A1(n406), .A2(n405), .ZN(n404) );
  NAND2_X1 U465 ( .A1(n407), .A2(KEYINPUT118), .ZN(n405) );
  OR2_X1 U466 ( .A1(n689), .A2(n576), .ZN(n361) );
  INV_X1 U467 ( .A(n500), .ZN(n641) );
  AND2_X1 U468 ( .A1(n429), .A2(n432), .ZN(n362) );
  AND2_X1 U469 ( .A1(n707), .A2(KEYINPUT2), .ZN(n363) );
  XOR2_X1 U470 ( .A(KEYINPUT79), .B(KEYINPUT34), .Z(n364) );
  XOR2_X1 U471 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n365) );
  XNOR2_X1 U472 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n366) );
  AND2_X1 U473 ( .A1(n559), .A2(KEYINPUT88), .ZN(n367) );
  XNOR2_X1 U474 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n368) );
  INV_X1 U475 ( .A(KEYINPUT118), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n378), .B(KEYINPUT45), .ZN(n645) );
  BUF_X1 U477 ( .A(n645), .Z(n668) );
  NAND2_X1 U478 ( .A1(n372), .A2(n369), .ZN(n377) );
  NOR2_X1 U479 ( .A1(n604), .A2(n375), .ZN(n370) );
  INV_X1 U480 ( .A(n572), .ZN(n371) );
  NAND2_X1 U481 ( .A1(n572), .A2(n375), .ZN(n374) );
  INV_X1 U482 ( .A(KEYINPUT105), .ZN(n375) );
  XNOR2_X1 U483 ( .A(n376), .B(n387), .ZN(n383) );
  NAND2_X1 U484 ( .A1(n377), .A2(n666), .ZN(n376) );
  BUF_X2 U485 ( .A(n566), .Z(n567) );
  NAND2_X1 U486 ( .A1(n390), .A2(n389), .ZN(n378) );
  BUF_X1 U487 ( .A(n663), .Z(n380) );
  NAND2_X1 U488 ( .A1(n614), .A2(n613), .ZN(n381) );
  NOR2_X2 U489 ( .A1(n663), .A2(n757), .ZN(n572) );
  OR2_X2 U490 ( .A1(n702), .A2(G902), .ZN(n395) );
  NAND2_X1 U491 ( .A1(n383), .A2(n416), .ZN(n391) );
  INV_X1 U492 ( .A(n717), .ZN(n385) );
  INV_X1 U493 ( .A(n556), .ZN(n553) );
  NAND2_X1 U494 ( .A1(n556), .A2(n552), .ZN(n425) );
  XNOR2_X2 U495 ( .A(n548), .B(n366), .ZN(n556) );
  XNOR2_X1 U496 ( .A(n538), .B(n522), .ZN(n488) );
  XNOR2_X2 U497 ( .A(G122), .B(G113), .ZN(n538) );
  NAND2_X1 U498 ( .A1(n577), .A2(KEYINPUT65), .ZN(n416) );
  AND2_X2 U499 ( .A1(n429), .A2(n427), .ZN(n426) );
  XNOR2_X2 U500 ( .A(KEYINPUT104), .B(n569), .ZN(n768) );
  AND2_X1 U501 ( .A1(n609), .A2(n608), .ZN(n614) );
  AND2_X2 U502 ( .A1(n708), .A2(n707), .ZN(n644) );
  NAND2_X1 U503 ( .A1(n628), .A2(n734), .ZN(n403) );
  NOR2_X1 U504 ( .A1(n656), .A2(G902), .ZN(n543) );
  XNOR2_X1 U505 ( .A(n541), .B(n542), .ZN(n656) );
  OR2_X2 U506 ( .A1(n737), .A2(n722), .ZN(n547) );
  NAND2_X1 U507 ( .A1(n393), .A2(n392), .ZN(n390) );
  OR2_X2 U508 ( .A1(n563), .A2(n562), .ZN(n393) );
  NOR2_X2 U509 ( .A1(n551), .A2(n720), .ZN(n565) );
  XNOR2_X2 U510 ( .A(n394), .B(KEYINPUT69), .ZN(n720) );
  NOR2_X2 U511 ( .A1(n550), .A2(n722), .ZN(n394) );
  XNOR2_X2 U512 ( .A(n469), .B(n468), .ZN(n550) );
  XNOR2_X2 U513 ( .A(n395), .B(n447), .ZN(n599) );
  NAND2_X1 U514 ( .A1(n732), .A2(n364), .ZN(n397) );
  NAND2_X1 U515 ( .A1(n567), .A2(n364), .ZN(n401) );
  NAND2_X1 U516 ( .A1(n639), .A2(n768), .ZN(n615) );
  XNOR2_X2 U517 ( .A(n403), .B(n365), .ZN(n639) );
  XNOR2_X1 U518 ( .A(n404), .B(n368), .ZN(G75) );
  INV_X1 U519 ( .A(n754), .ZN(n407) );
  NAND2_X1 U520 ( .A1(n754), .A2(n412), .ZN(n411) );
  AND2_X1 U521 ( .A1(n753), .A2(n414), .ZN(n412) );
  INV_X4 U522 ( .A(G953), .ZN(n413) );
  NAND2_X1 U523 ( .A1(n708), .A2(n363), .ZN(n415) );
  OR2_X1 U524 ( .A1(n718), .A2(n717), .ZN(n754) );
  NOR2_X1 U525 ( .A1(n714), .A2(n775), .ZN(n709) );
  XNOR2_X2 U526 ( .A(n492), .B(n442), .ZN(n518) );
  XNOR2_X2 U527 ( .A(n518), .B(n443), .ZN(n777) );
  AND2_X1 U528 ( .A1(n553), .A2(n549), .ZN(n436) );
  NAND2_X1 U529 ( .A1(n553), .A2(n418), .ZN(n417) );
  INV_X1 U530 ( .A(n552), .ZN(n420) );
  NAND2_X1 U531 ( .A1(n424), .A2(n552), .ZN(n423) );
  NAND2_X1 U532 ( .A1(n435), .A2(n549), .ZN(n424) );
  XNOR2_X1 U533 ( .A(n499), .B(n498), .ZN(n647) );
  OR2_X2 U534 ( .A1(n647), .A2(n430), .ZN(n429) );
  NAND2_X1 U535 ( .A1(n362), .A2(n433), .ZN(n591) );
  NAND2_X2 U536 ( .A1(n426), .A2(n433), .ZN(n509) );
  INV_X1 U537 ( .A(n432), .ZN(n428) );
  NAND2_X1 U538 ( .A1(n647), .A2(n504), .ZN(n433) );
  INV_X1 U539 ( .A(n684), .ZN(n685) );
  XNOR2_X1 U540 ( .A(n458), .B(n457), .ZN(n461) );
  XNOR2_X2 U541 ( .A(KEYINPUT68), .B(G101), .ZN(n476) );
  XNOR2_X2 U542 ( .A(G110), .B(G104), .ZN(n675) );
  XNOR2_X2 U543 ( .A(G143), .B(G128), .ZN(n492) );
  XNOR2_X2 U544 ( .A(G116), .B(G107), .ZN(n522) );
  XOR2_X1 U545 ( .A(n440), .B(n439), .Z(n434) );
  AND2_X1 U546 ( .A1(n723), .A2(n573), .ZN(n435) );
  INV_X1 U547 ( .A(KEYINPUT107), .ZN(n470) );
  XNOR2_X1 U548 ( .A(KEYINPUT48), .B(KEYINPUT70), .ZN(n633) );
  INV_X1 U549 ( .A(KEYINPUT23), .ZN(n455) );
  BUF_X1 U550 ( .A(n732), .Z(n750) );
  INV_X1 U551 ( .A(n463), .ZN(n440) );
  NAND2_X1 U552 ( .A1(n413), .A2(G227), .ZN(n438) );
  XOR2_X1 U553 ( .A(n358), .B(n497), .Z(n441) );
  XNOR2_X1 U554 ( .A(n434), .B(n441), .ZN(n444) );
  XNOR2_X1 U555 ( .A(n444), .B(n480), .ZN(n702) );
  XNOR2_X1 U556 ( .A(G469), .B(KEYINPUT73), .ZN(n446) );
  XNOR2_X1 U557 ( .A(n446), .B(KEYINPUT72), .ZN(n447) );
  NAND2_X1 U558 ( .A1(G234), .A2(n500), .ZN(n448) );
  XNOR2_X1 U559 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U560 ( .A(KEYINPUT94), .B(n450), .ZN(n465) );
  NAND2_X1 U561 ( .A1(n465), .A2(G221), .ZN(n452) );
  XNOR2_X1 U562 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n451) );
  XNOR2_X1 U563 ( .A(n452), .B(n451), .ZN(n722) );
  XOR2_X1 U564 ( .A(KEYINPUT24), .B(KEYINPUT83), .Z(n454) );
  XNOR2_X1 U565 ( .A(G110), .B(KEYINPUT92), .ZN(n453) );
  XNOR2_X1 U566 ( .A(n454), .B(n453), .ZN(n458) );
  AND2_X1 U567 ( .A1(G234), .A2(n413), .ZN(n459) );
  XNOR2_X1 U568 ( .A(KEYINPUT8), .B(n459), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n517), .A2(G221), .ZN(n460) );
  XNOR2_X1 U570 ( .A(n461), .B(n460), .ZN(n464) );
  XNOR2_X1 U571 ( .A(n495), .B(n462), .ZN(n540) );
  XNOR2_X1 U572 ( .A(n463), .B(n540), .ZN(n776) );
  XNOR2_X1 U573 ( .A(n464), .B(n776), .ZN(n696) );
  NAND2_X1 U574 ( .A1(n696), .A2(n445), .ZN(n469) );
  NAND2_X1 U575 ( .A1(n465), .A2(G217), .ZN(n467) );
  XOR2_X1 U576 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n466) );
  XNOR2_X1 U577 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U578 ( .A(n565), .B(n470), .ZN(n483) );
  NAND2_X1 U579 ( .A1(G210), .A2(n532), .ZN(n471) );
  XNOR2_X1 U580 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X2 U581 ( .A(KEYINPUT3), .B(G119), .ZN(n486) );
  XNOR2_X1 U582 ( .A(n486), .B(n473), .ZN(n478) );
  XNOR2_X1 U583 ( .A(KEYINPUT76), .B(n474), .ZN(n475) );
  XNOR2_X1 U584 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U585 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U586 ( .A(n480), .B(n479), .ZN(n690) );
  INV_X1 U587 ( .A(G472), .ZN(n481) );
  XNOR2_X2 U588 ( .A(n482), .B(n481), .ZN(n564) );
  XNOR2_X1 U589 ( .A(n564), .B(KEYINPUT6), .ZN(n589) );
  NAND2_X1 U590 ( .A1(n483), .A2(n589), .ZN(n485) );
  XOR2_X1 U591 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n484) );
  XNOR2_X1 U592 ( .A(n486), .B(KEYINPUT16), .ZN(n487) );
  XNOR2_X1 U593 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n490) );
  NAND2_X1 U594 ( .A1(n413), .A2(G224), .ZN(n489) );
  XNOR2_X1 U595 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U596 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U597 ( .A(n677), .B(n493), .ZN(n499) );
  XNOR2_X1 U598 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U599 ( .A(n497), .B(n496), .ZN(n498) );
  NAND2_X1 U600 ( .A1(n445), .A2(n501), .ZN(n505) );
  NAND2_X1 U601 ( .A1(n505), .A2(G210), .ZN(n503) );
  XNOR2_X1 U602 ( .A(KEYINPUT80), .B(KEYINPUT90), .ZN(n502) );
  XNOR2_X1 U603 ( .A(n503), .B(n502), .ZN(n504) );
  NAND2_X1 U604 ( .A1(n505), .A2(G214), .ZN(n733) );
  INV_X1 U605 ( .A(n733), .ZN(n506) );
  INV_X1 U606 ( .A(KEYINPUT67), .ZN(n507) );
  XNOR2_X1 U607 ( .A(n507), .B(KEYINPUT19), .ZN(n508) );
  XNOR2_X1 U608 ( .A(n510), .B(KEYINPUT14), .ZN(n746) );
  INV_X1 U609 ( .A(G898), .ZN(n511) );
  NAND2_X1 U610 ( .A1(n512), .A2(n511), .ZN(n513) );
  NAND2_X1 U611 ( .A1(n413), .A2(G952), .ZN(n582) );
  NAND2_X1 U612 ( .A1(n513), .A2(n582), .ZN(n514) );
  AND2_X1 U613 ( .A1(n746), .A2(n514), .ZN(n515) );
  NAND2_X1 U614 ( .A1(n602), .A2(n515), .ZN(n516) );
  XNOR2_X1 U615 ( .A(KEYINPUT103), .B(KEYINPUT102), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n517), .A2(G217), .ZN(n519) );
  XNOR2_X1 U617 ( .A(n519), .B(n518), .ZN(n526) );
  XNOR2_X1 U618 ( .A(n521), .B(n520), .ZN(n524) );
  XOR2_X1 U619 ( .A(KEYINPUT100), .B(n522), .Z(n523) );
  XNOR2_X1 U620 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U621 ( .A(n526), .B(n525), .ZN(n684) );
  NOR2_X1 U622 ( .A1(n684), .A2(G902), .ZN(n527) );
  XNOR2_X1 U623 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U624 ( .A(n529), .B(G478), .ZN(n570) );
  INV_X1 U625 ( .A(n570), .ZN(n546) );
  XNOR2_X1 U626 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n544) );
  XNOR2_X1 U627 ( .A(n531), .B(n530), .ZN(n536) );
  NAND2_X1 U628 ( .A1(n532), .A2(G214), .ZN(n533) );
  XNOR2_X1 U629 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U630 ( .A(n535), .B(n536), .ZN(n542) );
  XNOR2_X1 U631 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U632 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U633 ( .A1(n546), .A2(n571), .ZN(n625) );
  XNOR2_X2 U634 ( .A(n545), .B(KEYINPUT35), .ZN(n689) );
  NAND2_X1 U635 ( .A1(n546), .A2(n571), .ZN(n737) );
  NOR2_X2 U636 ( .A1(n566), .A2(n547), .ZN(n548) );
  INV_X1 U637 ( .A(n589), .ZN(n549) );
  BUF_X1 U638 ( .A(n550), .Z(n723) );
  BUF_X2 U639 ( .A(n551), .Z(n719) );
  INV_X1 U640 ( .A(n719), .ZN(n573) );
  AND2_X1 U641 ( .A1(n723), .A2(n719), .ZN(n554) );
  NAND2_X1 U642 ( .A1(n554), .A2(n564), .ZN(n555) );
  OR2_X1 U643 ( .A1(n556), .A2(n555), .ZN(n665) );
  NAND2_X1 U644 ( .A1(n682), .A2(n665), .ZN(n558) );
  INV_X1 U645 ( .A(KEYINPUT89), .ZN(n557) );
  NOR2_X1 U646 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n559) );
  NAND2_X1 U647 ( .A1(n689), .A2(KEYINPUT88), .ZN(n560) );
  NAND2_X1 U648 ( .A1(n560), .A2(KEYINPUT44), .ZN(n563) );
  INV_X1 U649 ( .A(KEYINPUT65), .ZN(n561) );
  NOR2_X1 U650 ( .A1(n689), .A2(KEYINPUT88), .ZN(n575) );
  INV_X1 U651 ( .A(n564), .ZN(n610) );
  NAND2_X1 U652 ( .A1(n565), .A2(n610), .ZN(n728) );
  NOR2_X1 U653 ( .A1(n720), .A2(n599), .ZN(n609) );
  NAND2_X1 U654 ( .A1(n609), .A2(n564), .ZN(n568) );
  NOR2_X1 U655 ( .A1(n568), .A2(n567), .ZN(n757) );
  NOR2_X1 U656 ( .A1(n571), .A2(n570), .ZN(n569) );
  AND2_X1 U657 ( .A1(n571), .A2(n570), .ZN(n762) );
  NOR2_X1 U658 ( .A1(n768), .A2(n762), .ZN(n739) );
  XNOR2_X1 U659 ( .A(n739), .B(KEYINPUT82), .ZN(n604) );
  NOR2_X1 U660 ( .A1(n723), .A2(n573), .ZN(n574) );
  NAND2_X1 U661 ( .A1(n436), .A2(n574), .ZN(n666) );
  INV_X1 U662 ( .A(n576), .ZN(n577) );
  NAND2_X1 U663 ( .A1(n645), .A2(n641), .ZN(n578) );
  XNOR2_X1 U664 ( .A(n578), .B(KEYINPUT85), .ZN(n640) );
  NAND2_X1 U665 ( .A1(G902), .A2(n746), .ZN(n579) );
  NOR2_X1 U666 ( .A1(G900), .A2(n579), .ZN(n580) );
  NAND2_X1 U667 ( .A1(G953), .A2(n580), .ZN(n581) );
  XOR2_X1 U668 ( .A(KEYINPUT108), .B(n581), .Z(n585) );
  INV_X1 U669 ( .A(n746), .ZN(n583) );
  NOR2_X1 U670 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U671 ( .A1(n585), .A2(n584), .ZN(n607) );
  NOR2_X1 U672 ( .A1(n607), .A2(n722), .ZN(n586) );
  XOR2_X1 U673 ( .A(KEYINPUT71), .B(n586), .Z(n596) );
  NAND2_X1 U674 ( .A1(n596), .A2(n733), .ZN(n588) );
  NAND2_X1 U675 ( .A1(n723), .A2(n768), .ZN(n587) );
  NOR2_X1 U676 ( .A1(n588), .A2(n587), .ZN(n590) );
  AND2_X1 U677 ( .A1(n590), .A2(n589), .ZN(n635) );
  INV_X1 U678 ( .A(n591), .ZN(n592) );
  NAND2_X1 U679 ( .A1(n635), .A2(n592), .ZN(n593) );
  XNOR2_X1 U680 ( .A(n593), .B(KEYINPUT36), .ZN(n594) );
  XNOR2_X1 U681 ( .A(n594), .B(KEYINPUT112), .ZN(n595) );
  NOR2_X1 U682 ( .A1(n719), .A2(n595), .ZN(n771) );
  NAND2_X1 U683 ( .A1(n723), .A2(n596), .ZN(n597) );
  NOR2_X1 U684 ( .A1(n564), .A2(n597), .ZN(n598) );
  XNOR2_X1 U685 ( .A(n598), .B(KEYINPUT28), .ZN(n601) );
  INV_X1 U686 ( .A(n599), .ZN(n600) );
  NAND2_X1 U687 ( .A1(n601), .A2(n600), .ZN(n619) );
  INV_X1 U688 ( .A(n619), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n603), .A2(n360), .ZN(n761) );
  OR2_X1 U690 ( .A1(n604), .A2(n761), .ZN(n605) );
  NOR2_X1 U691 ( .A1(KEYINPUT47), .A2(n605), .ZN(n606) );
  NOR2_X1 U692 ( .A1(n771), .A2(n606), .ZN(n623) );
  INV_X1 U693 ( .A(KEYINPUT40), .ZN(n616) );
  INV_X1 U694 ( .A(n607), .ZN(n608) );
  XOR2_X1 U695 ( .A(KEYINPUT30), .B(KEYINPUT110), .Z(n612) );
  NAND2_X1 U696 ( .A1(n610), .A2(n733), .ZN(n611) );
  XNOR2_X1 U697 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U698 ( .A(n591), .B(KEYINPUT38), .ZN(n734) );
  NAND2_X1 U699 ( .A1(n734), .A2(n733), .ZN(n738) );
  NOR2_X1 U700 ( .A1(n738), .A2(n737), .ZN(n618) );
  XOR2_X1 U701 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n617) );
  XNOR2_X1 U702 ( .A(n618), .B(n617), .ZN(n749) );
  NOR2_X1 U703 ( .A1(n619), .A2(n749), .ZN(n620) );
  XNOR2_X1 U704 ( .A(KEYINPUT42), .B(n620), .ZN(n787) );
  XNOR2_X1 U705 ( .A(n621), .B(KEYINPUT46), .ZN(n622) );
  NAND2_X1 U706 ( .A1(n622), .A2(n623), .ZN(n632) );
  OR2_X1 U707 ( .A1(n761), .A2(n739), .ZN(n624) );
  NAND2_X1 U708 ( .A1(n624), .A2(KEYINPUT47), .ZN(n629) );
  INV_X1 U709 ( .A(n625), .ZN(n626) );
  NOR2_X1 U710 ( .A1(n626), .A2(n591), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n767) );
  NAND2_X1 U712 ( .A1(n629), .A2(n767), .ZN(n630) );
  XOR2_X1 U713 ( .A(n630), .B(KEYINPUT81), .Z(n631) );
  NOR2_X2 U714 ( .A1(n632), .A2(n631), .ZN(n634) );
  XOR2_X1 U715 ( .A(KEYINPUT109), .B(n635), .Z(n636) );
  NAND2_X1 U716 ( .A1(n636), .A2(n719), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n637), .B(KEYINPUT43), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n638), .A2(n591), .ZN(n667) );
  NAND2_X1 U719 ( .A1(n762), .A2(n359), .ZN(n773) );
  AND2_X1 U720 ( .A1(n667), .A2(n773), .ZN(n707) );
  NAND2_X1 U721 ( .A1(n640), .A2(n644), .ZN(n643) );
  INV_X1 U722 ( .A(n668), .ZN(n714) );
  NAND2_X1 U723 ( .A1(n699), .A2(G210), .ZN(n651) );
  BUF_X1 U724 ( .A(n647), .Z(n648) );
  XNOR2_X1 U725 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n649) );
  XNOR2_X1 U726 ( .A(n651), .B(n650), .ZN(n653) );
  INV_X1 U727 ( .A(G952), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n697), .ZN(n655) );
  INV_X1 U729 ( .A(KEYINPUT56), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n655), .B(n654), .ZN(G51) );
  NAND2_X1 U731 ( .A1(n699), .A2(G475), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n659), .A2(n697), .ZN(n661) );
  INV_X1 U734 ( .A(KEYINPUT60), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n661), .B(n660), .ZN(G60) );
  NAND2_X1 U736 ( .A1(n380), .A2(n762), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n662), .B(G116), .ZN(G18) );
  NAND2_X1 U738 ( .A1(n380), .A2(n768), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n664), .B(G113), .ZN(G15) );
  XNOR2_X1 U740 ( .A(n665), .B(G110), .ZN(G12) );
  XNOR2_X1 U741 ( .A(n666), .B(G101), .ZN(G3) );
  XNOR2_X1 U742 ( .A(n667), .B(G140), .ZN(G42) );
  NAND2_X1 U743 ( .A1(n668), .A2(n413), .ZN(n673) );
  NAND2_X1 U744 ( .A1(G953), .A2(G224), .ZN(n669) );
  XNOR2_X1 U745 ( .A(KEYINPUT61), .B(n669), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n670), .A2(G898), .ZN(n671) );
  XNOR2_X1 U747 ( .A(n671), .B(KEYINPUT122), .ZN(n672) );
  NAND2_X1 U748 ( .A1(n673), .A2(n672), .ZN(n681) );
  XOR2_X1 U749 ( .A(G101), .B(KEYINPUT123), .Z(n674) );
  XNOR2_X1 U750 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U751 ( .A(n677), .B(n676), .ZN(n679) );
  NOR2_X1 U752 ( .A1(n413), .A2(G898), .ZN(n678) );
  NOR2_X1 U753 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U754 ( .A(n681), .B(n680), .ZN(G69) );
  BUF_X1 U755 ( .A(n682), .Z(n683) );
  XNOR2_X1 U756 ( .A(n683), .B(G119), .ZN(G21) );
  NAND2_X1 U757 ( .A1(n699), .A2(G478), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U759 ( .A1(n687), .A2(n697), .ZN(n688) );
  XNOR2_X1 U760 ( .A(n688), .B(KEYINPUT121), .ZN(G63) );
  XOR2_X1 U761 ( .A(n689), .B(G122), .Z(G24) );
  NAND2_X1 U762 ( .A1(n699), .A2(G472), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n692), .B(n691), .ZN(n693) );
  NAND2_X1 U764 ( .A1(n693), .A2(n697), .ZN(n694) );
  XNOR2_X1 U765 ( .A(n694), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U766 ( .A1(n699), .A2(G217), .ZN(n695) );
  XOR2_X1 U767 ( .A(n696), .B(n695), .Z(n698) );
  INV_X1 U768 ( .A(n697), .ZN(n705) );
  NOR2_X1 U769 ( .A1(n698), .A2(n705), .ZN(G66) );
  NAND2_X1 U770 ( .A1(n699), .A2(G469), .ZN(n704) );
  XOR2_X1 U771 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n700) );
  XNOR2_X1 U772 ( .A(n700), .B(KEYINPUT58), .ZN(n701) );
  XNOR2_X1 U773 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U774 ( .A(n704), .B(n703), .ZN(n706) );
  NOR2_X1 U775 ( .A1(n706), .A2(n705), .ZN(G54) );
  NAND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n775) );
  NOR2_X1 U777 ( .A1(n709), .A2(KEYINPUT2), .ZN(n711) );
  INV_X1 U778 ( .A(KEYINPUT84), .ZN(n710) );
  NOR2_X1 U779 ( .A1(n711), .A2(n710), .ZN(n716) );
  NOR2_X1 U780 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n775), .A2(n712), .ZN(n713) );
  NOR2_X1 U782 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n718) );
  NAND2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U785 ( .A(n721), .B(KEYINPUT50), .ZN(n727) );
  NAND2_X1 U786 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U787 ( .A(KEYINPUT49), .B(n724), .ZN(n725) );
  NOR2_X1 U788 ( .A1(n610), .A2(n725), .ZN(n726) );
  NAND2_X1 U789 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U790 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U791 ( .A(KEYINPUT51), .B(n730), .ZN(n731) );
  NOR2_X1 U792 ( .A1(n749), .A2(n731), .ZN(n744) );
  NOR2_X1 U793 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U794 ( .A(KEYINPUT117), .B(n735), .Z(n736) );
  NOR2_X1 U795 ( .A1(n737), .A2(n736), .ZN(n741) );
  NOR2_X1 U796 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U797 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U798 ( .A1(n750), .A2(n742), .ZN(n743) );
  NOR2_X1 U799 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U800 ( .A(n745), .B(KEYINPUT52), .ZN(n748) );
  NAND2_X1 U801 ( .A1(n746), .A2(G952), .ZN(n747) );
  NOR2_X1 U802 ( .A1(n748), .A2(n747), .ZN(n752) );
  NOR2_X1 U803 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U804 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U805 ( .A(G104), .B(KEYINPUT113), .Z(n756) );
  NAND2_X1 U806 ( .A1(n757), .A2(n768), .ZN(n755) );
  XNOR2_X1 U807 ( .A(n756), .B(n755), .ZN(G6) );
  XOR2_X1 U808 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n759) );
  NAND2_X1 U809 ( .A1(n757), .A2(n762), .ZN(n758) );
  XNOR2_X1 U810 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U811 ( .A(n358), .B(n760), .ZN(G9) );
  XOR2_X1 U812 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n764) );
  INV_X1 U813 ( .A(n761), .ZN(n769) );
  NAND2_X1 U814 ( .A1(n769), .A2(n762), .ZN(n763) );
  XNOR2_X1 U815 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U816 ( .A(G128), .B(n765), .ZN(G30) );
  XOR2_X1 U817 ( .A(G143), .B(KEYINPUT115), .Z(n766) );
  XNOR2_X1 U818 ( .A(n767), .B(n766), .ZN(G45) );
  NAND2_X1 U819 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U820 ( .A(n770), .B(G146), .ZN(G48) );
  XNOR2_X1 U821 ( .A(G125), .B(n771), .ZN(n772) );
  XNOR2_X1 U822 ( .A(n772), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U823 ( .A(G134), .B(KEYINPUT116), .ZN(n774) );
  XNOR2_X1 U824 ( .A(n774), .B(n773), .ZN(G36) );
  XNOR2_X1 U825 ( .A(n776), .B(KEYINPUT124), .ZN(n778) );
  XNOR2_X1 U826 ( .A(n778), .B(n777), .ZN(n780) );
  XOR2_X1 U827 ( .A(n644), .B(n780), .Z(n779) );
  NAND2_X1 U828 ( .A1(n779), .A2(n413), .ZN(n785) );
  XNOR2_X1 U829 ( .A(G227), .B(n780), .ZN(n781) );
  NAND2_X1 U830 ( .A1(n781), .A2(G900), .ZN(n782) );
  NAND2_X1 U831 ( .A1(G953), .A2(n782), .ZN(n783) );
  XOR2_X1 U832 ( .A(KEYINPUT125), .B(n783), .Z(n784) );
  NAND2_X1 U833 ( .A1(n785), .A2(n784), .ZN(G72) );
  XOR2_X1 U834 ( .A(G137), .B(KEYINPUT126), .Z(n786) );
  XNOR2_X1 U835 ( .A(n787), .B(n786), .ZN(G39) );
  XNOR2_X1 U836 ( .A(G131), .B(KEYINPUT127), .ZN(n789) );
  XNOR2_X1 U837 ( .A(n789), .B(n788), .ZN(G33) );
endmodule

