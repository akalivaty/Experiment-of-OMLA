

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U557 ( .A1(n543), .A2(n542), .ZN(G160) );
  INV_X1 U558 ( .A(KEYINPUT109), .ZN(n621) );
  INV_X1 U559 ( .A(KEYINPUT31), .ZN(n632) );
  XNOR2_X1 U560 ( .A(KEYINPUT104), .B(KEYINPUT27), .ZN(n636) );
  XNOR2_X1 U561 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U562 ( .A(n620), .ZN(n669) );
  XNOR2_X1 U563 ( .A(n683), .B(KEYINPUT29), .ZN(n684) );
  XNOR2_X1 U564 ( .A(n685), .B(n684), .ZN(n686) );
  XOR2_X1 U565 ( .A(KEYINPUT17), .B(n532), .Z(n915) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n817) );
  INV_X1 U567 ( .A(G651), .ZN(n527) );
  NOR2_X1 U568 ( .A1(G543), .A2(n527), .ZN(n524) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n524), .Z(n813) );
  NAND2_X1 U570 ( .A1(G60), .A2(n813), .ZN(n526) );
  XOR2_X1 U571 ( .A(KEYINPUT0), .B(G543), .Z(n590) );
  NOR2_X1 U572 ( .A1(G651), .A2(n590), .ZN(n814) );
  NAND2_X1 U573 ( .A1(G47), .A2(n814), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n526), .A2(n525), .ZN(n531) );
  NAND2_X1 U575 ( .A1(G85), .A2(n817), .ZN(n529) );
  NOR2_X1 U576 ( .A1(n590), .A2(n527), .ZN(n812) );
  NAND2_X1 U577 ( .A1(G72), .A2(n812), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  OR2_X1 U579 ( .A1(n531), .A2(n530), .ZN(G290) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n532) );
  NAND2_X1 U581 ( .A1(G137), .A2(n915), .ZN(n534) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n912) );
  NAND2_X1 U583 ( .A1(G113), .A2(n912), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n534), .A2(n533), .ZN(n543) );
  INV_X1 U585 ( .A(G2104), .ZN(n537) );
  NOR2_X1 U586 ( .A1(n537), .A2(G2105), .ZN(n535) );
  XNOR2_X2 U587 ( .A(n535), .B(KEYINPUT64), .ZN(n917) );
  NAND2_X1 U588 ( .A1(G101), .A2(n917), .ZN(n536) );
  XOR2_X1 U589 ( .A(n536), .B(KEYINPUT23), .Z(n539) );
  AND2_X1 U590 ( .A1(n537), .A2(G2105), .ZN(n911) );
  NAND2_X1 U591 ( .A1(n911), .A2(G125), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n541) );
  INV_X1 U593 ( .A(KEYINPUT65), .ZN(n540) );
  XNOR2_X1 U594 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U595 ( .A1(G138), .A2(n915), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G102), .A2(n917), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U598 ( .A1(G126), .A2(n911), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G114), .A2(n912), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U601 ( .A1(n549), .A2(n548), .ZN(G164) );
  NAND2_X1 U602 ( .A1(n817), .A2(G89), .ZN(n550) );
  XNOR2_X1 U603 ( .A(KEYINPUT4), .B(n550), .ZN(n553) );
  NAND2_X1 U604 ( .A1(n812), .A2(G76), .ZN(n551) );
  XOR2_X1 U605 ( .A(KEYINPUT79), .B(n551), .Z(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U607 ( .A(n554), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U608 ( .A1(G63), .A2(n813), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G51), .A2(n814), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U611 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U612 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U613 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U614 ( .A1(n814), .A2(G52), .ZN(n561) );
  XNOR2_X1 U615 ( .A(n561), .B(KEYINPUT66), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G64), .A2(n813), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U618 ( .A(KEYINPUT67), .B(n564), .Z(n569) );
  NAND2_X1 U619 ( .A1(G90), .A2(n817), .ZN(n566) );
  NAND2_X1 U620 ( .A1(G77), .A2(n812), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  NOR2_X1 U623 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U624 ( .A(KEYINPUT68), .B(n570), .ZN(G171) );
  NAND2_X1 U625 ( .A1(n813), .A2(G65), .ZN(n571) );
  XOR2_X1 U626 ( .A(KEYINPUT69), .B(n571), .Z(n573) );
  NAND2_X1 U627 ( .A1(n814), .A2(G53), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U629 ( .A(KEYINPUT70), .B(n574), .Z(n578) );
  NAND2_X1 U630 ( .A1(G91), .A2(n817), .ZN(n576) );
  NAND2_X1 U631 ( .A1(G78), .A2(n812), .ZN(n575) );
  AND2_X1 U632 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n578), .A2(n577), .ZN(G299) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G50), .A2(n814), .ZN(n579) );
  XNOR2_X1 U636 ( .A(n579), .B(KEYINPUT84), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G75), .A2(n812), .ZN(n580) );
  XOR2_X1 U638 ( .A(KEYINPUT85), .B(n580), .Z(n581) );
  NAND2_X1 U639 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U640 ( .A1(G62), .A2(n813), .ZN(n584) );
  NAND2_X1 U641 ( .A1(G88), .A2(n817), .ZN(n583) );
  NAND2_X1 U642 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U643 ( .A1(n586), .A2(n585), .ZN(G166) );
  XOR2_X1 U644 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NAND2_X1 U645 ( .A1(G49), .A2(n814), .ZN(n588) );
  NAND2_X1 U646 ( .A1(G74), .A2(G651), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U648 ( .A1(n813), .A2(n589), .ZN(n592) );
  NAND2_X1 U649 ( .A1(n590), .A2(G87), .ZN(n591) );
  NAND2_X1 U650 ( .A1(n592), .A2(n591), .ZN(G288) );
  NAND2_X1 U651 ( .A1(G61), .A2(n813), .ZN(n594) );
  NAND2_X1 U652 ( .A1(G48), .A2(n814), .ZN(n593) );
  NAND2_X1 U653 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U654 ( .A1(n812), .A2(G73), .ZN(n595) );
  XOR2_X1 U655 ( .A(KEYINPUT2), .B(n595), .Z(n596) );
  NOR2_X1 U656 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U657 ( .A1(n817), .A2(G86), .ZN(n598) );
  NAND2_X1 U658 ( .A1(n599), .A2(n598), .ZN(G305) );
  XNOR2_X1 U659 ( .A(G1986), .B(G290), .ZN(n985) );
  NAND2_X1 U660 ( .A1(G160), .A2(G40), .ZN(n617) );
  NOR2_X1 U661 ( .A1(G164), .A2(G1384), .ZN(n618) );
  NOR2_X1 U662 ( .A1(n617), .A2(n618), .ZN(n600) );
  XOR2_X1 U663 ( .A(n600), .B(KEYINPUT91), .Z(n769) );
  NAND2_X1 U664 ( .A1(n985), .A2(n769), .ZN(n601) );
  XNOR2_X1 U665 ( .A(n601), .B(KEYINPUT92), .ZN(n616) );
  XNOR2_X1 U666 ( .A(KEYINPUT95), .B(KEYINPUT36), .ZN(n612) );
  NAND2_X1 U667 ( .A1(G128), .A2(n911), .ZN(n603) );
  NAND2_X1 U668 ( .A1(G116), .A2(n912), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U670 ( .A(KEYINPUT35), .B(n604), .ZN(n610) );
  NAND2_X1 U671 ( .A1(G140), .A2(n915), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G104), .A2(n917), .ZN(n605) );
  NAND2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n608) );
  XOR2_X1 U674 ( .A(KEYINPUT94), .B(KEYINPUT34), .Z(n607) );
  XNOR2_X1 U675 ( .A(n608), .B(n607), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U677 ( .A(n612), .B(n611), .Z(n908) );
  XOR2_X1 U678 ( .A(G2067), .B(KEYINPUT37), .Z(n613) );
  XOR2_X1 U679 ( .A(KEYINPUT93), .B(n613), .Z(n767) );
  NAND2_X1 U680 ( .A1(n908), .A2(n767), .ZN(n614) );
  XNOR2_X1 U681 ( .A(n614), .B(KEYINPUT96), .ZN(n765) );
  INV_X1 U682 ( .A(n765), .ZN(n954) );
  NAND2_X1 U683 ( .A1(n954), .A2(n769), .ZN(n615) );
  NAND2_X1 U684 ( .A1(n616), .A2(n615), .ZN(n735) );
  XOR2_X1 U685 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n625) );
  INV_X1 U686 ( .A(n617), .ZN(n619) );
  NAND2_X1 U687 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U688 ( .A1(G2084), .A2(n620), .ZN(n693) );
  NAND2_X1 U689 ( .A1(G8), .A2(n620), .ZN(n729) );
  NOR2_X1 U690 ( .A1(G1966), .A2(n729), .ZN(n690) );
  NOR2_X1 U691 ( .A1(n693), .A2(n690), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n623), .A2(G8), .ZN(n624) );
  XOR2_X1 U694 ( .A(n625), .B(n624), .Z(n626) );
  NOR2_X1 U695 ( .A1(G168), .A2(n626), .ZN(n631) );
  INV_X1 U696 ( .A(G1961), .ZN(n986) );
  NAND2_X1 U697 ( .A1(n620), .A2(n986), .ZN(n628) );
  XNOR2_X1 U698 ( .A(G2078), .B(KEYINPUT25), .ZN(n965) );
  NAND2_X1 U699 ( .A1(n669), .A2(n965), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n634) );
  NOR2_X1 U701 ( .A1(G171), .A2(n634), .ZN(n629) );
  XOR2_X1 U702 ( .A(KEYINPUT111), .B(n629), .Z(n630) );
  NOR2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n633), .B(n632), .ZN(n689) );
  AND2_X1 U705 ( .A1(G171), .A2(n634), .ZN(n635) );
  XNOR2_X1 U706 ( .A(KEYINPUT103), .B(n635), .ZN(n687) );
  NAND2_X1 U707 ( .A1(G2072), .A2(n669), .ZN(n637) );
  INV_X1 U708 ( .A(G1956), .ZN(n1007) );
  NOR2_X1 U709 ( .A1(n669), .A2(n1007), .ZN(n638) );
  NOR2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n642) );
  INV_X1 U711 ( .A(G299), .ZN(n988) );
  NOR2_X1 U712 ( .A1(n642), .A2(n988), .ZN(n641) );
  XNOR2_X1 U713 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(n682) );
  NAND2_X1 U715 ( .A1(n642), .A2(n988), .ZN(n680) );
  XNOR2_X1 U716 ( .A(KEYINPUT26), .B(KEYINPUT106), .ZN(n670) );
  NOR2_X1 U717 ( .A1(G1996), .A2(n670), .ZN(n654) );
  XOR2_X1 U718 ( .A(KEYINPUT14), .B(KEYINPUT73), .Z(n644) );
  NAND2_X1 U719 ( .A1(G56), .A2(n813), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n644), .B(n643), .ZN(n653) );
  NAND2_X1 U721 ( .A1(G43), .A2(n814), .ZN(n645) );
  XOR2_X1 U722 ( .A(KEYINPUT74), .B(n645), .Z(n651) );
  NAND2_X1 U723 ( .A1(n817), .A2(G81), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n646), .B(KEYINPUT12), .ZN(n648) );
  NAND2_X1 U725 ( .A1(G68), .A2(n812), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U727 ( .A(KEYINPUT13), .B(n649), .Z(n650) );
  NOR2_X1 U728 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n979) );
  NOR2_X1 U730 ( .A1(n654), .A2(n979), .ZN(n667) );
  NAND2_X1 U731 ( .A1(G92), .A2(n817), .ZN(n655) );
  XNOR2_X1 U732 ( .A(n655), .B(KEYINPUT76), .ZN(n662) );
  NAND2_X1 U733 ( .A1(G66), .A2(n813), .ZN(n657) );
  NAND2_X1 U734 ( .A1(G54), .A2(n814), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U736 ( .A1(G79), .A2(n812), .ZN(n658) );
  XNOR2_X1 U737 ( .A(KEYINPUT77), .B(n658), .ZN(n659) );
  NOR2_X1 U738 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U740 ( .A(KEYINPUT15), .B(n663), .Z(n991) );
  NAND2_X1 U741 ( .A1(G1348), .A2(n620), .ZN(n665) );
  NAND2_X1 U742 ( .A1(G2067), .A2(n669), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n676) );
  NAND2_X1 U744 ( .A1(n991), .A2(n676), .ZN(n666) );
  NAND2_X1 U745 ( .A1(n667), .A2(n666), .ZN(n675) );
  INV_X1 U746 ( .A(G1341), .ZN(n1008) );
  NAND2_X1 U747 ( .A1(n1008), .A2(n670), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n668), .A2(n620), .ZN(n673) );
  AND2_X1 U749 ( .A1(G1996), .A2(n669), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U752 ( .A1(n675), .A2(n674), .ZN(n678) );
  NOR2_X1 U753 ( .A1(n676), .A2(n991), .ZN(n677) );
  NOR2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U755 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U756 ( .A1(n682), .A2(n681), .ZN(n685) );
  XNOR2_X1 U757 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n683) );
  NAND2_X1 U758 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n697) );
  INV_X1 U760 ( .A(n697), .ZN(n691) );
  NOR2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U762 ( .A(n692), .B(KEYINPUT112), .ZN(n695) );
  NAND2_X1 U763 ( .A1(n693), .A2(G8), .ZN(n694) );
  NAND2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n707) );
  AND2_X1 U765 ( .A1(G286), .A2(G8), .ZN(n696) );
  NAND2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n704) );
  INV_X1 U767 ( .A(G8), .ZN(n702) );
  NOR2_X1 U768 ( .A1(G1971), .A2(n729), .ZN(n699) );
  NOR2_X1 U769 ( .A1(G2090), .A2(n620), .ZN(n698) );
  NOR2_X1 U770 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U771 ( .A1(n700), .A2(G303), .ZN(n701) );
  OR2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U774 ( .A(n705), .B(KEYINPUT32), .ZN(n706) );
  NAND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n724) );
  NOR2_X1 U776 ( .A1(G1976), .A2(G288), .ZN(n715) );
  NOR2_X1 U777 ( .A1(G303), .A2(G1971), .ZN(n708) );
  NOR2_X1 U778 ( .A1(n715), .A2(n708), .ZN(n983) );
  NAND2_X1 U779 ( .A1(n724), .A2(n983), .ZN(n711) );
  AND2_X1 U780 ( .A1(G1976), .A2(G288), .ZN(n981) );
  OR2_X1 U781 ( .A1(n981), .A2(n729), .ZN(n709) );
  NOR2_X1 U782 ( .A1(n709), .A2(KEYINPUT113), .ZN(n710) );
  AND2_X1 U783 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U784 ( .A1(KEYINPUT33), .A2(n712), .ZN(n720) );
  INV_X1 U785 ( .A(KEYINPUT113), .ZN(n714) );
  NAND2_X1 U786 ( .A1(n715), .A2(KEYINPUT33), .ZN(n713) );
  NAND2_X1 U787 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U788 ( .A1(n715), .A2(KEYINPUT113), .ZN(n716) );
  NAND2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U790 ( .A1(n729), .A2(n718), .ZN(n719) );
  NOR2_X1 U791 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U792 ( .A(G1981), .B(G305), .Z(n996) );
  NAND2_X1 U793 ( .A1(n721), .A2(n996), .ZN(n733) );
  NOR2_X1 U794 ( .A1(G303), .A2(G2090), .ZN(n722) );
  NAND2_X1 U795 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U796 ( .A(n723), .B(KEYINPUT114), .ZN(n725) );
  NAND2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n726) );
  AND2_X1 U798 ( .A1(n726), .A2(n729), .ZN(n731) );
  NOR2_X1 U799 ( .A1(G1981), .A2(G305), .ZN(n727) );
  XOR2_X1 U800 ( .A(n727), .B(KEYINPUT24), .Z(n728) );
  NOR2_X1 U801 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U802 ( .A1(n731), .A2(n730), .ZN(n732) );
  AND2_X1 U803 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U804 ( .A1(n735), .A2(n734), .ZN(n758) );
  NAND2_X1 U805 ( .A1(G131), .A2(n915), .ZN(n737) );
  NAND2_X1 U806 ( .A1(G95), .A2(n917), .ZN(n736) );
  NAND2_X1 U807 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U808 ( .A(KEYINPUT99), .B(n738), .ZN(n744) );
  NAND2_X1 U809 ( .A1(G119), .A2(n911), .ZN(n739) );
  XNOR2_X1 U810 ( .A(n739), .B(KEYINPUT97), .ZN(n742) );
  NAND2_X1 U811 ( .A1(G107), .A2(n912), .ZN(n740) );
  XOR2_X1 U812 ( .A(KEYINPUT98), .B(n740), .Z(n741) );
  NOR2_X1 U813 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U814 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U815 ( .A(KEYINPUT100), .B(n745), .ZN(n895) );
  AND2_X1 U816 ( .A1(G1991), .A2(n895), .ZN(n755) );
  NAND2_X1 U817 ( .A1(n917), .A2(G105), .ZN(n746) );
  XNOR2_X1 U818 ( .A(n746), .B(KEYINPUT38), .ZN(n753) );
  NAND2_X1 U819 ( .A1(G129), .A2(n911), .ZN(n748) );
  NAND2_X1 U820 ( .A1(G117), .A2(n912), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n751) );
  NAND2_X1 U822 ( .A1(G141), .A2(n915), .ZN(n749) );
  XNOR2_X1 U823 ( .A(KEYINPUT101), .B(n749), .ZN(n750) );
  NOR2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n907) );
  AND2_X1 U826 ( .A1(n907), .A2(G1996), .ZN(n754) );
  NOR2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n939) );
  INV_X1 U828 ( .A(n769), .ZN(n756) );
  NOR2_X1 U829 ( .A1(n939), .A2(n756), .ZN(n762) );
  XOR2_X1 U830 ( .A(KEYINPUT102), .B(n762), .Z(n757) );
  NAND2_X1 U831 ( .A1(n758), .A2(n757), .ZN(n772) );
  NOR2_X1 U832 ( .A1(G1996), .A2(n907), .ZN(n943) );
  NOR2_X1 U833 ( .A1(G1986), .A2(G290), .ZN(n759) );
  XOR2_X1 U834 ( .A(n759), .B(KEYINPUT115), .Z(n760) );
  NOR2_X1 U835 ( .A1(G1991), .A2(n895), .ZN(n938) );
  NOR2_X1 U836 ( .A1(n760), .A2(n938), .ZN(n761) );
  NOR2_X1 U837 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U838 ( .A1(n943), .A2(n763), .ZN(n764) );
  XNOR2_X1 U839 ( .A(KEYINPUT39), .B(n764), .ZN(n766) );
  NAND2_X1 U840 ( .A1(n766), .A2(n765), .ZN(n768) );
  OR2_X1 U841 ( .A1(n767), .A2(n908), .ZN(n947) );
  NAND2_X1 U842 ( .A1(n768), .A2(n947), .ZN(n770) );
  NAND2_X1 U843 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U844 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U845 ( .A(n773), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U846 ( .A(G2443), .B(KEYINPUT118), .Z(n775) );
  XNOR2_X1 U847 ( .A(G2451), .B(G2427), .ZN(n774) );
  XNOR2_X1 U848 ( .A(n775), .B(n774), .ZN(n779) );
  XOR2_X1 U849 ( .A(G2435), .B(G2438), .Z(n777) );
  XNOR2_X1 U850 ( .A(G2454), .B(KEYINPUT117), .ZN(n776) );
  XNOR2_X1 U851 ( .A(n777), .B(n776), .ZN(n778) );
  XOR2_X1 U852 ( .A(n779), .B(n778), .Z(n781) );
  XNOR2_X1 U853 ( .A(G2446), .B(KEYINPUT116), .ZN(n780) );
  XNOR2_X1 U854 ( .A(n781), .B(n780), .ZN(n784) );
  XNOR2_X1 U855 ( .A(G1348), .B(G2430), .ZN(n782) );
  XNOR2_X1 U856 ( .A(n782), .B(n1008), .ZN(n783) );
  XOR2_X1 U857 ( .A(n784), .B(n783), .Z(n785) );
  AND2_X1 U858 ( .A1(G14), .A2(n785), .ZN(G401) );
  AND2_X1 U859 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U860 ( .A1(n911), .A2(G123), .ZN(n786) );
  XNOR2_X1 U861 ( .A(n786), .B(KEYINPUT18), .ZN(n788) );
  NAND2_X1 U862 ( .A1(G111), .A2(n912), .ZN(n787) );
  NAND2_X1 U863 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U864 ( .A1(G135), .A2(n915), .ZN(n790) );
  NAND2_X1 U865 ( .A1(G99), .A2(n917), .ZN(n789) );
  NAND2_X1 U866 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U867 ( .A1(n792), .A2(n791), .ZN(n946) );
  XNOR2_X1 U868 ( .A(n946), .B(G2096), .ZN(n793) );
  XNOR2_X1 U869 ( .A(n793), .B(KEYINPUT81), .ZN(n794) );
  OR2_X1 U870 ( .A1(G2100), .A2(n794), .ZN(G156) );
  INV_X1 U871 ( .A(G120), .ZN(G236) );
  INV_X1 U872 ( .A(G69), .ZN(G235) );
  INV_X1 U873 ( .A(G108), .ZN(G238) );
  INV_X1 U874 ( .A(G132), .ZN(G219) );
  INV_X1 U875 ( .A(G82), .ZN(G220) );
  XOR2_X1 U876 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n796) );
  NAND2_X1 U877 ( .A1(G7), .A2(G661), .ZN(n795) );
  XNOR2_X1 U878 ( .A(n796), .B(n795), .ZN(G223) );
  INV_X1 U879 ( .A(G567), .ZN(n845) );
  NOR2_X1 U880 ( .A1(G223), .A2(n845), .ZN(n798) );
  XNOR2_X1 U881 ( .A(KEYINPUT11), .B(KEYINPUT72), .ZN(n797) );
  XNOR2_X1 U882 ( .A(n798), .B(n797), .ZN(G234) );
  INV_X1 U883 ( .A(G860), .ZN(n859) );
  OR2_X1 U884 ( .A1(n979), .A2(n859), .ZN(G153) );
  XNOR2_X1 U885 ( .A(KEYINPUT75), .B(G171), .ZN(G301) );
  INV_X1 U886 ( .A(G868), .ZN(n830) );
  NAND2_X1 U887 ( .A1(n991), .A2(n830), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n799), .B(KEYINPUT78), .ZN(n801) );
  NAND2_X1 U889 ( .A1(G301), .A2(G868), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n801), .A2(n800), .ZN(G284) );
  NOR2_X1 U891 ( .A1(G286), .A2(n830), .ZN(n803) );
  NOR2_X1 U892 ( .A1(G868), .A2(G299), .ZN(n802) );
  NOR2_X1 U893 ( .A1(n803), .A2(n802), .ZN(G297) );
  NAND2_X1 U894 ( .A1(n859), .A2(G559), .ZN(n804) );
  INV_X1 U895 ( .A(n991), .ZN(n810) );
  NAND2_X1 U896 ( .A1(n804), .A2(n810), .ZN(n805) );
  XNOR2_X1 U897 ( .A(n805), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U898 ( .A1(n991), .A2(n830), .ZN(n806) );
  XOR2_X1 U899 ( .A(KEYINPUT80), .B(n806), .Z(n807) );
  NOR2_X1 U900 ( .A1(G559), .A2(n807), .ZN(n809) );
  NOR2_X1 U901 ( .A1(G868), .A2(n979), .ZN(n808) );
  NOR2_X1 U902 ( .A1(n809), .A2(n808), .ZN(G282) );
  NAND2_X1 U903 ( .A1(G559), .A2(n810), .ZN(n811) );
  XOR2_X1 U904 ( .A(n979), .B(n811), .Z(n858) );
  NAND2_X1 U905 ( .A1(G80), .A2(n812), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G67), .A2(n813), .ZN(n816) );
  NAND2_X1 U907 ( .A1(G55), .A2(n814), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n817), .A2(G93), .ZN(n818) );
  XOR2_X1 U910 ( .A(KEYINPUT82), .B(n818), .Z(n819) );
  NOR2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U912 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U913 ( .A(n823), .B(KEYINPUT83), .Z(n860) );
  XOR2_X1 U914 ( .A(KEYINPUT19), .B(n860), .Z(n825) );
  XNOR2_X1 U915 ( .A(G290), .B(G166), .ZN(n824) );
  XNOR2_X1 U916 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U917 ( .A(n826), .B(G305), .Z(n827) );
  XNOR2_X1 U918 ( .A(G288), .B(n827), .ZN(n828) );
  XNOR2_X1 U919 ( .A(n988), .B(n828), .ZN(n862) );
  XNOR2_X1 U920 ( .A(n858), .B(n862), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n829), .A2(G868), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n830), .A2(n860), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(G295) );
  NAND2_X1 U924 ( .A1(G2084), .A2(G2078), .ZN(n834) );
  XOR2_X1 U925 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n833) );
  XNOR2_X1 U926 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U927 ( .A1(G2090), .A2(n835), .ZN(n836) );
  XNOR2_X1 U928 ( .A(KEYINPUT21), .B(n836), .ZN(n837) );
  NAND2_X1 U929 ( .A1(n837), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U930 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U931 ( .A1(G220), .A2(G219), .ZN(n838) );
  XOR2_X1 U932 ( .A(KEYINPUT22), .B(n838), .Z(n839) );
  NOR2_X1 U933 ( .A1(G218), .A2(n839), .ZN(n840) );
  NAND2_X1 U934 ( .A1(G96), .A2(n840), .ZN(n855) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n855), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n841), .B(KEYINPUT87), .ZN(n847) );
  NOR2_X1 U937 ( .A1(G235), .A2(G236), .ZN(n842) );
  XNOR2_X1 U938 ( .A(KEYINPUT88), .B(n842), .ZN(n843) );
  NAND2_X1 U939 ( .A1(n843), .A2(G57), .ZN(n844) );
  NOR2_X1 U940 ( .A1(G238), .A2(n844), .ZN(n857) );
  NOR2_X1 U941 ( .A1(n845), .A2(n857), .ZN(n846) );
  NOR2_X1 U942 ( .A1(n847), .A2(n846), .ZN(G319) );
  INV_X1 U943 ( .A(G319), .ZN(n928) );
  NAND2_X1 U944 ( .A1(G483), .A2(G661), .ZN(n848) );
  NOR2_X1 U945 ( .A1(n928), .A2(n848), .ZN(n854) );
  NAND2_X1 U946 ( .A1(G36), .A2(n854), .ZN(n849) );
  XOR2_X1 U947 ( .A(KEYINPUT89), .B(n849), .Z(G176) );
  INV_X1 U948 ( .A(G223), .ZN(n850) );
  NAND2_X1 U949 ( .A1(G2106), .A2(n850), .ZN(G217) );
  AND2_X1 U950 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U951 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U952 ( .A1(G3), .A2(G1), .ZN(n852) );
  XOR2_X1 U953 ( .A(KEYINPUT119), .B(n852), .Z(n853) );
  NAND2_X1 U954 ( .A1(n854), .A2(n853), .ZN(G188) );
  INV_X1 U956 ( .A(G96), .ZN(G221) );
  INV_X1 U957 ( .A(G57), .ZN(G237) );
  INV_X1 U958 ( .A(n855), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(G261) );
  INV_X1 U960 ( .A(G261), .ZN(G325) );
  NAND2_X1 U961 ( .A1(n859), .A2(n858), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(G145) );
  XNOR2_X1 U963 ( .A(n862), .B(n991), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n863), .B(n979), .ZN(n865) );
  INV_X1 U965 ( .A(G171), .ZN(n987) );
  XNOR2_X1 U966 ( .A(G286), .B(n987), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n866) );
  NOR2_X1 U968 ( .A1(G37), .A2(n866), .ZN(G397) );
  XOR2_X1 U969 ( .A(KEYINPUT120), .B(G1981), .Z(n868) );
  XNOR2_X1 U970 ( .A(G1966), .B(G1956), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U972 ( .A(n869), .B(KEYINPUT41), .Z(n871) );
  XNOR2_X1 U973 ( .A(G1996), .B(G1991), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U975 ( .A(G1976), .B(G1971), .Z(n873) );
  XNOR2_X1 U976 ( .A(G1986), .B(G1961), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U978 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U979 ( .A(KEYINPUT121), .B(G2474), .ZN(n876) );
  XNOR2_X1 U980 ( .A(n877), .B(n876), .ZN(G229) );
  XOR2_X1 U981 ( .A(G2100), .B(G2096), .Z(n879) );
  XNOR2_X1 U982 ( .A(KEYINPUT42), .B(G2678), .ZN(n878) );
  XNOR2_X1 U983 ( .A(n879), .B(n878), .ZN(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT43), .B(G2090), .Z(n881) );
  XNOR2_X1 U985 ( .A(G2067), .B(G2072), .ZN(n880) );
  XNOR2_X1 U986 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U987 ( .A(n883), .B(n882), .Z(n885) );
  XNOR2_X1 U988 ( .A(G2084), .B(G2078), .ZN(n884) );
  XNOR2_X1 U989 ( .A(n885), .B(n884), .ZN(G227) );
  NAND2_X1 U990 ( .A1(n911), .A2(G124), .ZN(n886) );
  XNOR2_X1 U991 ( .A(n886), .B(KEYINPUT44), .ZN(n888) );
  NAND2_X1 U992 ( .A1(G112), .A2(n912), .ZN(n887) );
  NAND2_X1 U993 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U994 ( .A1(G136), .A2(n915), .ZN(n890) );
  NAND2_X1 U995 ( .A1(G100), .A2(n917), .ZN(n889) );
  NAND2_X1 U996 ( .A1(n890), .A2(n889), .ZN(n891) );
  NOR2_X1 U997 ( .A1(n892), .A2(n891), .ZN(G162) );
  XOR2_X1 U998 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n894) );
  XNOR2_X1 U999 ( .A(G162), .B(n946), .ZN(n893) );
  XNOR2_X1 U1000 ( .A(n894), .B(n893), .ZN(n896) );
  XOR2_X1 U1001 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U1002 ( .A(G164), .B(G160), .ZN(n897) );
  XNOR2_X1 U1003 ( .A(n898), .B(n897), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(G139), .A2(n915), .ZN(n900) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n917), .ZN(n899) );
  NAND2_X1 U1006 ( .A1(n900), .A2(n899), .ZN(n905) );
  NAND2_X1 U1007 ( .A1(G127), .A2(n911), .ZN(n902) );
  NAND2_X1 U1008 ( .A1(G115), .A2(n912), .ZN(n901) );
  NAND2_X1 U1009 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1010 ( .A(KEYINPUT47), .B(n903), .Z(n904) );
  NOR2_X1 U1011 ( .A1(n905), .A2(n904), .ZN(n933) );
  XOR2_X1 U1012 ( .A(n906), .B(n933), .Z(n910) );
  XOR2_X1 U1013 ( .A(n908), .B(n907), .Z(n909) );
  XNOR2_X1 U1014 ( .A(n910), .B(n909), .ZN(n924) );
  NAND2_X1 U1015 ( .A1(G130), .A2(n911), .ZN(n914) );
  NAND2_X1 U1016 ( .A1(G118), .A2(n912), .ZN(n913) );
  NAND2_X1 U1017 ( .A1(n914), .A2(n913), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n915), .A2(G142), .ZN(n916) );
  XNOR2_X1 U1019 ( .A(n916), .B(KEYINPUT122), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(G106), .A2(n917), .ZN(n918) );
  NAND2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1022 ( .A(n920), .B(KEYINPUT45), .Z(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1024 ( .A(n924), .B(n923), .Z(n925) );
  NOR2_X1 U1025 ( .A1(G37), .A2(n925), .ZN(G395) );
  NOR2_X1 U1026 ( .A1(G229), .A2(G227), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(KEYINPUT49), .B(n926), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(G397), .A2(n927), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(G401), .A2(n928), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT123), .B(n929), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(G395), .A2(n930), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(G225) );
  INV_X1 U1033 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1034 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n936), .Z(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n952) );
  XNOR2_X1 U1039 ( .A(G160), .B(G2084), .ZN(n940) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n950) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n941) );
  XNOR2_X1 U1042 ( .A(KEYINPUT124), .B(n941), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT51), .B(n944), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT52), .B(n955), .ZN(n956) );
  INV_X1 U1051 ( .A(KEYINPUT55), .ZN(n975) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n975), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n957), .A2(G29), .ZN(n1037) );
  XNOR2_X1 U1054 ( .A(G2090), .B(G35), .ZN(n970) );
  XNOR2_X1 U1055 ( .A(G1996), .B(G32), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(G33), .B(G2072), .ZN(n958) );
  NOR2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n964) );
  XOR2_X1 U1058 ( .A(G25), .B(G1991), .Z(n960) );
  NAND2_X1 U1059 ( .A1(n960), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(G26), .B(G2067), .ZN(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1063 ( .A(G27), .B(n965), .Z(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n968), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1067 ( .A(G2084), .B(G34), .Z(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT54), .B(n971), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n975), .B(n974), .ZN(n977) );
  INV_X1 U1071 ( .A(G29), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n978), .ZN(n1035) );
  XNOR2_X1 U1074 ( .A(G16), .B(KEYINPUT56), .ZN(n1005) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n979), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n1003) );
  XNOR2_X1 U1079 ( .A(n987), .B(n986), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(n988), .B(G1956), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(G1971), .A2(G303), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(G1348), .B(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G168), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n998), .B(KEYINPUT125), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n999), .B(KEYINPUT57), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1033) );
  INV_X1 U1093 ( .A(G16), .ZN(n1031) );
  XNOR2_X1 U1094 ( .A(KEYINPUT127), .B(G1966), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1006), .B(G21), .ZN(n1026) );
  XNOR2_X1 U1096 ( .A(n1007), .B(G20), .ZN(n1016) );
  XNOR2_X1 U1097 ( .A(n1008), .B(G19), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(G1981), .B(G6), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT126), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(KEYINPUT59), .B(G1348), .Z(n1012) );
  XNOR2_X1 U1102 ( .A(G4), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(n1017), .B(KEYINPUT60), .ZN(n1024) );
  XNOR2_X1 U1106 ( .A(G1986), .B(G24), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(G1971), .B(G22), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XOR2_X1 U1109 ( .A(G1976), .B(G23), .Z(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(G5), .B(G1961), .ZN(n1027) );
  NOR2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(KEYINPUT61), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1120 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1038), .Z(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

