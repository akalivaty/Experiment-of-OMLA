//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT79), .B1(new_n191), .B2(G104), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(new_n188), .A3(G107), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n189), .A2(new_n194), .A3(new_n192), .A4(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G101), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT4), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n204), .A3(G101), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n199), .A2(new_n201), .A3(KEYINPUT80), .A4(KEYINPUT4), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT65), .B1(new_n211), .B2(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n210), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT0), .A3(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(KEYINPUT69), .A3(new_n221), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n206), .A2(new_n207), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n191), .A2(KEYINPUT81), .A3(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n188), .A2(G107), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT81), .B1(new_n191), .B2(G104), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(G101), .B2(new_n200), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT82), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n214), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n216), .A2(new_n234), .A3(new_n235), .A4(G128), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n220), .A2(new_n238), .A3(new_n235), .A4(G128), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G128), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n217), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n199), .A2(new_n245), .A3(new_n231), .ZN(new_n246));
  AND4_X1   g060(.A1(KEYINPUT10), .A2(new_n233), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n232), .ZN(new_n248));
  INV_X1    g062(.A(new_n220), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n240), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT10), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n226), .A2(new_n247), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G137), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(G137), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n253), .A2(KEYINPUT83), .A3(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n199), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n205), .A2(new_n203), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n207), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n224), .A2(new_n225), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n252), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n246), .A4(new_n244), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n262), .A4(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT83), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n262), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n263), .A2(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(G110), .B(G140), .Z(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT78), .ZN(new_n278));
  INV_X1    g092(.A(G227), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G953), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n278), .B(new_n280), .Z(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n187), .B1(new_n276), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n275), .A2(new_n274), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT83), .B1(new_n253), .B2(new_n262), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n271), .A2(new_n272), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT84), .A3(new_n281), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n281), .B1(new_n263), .B2(new_n273), .ZN(new_n289));
  INV_X1    g103(.A(new_n251), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(new_n232), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n248), .A2(new_n244), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n274), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n293), .B(KEYINPUT12), .Z(new_n294));
  NAND2_X1  g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n283), .A2(new_n288), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G469), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n294), .B1(new_n285), .B2(new_n286), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n300), .A2(new_n281), .B1(new_n289), .B2(new_n284), .ZN(new_n301));
  OAI21_X1  g115(.A(G469), .B1(new_n301), .B2(G902), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT9), .B(G234), .Z(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G221), .B1(new_n305), .B2(G902), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT77), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G237), .ZN(new_n309));
  INV_X1    g123(.A(G953), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G214), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n211), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n309), .A2(new_n310), .A3(G143), .A4(G214), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT18), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(new_n261), .ZN(new_n316));
  OR2_X1    g130(.A1(G125), .A2(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(G125), .A2(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(new_n214), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n312), .A2(new_n313), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT18), .A3(G131), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n316), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n317), .B2(new_n318), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n327), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n326), .A2(new_n214), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT93), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n319), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT19), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n319), .B2(new_n330), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n336), .B2(new_n332), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n329), .B1(new_n337), .B2(new_n214), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT92), .B1(new_n314), .B2(new_n261), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT92), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n321), .A2(new_n340), .A3(G131), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n314), .A2(new_n261), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n324), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G113), .B(G122), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n188), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT95), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT95), .ZN(new_n349));
  INV_X1    g163(.A(new_n347), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n339), .A2(new_n341), .B1(new_n261), .B2(new_n314), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n317), .A2(new_n318), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT93), .B1(new_n352), .B2(KEYINPUT94), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n335), .ZN(new_n354));
  AOI21_X1  g168(.A(G146), .B1(new_n354), .B2(new_n334), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n351), .A2(new_n355), .A3(new_n329), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n349), .B(new_n350), .C1(new_n356), .C2(new_n324), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT96), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT17), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n342), .A2(new_n358), .A3(new_n359), .A4(new_n343), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n340), .B1(new_n321), .B2(G131), .ZN(new_n361));
  AOI211_X1 g175(.A(KEYINPUT92), .B(new_n261), .C1(new_n312), .C2(new_n313), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n359), .B(new_n343), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT96), .ZN(new_n364));
  OR3_X1    g178(.A1(new_n326), .A2(new_n214), .A3(new_n328), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n214), .B1(new_n326), .B2(new_n328), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n361), .A2(new_n362), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(KEYINPUT17), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n347), .A3(new_n323), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n348), .A2(new_n357), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G475), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n298), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n372), .A2(KEYINPUT97), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(KEYINPUT20), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT20), .B1(new_n372), .B2(KEYINPUT97), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(new_n373), .A3(new_n298), .A4(new_n372), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G128), .B(G143), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n255), .ZN(new_n381));
  INV_X1    g195(.A(G116), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT14), .A3(G122), .ZN(new_n383));
  XNOR2_X1  g197(.A(G116), .B(G122), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(G107), .B(new_n383), .C1(new_n385), .C2(KEYINPUT14), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n381), .B(new_n386), .C1(G107), .C2(new_n385), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT99), .B(KEYINPUT13), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n380), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n211), .A2(G128), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n389), .B(G134), .C1(new_n390), .C2(new_n388), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n384), .B(new_n191), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n380), .A2(new_n255), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n304), .A2(G217), .A3(new_n310), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n298), .ZN(new_n398));
  INV_X1    g212(.A(G478), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(KEYINPUT15), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n398), .B(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT98), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n370), .A2(new_n323), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n350), .ZN(new_n404));
  AOI211_X1 g218(.A(KEYINPUT98), .B(new_n347), .C1(new_n370), .C2(new_n323), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n371), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n298), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n401), .B1(new_n407), .B2(G475), .ZN(new_n408));
  NAND2_X1  g222(.A1(G234), .A2(G237), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(G952), .A3(new_n310), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT21), .B(G898), .Z(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(G902), .A3(G953), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n379), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n308), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT67), .B(G119), .ZN(new_n416));
  INV_X1    g230(.A(G128), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT23), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G119), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(G128), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n416), .B2(new_n417), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n418), .B1(KEYINPUT23), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G110), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT72), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(KEYINPUT67), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT67), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G119), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n420), .B1(new_n429), .B2(G128), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT24), .B(G110), .Z(new_n431));
  AOI22_X1  g245(.A1(new_n365), .A2(new_n366), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT23), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n429), .B2(G128), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n430), .B2(new_n433), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT72), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(G110), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n425), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  OAI22_X1  g252(.A1(new_n435), .A2(G110), .B1(new_n430), .B2(new_n431), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n329), .B1(new_n214), .B2(new_n319), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n310), .A2(G221), .A3(G234), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT22), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(new_n258), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT22), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n442), .B(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(G137), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n438), .A2(new_n441), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT73), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n444), .B2(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(G137), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n443), .A2(new_n258), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT73), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n438), .B2(new_n441), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT76), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G217), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(G234), .B2(new_n298), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G902), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n438), .A2(new_n441), .ZN(new_n464));
  INV_X1    g278(.A(new_n455), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n438), .A2(new_n441), .A3(new_n448), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT74), .B(KEYINPUT25), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(new_n298), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n449), .A2(new_n456), .A3(G902), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(KEYINPUT74), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n461), .B(new_n469), .C1(new_n470), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT75), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n466), .A2(new_n298), .A3(new_n467), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n472), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(KEYINPUT75), .A3(new_n461), .A4(new_n469), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n463), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n237), .A2(new_n239), .B1(new_n242), .B2(new_n217), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n260), .A2(G131), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n258), .A2(G134), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n261), .B1(new_n257), .B2(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n262), .A2(new_n222), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT2), .B(G113), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n427), .A2(G119), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n419), .A2(KEYINPUT67), .ZN(new_n492));
  OAI21_X1  g306(.A(G116), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n419), .A2(G116), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n490), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n382), .B1(new_n426), .B2(new_n428), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n497), .A2(new_n489), .A3(new_n494), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n488), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n490), .A3(new_n495), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n489), .B1(new_n497), .B2(new_n494), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT68), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n487), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT28), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n485), .B1(new_n267), .B2(new_n274), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n507), .B2(new_n503), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n219), .A2(KEYINPUT69), .A3(new_n221), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT69), .B1(new_n219), .B2(new_n221), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n274), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n484), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n244), .B(new_n512), .C1(G131), .C2(new_n260), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n511), .A2(new_n513), .A3(new_n506), .A4(new_n503), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n505), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT70), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(G101), .ZN(new_n519));
  INV_X1    g333(.A(G210), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n520), .A2(G237), .A3(G953), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n519), .B(new_n521), .Z(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n516), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n511), .A2(new_n503), .A3(new_n513), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT28), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n504), .B1(new_n526), .B2(new_n514), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT70), .B1(new_n527), .B2(new_n522), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n511), .A2(KEYINPUT30), .A3(new_n513), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n485), .B2(new_n486), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n499), .A2(new_n502), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n525), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT31), .B1(new_n534), .B2(new_n523), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT31), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n533), .A2(new_n536), .A3(new_n525), .A4(new_n522), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n524), .A2(new_n528), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G472), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n298), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT32), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT32), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n538), .A2(new_n542), .A3(new_n539), .A4(new_n298), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n507), .A2(new_n503), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n526), .B2(new_n514), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n523), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(G902), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n523), .B1(new_n527), .B2(KEYINPUT71), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n522), .B1(new_n507), .B2(new_n503), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n551), .A2(new_n533), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n547), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT71), .B1(new_n527), .B2(new_n522), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G472), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n480), .B1(new_n544), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G214), .B1(G237), .B2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n327), .B1(new_n219), .B2(new_n221), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT89), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n481), .A2(new_n327), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G224), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G953), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n563), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(G110), .B(G122), .Z(new_n567));
  AOI21_X1  g381(.A(new_n503), .B1(new_n206), .B2(new_n207), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n569));
  OR3_X1    g383(.A1(new_n497), .A2(new_n494), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G113), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n497), .B2(new_n569), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n498), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n233), .A3(new_n246), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n567), .B1(new_n568), .B2(new_n575), .ZN(new_n576));
  OR3_X1    g390(.A1(new_n576), .A2(KEYINPUT88), .A3(KEYINPUT6), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT88), .B1(new_n576), .B2(KEYINPUT6), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n568), .A2(new_n575), .A3(new_n567), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(KEYINPUT86), .B2(new_n576), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT6), .ZN(new_n582));
  INV_X1    g396(.A(new_n567), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n266), .A2(new_n532), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(new_n574), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT86), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT87), .B1(new_n581), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(new_n574), .A3(new_n583), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n585), .B2(new_n586), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n586), .B(new_n567), .C1(new_n568), .C2(new_n575), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT6), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT87), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n566), .B(new_n579), .C1(new_n588), .C2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT7), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n563), .B1(new_n596), .B2(new_n565), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT90), .B(KEYINPUT8), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n567), .B(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n493), .A2(KEYINPUT5), .A3(new_n495), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n498), .B(new_n232), .C1(new_n572), .C2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n573), .A2(new_n248), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n565), .A2(new_n596), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n561), .A2(new_n604), .A3(new_n562), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n597), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n580), .B1(new_n606), .B2(KEYINPUT91), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(KEYINPUT91), .B2(new_n606), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n595), .A2(new_n298), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G210), .B1(G237), .B2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n595), .A2(new_n298), .A3(new_n610), .A4(new_n608), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n559), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n415), .A2(new_n557), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  AOI22_X1  g430(.A1(new_n376), .A2(new_n378), .B1(new_n407), .B2(G475), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n397), .B(KEYINPUT33), .Z(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G478), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n397), .A2(new_n399), .A3(new_n298), .ZN(new_n620));
  NAND2_X1  g434(.A1(G478), .A2(G902), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n614), .A2(new_n413), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n538), .A2(new_n298), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(G472), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(new_n540), .ZN(new_n627));
  INV_X1    g441(.A(new_n307), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n628), .B(new_n480), .C1(new_n299), .C2(new_n302), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n624), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(new_n401), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n407), .B2(G475), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n374), .B(KEYINPUT20), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n614), .A2(new_n413), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n627), .ZN(new_n637));
  NOR4_X1   g451(.A1(new_n636), .A2(new_n308), .A3(new_n480), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT35), .B(G107), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n465), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n464), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n462), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n476), .A2(new_n479), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT100), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n476), .A2(new_n479), .A3(new_n646), .A4(new_n643), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  AOI211_X1 g462(.A(new_n559), .B(new_n648), .C1(new_n612), .C2(new_n613), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n415), .A3(new_n627), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT37), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n424), .ZN(G12));
  AOI22_X1  g466(.A1(new_n541), .A2(new_n543), .B1(G472), .B2(new_n555), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n308), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n410), .B1(new_n412), .B2(G900), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n635), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n656), .A2(new_n634), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n649), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  NAND2_X1  g473(.A1(new_n612), .A2(new_n613), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT38), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n534), .A2(new_n522), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n551), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n298), .B1(new_n664), .B2(new_n545), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n544), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n655), .B(KEYINPUT39), .Z(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n303), .A2(new_n307), .A3(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n617), .A2(new_n633), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n558), .B(new_n673), .C1(new_n671), .C2(KEYINPUT40), .ZN(new_n674));
  INV_X1    g488(.A(new_n648), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n668), .A2(new_n672), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT101), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n211), .ZN(G45));
  AND2_X1   g492(.A1(new_n623), .A2(new_n655), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n649), .A2(new_n654), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  NAND2_X1  g495(.A1(new_n544), .A2(new_n556), .ZN(new_n682));
  INV_X1    g496(.A(new_n480), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n296), .A2(new_n298), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n306), .A3(new_n299), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n624), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  AND3_X1   g505(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n693));
  INV_X1    g507(.A(new_n306), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n557), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n636), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  AOI21_X1  g512(.A(new_n414), .B1(new_n544), .B2(new_n556), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n695), .A2(new_n614), .A3(new_n699), .A4(new_n675), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  OAI21_X1  g515(.A(KEYINPUT103), .B1(new_n617), .B2(new_n633), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n593), .B1(new_n590), .B2(new_n592), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n576), .A2(KEYINPUT86), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n587), .A2(KEYINPUT87), .A3(new_n589), .A4(new_n704), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n703), .A2(new_n705), .B1(new_n578), .B2(new_n577), .ZN(new_n706));
  AOI21_X1  g520(.A(G902), .B1(new_n706), .B2(new_n566), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n610), .B1(new_n707), .B2(new_n608), .ZN(new_n708));
  INV_X1    g522(.A(new_n613), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n702), .B(new_n558), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n686), .A2(new_n306), .A3(new_n299), .A4(new_n413), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT102), .B(G472), .Z(new_n714));
  NAND2_X1  g528(.A1(new_n625), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n535), .A2(new_n537), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n546), .A2(new_n522), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n539), .B(new_n298), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n480), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n617), .A2(KEYINPUT103), .A3(new_n633), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n711), .A2(new_n713), .A3(new_n720), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  AND2_X1   g538(.A1(new_n715), .A2(new_n718), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n675), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT104), .B1(new_n648), .B2(new_n719), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n614), .A3(new_n679), .A4(new_n695), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT105), .B(G125), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G27));
  NAND3_X1  g546(.A1(new_n612), .A2(new_n558), .A3(new_n613), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n733), .A2(new_n480), .A3(new_n653), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n694), .B1(new_n299), .B2(new_n302), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n736));
  NAND4_X1  g550(.A1(new_n734), .A2(new_n679), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n612), .A2(new_n558), .A3(new_n613), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n679), .A3(new_n557), .A4(new_n735), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT42), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  NAND3_X1  g558(.A1(new_n734), .A2(new_n657), .A3(new_n735), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  INV_X1    g560(.A(new_n622), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n617), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT108), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT43), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n750), .A2(KEYINPUT109), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n648), .B1(new_n750), .B2(KEYINPUT109), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n637), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n733), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n300), .A2(new_n281), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n289), .A2(new_n284), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n301), .A2(KEYINPUT45), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(G469), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(G469), .A2(G902), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT107), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n767), .A3(KEYINPUT46), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n765), .A2(new_n766), .A3(new_n299), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n306), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n669), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n751), .A2(new_n752), .A3(KEYINPUT44), .A4(new_n637), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n755), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  AND2_X1   g588(.A1(new_n679), .A2(new_n480), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n733), .A2(new_n682), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n769), .A2(KEYINPUT47), .A3(new_n306), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT47), .B1(new_n769), .B2(new_n306), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n775), .B(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  INV_X1    g594(.A(G952), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n310), .ZN(new_n782));
  INV_X1    g596(.A(new_n644), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n735), .A2(new_n667), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n711), .A3(new_n655), .A4(new_n722), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n649), .B(new_n654), .C1(new_n657), .C2(new_n679), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n786), .A3(new_n730), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n785), .A2(new_n786), .A3(new_n730), .A4(KEYINPUT52), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n710), .A2(new_n712), .A3(new_n721), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n791), .A2(new_n720), .B1(new_n624), .B2(new_n688), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n700), .B1(new_n636), .B2(new_n696), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n743), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n789), .A2(new_n790), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n743), .A2(new_n792), .A3(new_n794), .A4(KEYINPUT112), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n729), .A2(new_n679), .A3(new_n735), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n675), .A2(new_n408), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n654), .A2(new_n656), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n738), .ZN(new_n804));
  INV_X1    g618(.A(new_n413), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n805), .B(new_n559), .C1(new_n612), .C2(new_n613), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n617), .A2(new_n401), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n617), .B2(new_n622), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n806), .A2(new_n629), .A3(new_n627), .A4(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n650), .A2(new_n615), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n804), .A2(new_n810), .A3(new_n745), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT111), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n804), .A2(new_n810), .A3(new_n813), .A4(new_n745), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n797), .A2(new_n799), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n789), .A2(new_n790), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n733), .B1(new_n800), .B2(new_n802), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n650), .A2(new_n615), .A3(new_n809), .ZN(new_n819));
  INV_X1    g633(.A(new_n745), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n795), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n815), .A2(new_n816), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT110), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n789), .B2(new_n790), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n823), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n795), .B1(new_n789), .B2(new_n790), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n831), .B(new_n821), .C1(new_n828), .C2(KEYINPUT53), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n816), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n826), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n410), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n750), .A2(new_n835), .A3(new_n720), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n614), .A3(new_n695), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n660), .B(KEYINPUT38), .Z(new_n838));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n687), .B2(new_n558), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n695), .A2(KEYINPUT115), .A3(new_n559), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n841), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT116), .B1(new_n844), .B2(new_n661), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n845), .A3(new_n836), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT50), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT50), .A4(new_n836), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n687), .A2(new_n733), .A3(new_n410), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n667), .A2(new_n480), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n617), .A3(new_n622), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n750), .A2(new_n851), .A3(new_n729), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n836), .A2(new_n738), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n777), .A2(new_n778), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n692), .A2(new_n693), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT113), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n628), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT114), .Z(new_n864));
  OAI21_X1  g678(.A(new_n859), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n850), .A2(KEYINPUT117), .A3(new_n855), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n858), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n834), .B(new_n837), .C1(KEYINPUT51), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n863), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n859), .B1(new_n860), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n855), .B2(KEYINPUT118), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n855), .A2(KEYINPUT118), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(new_n872), .A3(new_n850), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n851), .A2(new_n623), .A3(new_n852), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT48), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n750), .A2(new_n851), .ZN(new_n877));
  OAI211_X1 g691(.A(KEYINPUT119), .B(new_n876), .C1(new_n877), .C2(new_n684), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n684), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT119), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n781), .B(G953), .C1(new_n880), .C2(KEYINPUT48), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n874), .A2(new_n875), .A3(new_n878), .A4(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n782), .B1(new_n868), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT49), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n748), .B1(new_n861), .B2(new_n884), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n558), .A2(new_n838), .A3(new_n852), .A4(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n886), .B(new_n307), .C1(new_n884), .C2(new_n861), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n887), .ZN(G75));
  XOR2_X1   g702(.A(new_n706), .B(new_n566), .Z(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n298), .B1(new_n815), .B2(new_n825), .ZN(new_n893));
  AOI211_X1 g707(.A(KEYINPUT55), .B(new_n892), .C1(new_n893), .C2(G210), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT55), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n795), .A2(new_n796), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n817), .A2(new_n896), .A3(KEYINPUT53), .A4(new_n798), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n812), .A2(new_n814), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT53), .B1(new_n831), .B2(new_n821), .ZN(new_n900));
  OAI211_X1 g714(.A(G210), .B(G902), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n895), .B1(new_n901), .B2(new_n891), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n890), .B1(new_n894), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n310), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n520), .B(new_n298), .C1(new_n815), .C2(new_n825), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT55), .B1(new_n906), .B2(new_n892), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n901), .A2(new_n895), .A3(new_n891), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n908), .A3(new_n889), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n903), .A2(new_n905), .A3(new_n909), .ZN(G51));
  AOI211_X1 g724(.A(new_n298), .B(new_n761), .C1(new_n815), .C2(new_n825), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n762), .B(KEYINPUT57), .Z(new_n912));
  AOI21_X1  g726(.A(new_n816), .B1(new_n815), .B2(new_n825), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n826), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n914), .B2(new_n296), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT121), .B1(new_n915), .B2(new_n904), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n917));
  INV_X1    g731(.A(new_n296), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT54), .B1(new_n899), .B2(new_n900), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n815), .A2(new_n816), .A3(new_n825), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n921), .B2(new_n912), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n917), .B(new_n905), .C1(new_n922), .C2(new_n911), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n916), .A2(new_n923), .ZN(G54));
  AND3_X1   g738(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(new_n372), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n372), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n904), .ZN(G60));
  INV_X1    g742(.A(new_n618), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n621), .B(KEYINPUT59), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n921), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT122), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n826), .B2(new_n833), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n904), .B1(new_n933), .B2(new_n618), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n921), .A2(new_n935), .A3(new_n929), .A4(new_n930), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n932), .A2(new_n934), .A3(new_n936), .ZN(G63));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n815), .B2(new_n825), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n642), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n905), .B1(new_n941), .B2(new_n459), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n938), .B(KEYINPUT61), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n942), .B(new_n905), .C1(new_n459), .C2(new_n941), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT61), .B1(new_n947), .B2(new_n938), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n411), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n950), .B2(new_n564), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n792), .A2(new_n794), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(new_n819), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n953), .B2(G953), .ZN(new_n954));
  INV_X1    g768(.A(new_n706), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(G898), .B2(new_n310), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  NAND2_X1  g771(.A1(new_n529), .A2(new_n531), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n337), .ZN(new_n959));
  INV_X1    g773(.A(G900), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n279), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n773), .A2(new_n779), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n786), .A2(new_n730), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n676), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n808), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n671), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n808), .A2(new_n967), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n734), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n963), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n962), .B1(new_n972), .B2(new_n310), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n711), .A2(new_n722), .ZN(new_n974));
  NOR4_X1   g788(.A1(new_n770), .A2(new_n684), .A3(new_n669), .A4(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n743), .A2(new_n730), .A3(new_n786), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n963), .A2(new_n745), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n959), .B1(new_n979), .B2(new_n310), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n960), .B2(G227), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n973), .B1(new_n980), .B2(new_n981), .ZN(G72));
  XOR2_X1   g796(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n983));
  NOR2_X1   g797(.A1(new_n539), .A2(new_n298), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT126), .ZN(new_n986));
  INV_X1    g800(.A(new_n953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n978), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n904), .B1(new_n988), .B2(new_n552), .ZN(new_n989));
  AOI211_X1 g803(.A(new_n663), .B(new_n985), .C1(new_n830), .C2(new_n832), .ZN(new_n990));
  INV_X1    g804(.A(new_n552), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n963), .A2(new_n966), .A3(new_n953), .A4(new_n971), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n986), .ZN(new_n994));
  AOI21_X1  g808(.A(KEYINPUT127), .B1(new_n994), .B2(new_n663), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n996), .B(new_n662), .C1(new_n993), .C2(new_n986), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n989), .B(new_n992), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(G57));
endmodule


