//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1100,
    new_n1101, new_n1102, new_n1103;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  NOR3_X1   g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n461), .B2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n465), .A2(new_n469), .B1(new_n474), .B2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n460), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n466), .A2(new_n467), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(G160));
  INV_X1    g060(.A(new_n465), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(new_n481), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT72), .Z(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n481), .C2(G112), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n486), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT71), .Z(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(G138), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n476), .A2(new_n477), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n498), .A2(KEYINPUT4), .A3(G138), .A4(new_n499), .ZN(new_n509));
  NAND2_X1  g084(.A1(G126), .A2(G2105), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n509), .A2(new_n510), .B1(new_n462), .B2(new_n464), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n516), .A2(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT73), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n522), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n521), .A2(new_n526), .ZN(G166));
  XOR2_X1   g102(.A(KEYINPUT5), .B(G543), .Z(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT74), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n529), .A2(G63), .A3(G651), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(new_n519), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n517), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT75), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n532), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n529), .A2(G64), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n522), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n517), .A2(new_n542), .B1(new_n519), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n522), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n517), .A2(new_n548), .B1(new_n519), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G188));
  INV_X1    g133(.A(new_n519), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n528), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n515), .A2(new_n516), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(G651), .B1(new_n565), .B2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  OAI21_X1  g145(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n565), .A2(KEYINPUT77), .A3(G87), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n517), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n572), .A2(new_n575), .B1(G49), .B2(new_n559), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n571), .A2(new_n576), .ZN(G288));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n517), .A2(new_n578), .B1(new_n519), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n522), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(G47), .A2(new_n559), .B1(new_n565), .B2(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n522), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n565), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT78), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n528), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n559), .B2(G54), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n589), .B1(new_n600), .B2(new_n588), .ZN(G284));
  AOI21_X1  g176(.A(new_n589), .B1(new_n600), .B2(new_n588), .ZN(G321));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT80), .B1(new_n603), .B2(G868), .ZN(new_n604));
  NOR2_X1   g179(.A1(G168), .A2(new_n588), .ZN(new_n605));
  MUX2_X1   g180(.A(new_n604), .B(KEYINPUT80), .S(new_n605), .Z(G297));
  MUX2_X1   g181(.A(new_n604), .B(KEYINPUT80), .S(new_n605), .Z(G280));
  XOR2_X1   g182(.A(KEYINPUT81), .B(G559), .Z(new_n608));
  OAI21_X1  g183(.A(new_n600), .B1(G860), .B2(new_n608), .ZN(G148));
  NAND2_X1  g184(.A1(new_n600), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(KEYINPUT82), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(KEYINPUT82), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n612), .B(new_n613), .C1(G868), .C2(new_n551), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n487), .A2(G123), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n492), .A2(G135), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n620), .B(new_n621), .C1(G111), .C2(new_n481), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n616), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  INV_X1    g199(.A(new_n501), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n474), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT13), .Z(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT85), .Z(G156));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT89), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT88), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n637), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT87), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n645), .A2(new_n649), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT90), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT17), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n655), .B2(new_n657), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n656), .B2(new_n657), .ZN(new_n661));
  INV_X1    g236(.A(new_n657), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(new_n658), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n659), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n630), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT91), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT93), .ZN(new_n680));
  OR3_X1    g255(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G288), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n692), .B2(G23), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT33), .B(G1976), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n692), .A2(G22), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n692), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(G1971), .Z(new_n700));
  NOR2_X1   g275(.A1(G6), .A2(G16), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n583), .B2(G16), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT32), .B(G1981), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n696), .A2(new_n697), .A3(new_n700), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT34), .Z(new_n706));
  XNOR2_X1  g281(.A(G290), .B(KEYINPUT94), .ZN(new_n707));
  MUX2_X1   g282(.A(G24), .B(new_n707), .S(G16), .Z(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT95), .B(G1986), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n487), .A2(G119), .ZN(new_n713));
  OAI221_X1 g288(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n481), .C2(G107), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n492), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n718), .B2(new_n711), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  XOR2_X1   g295(.A(new_n719), .B(new_n720), .Z(new_n721));
  NOR3_X1   g296(.A1(new_n710), .A2(KEYINPUT96), .A3(new_n721), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n706), .B(new_n722), .C1(new_n708), .C2(new_n709), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n711), .A2(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n711), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G2090), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT102), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n692), .A2(G5), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G171), .B2(new_n692), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1961), .ZN(new_n734));
  INV_X1    g309(.A(G34), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(KEYINPUT24), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(KEYINPUT24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n711), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G160), .B2(new_n711), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2084), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n692), .A2(G20), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT23), .Z(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G299), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT103), .ZN(new_n745));
  INV_X1    g320(.A(G1956), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n741), .B(new_n747), .C1(new_n729), .C2(G2090), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT25), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n492), .A2(G139), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n625), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n750), .B(new_n751), .C1(new_n481), .C2(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G33), .B(new_n753), .S(G29), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2072), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n711), .A2(G32), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n492), .A2(G141), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n487), .A2(G129), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT26), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n474), .A2(G105), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n757), .A2(new_n758), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n756), .B1(new_n763), .B2(new_n711), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT27), .B(G1996), .Z(new_n765));
  AOI21_X1  g340(.A(new_n755), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n711), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  OAI221_X1 g343(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n481), .C2(G116), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT98), .ZN(new_n770));
  AOI22_X1  g345(.A1(G128), .A2(new_n487), .B1(new_n492), .B2(G140), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n768), .B1(new_n772), .B2(G29), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT99), .B(G2067), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n711), .A2(G27), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n711), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2078), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n551), .A2(new_n692), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n692), .B2(G19), .ZN(new_n781));
  INV_X1    g356(.A(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n692), .A2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G168), .B2(new_n692), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n781), .A2(new_n782), .B1(new_n784), .B2(G1966), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT31), .B(G11), .Z(new_n786));
  XOR2_X1   g361(.A(KEYINPUT100), .B(G28), .Z(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(KEYINPUT30), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(G29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(KEYINPUT30), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n791), .B1(new_n711), .B2(new_n623), .C1(new_n764), .C2(new_n765), .ZN(new_n792));
  INV_X1    g367(.A(new_n781), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(G1341), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n766), .A2(new_n779), .A3(new_n785), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G4), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n600), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1348), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n784), .A2(G1966), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT101), .Z(new_n800));
  NOR4_X1   g375(.A1(new_n748), .A2(new_n795), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n725), .A2(new_n726), .A3(new_n731), .A4(new_n801), .ZN(G150));
  INV_X1    g377(.A(G150), .ZN(G311));
  NAND2_X1  g378(.A1(new_n529), .A2(G67), .ZN(new_n804));
  NAND2_X1  g379(.A1(G80), .A2(G543), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n522), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G93), .ZN(new_n807));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n517), .A2(new_n807), .B1(new_n519), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G860), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n600), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n547), .A2(new_n550), .ZN(new_n816));
  INV_X1    g391(.A(new_n810), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n551), .A2(new_n810), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n815), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT39), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT104), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(new_n811), .C1(new_n822), .C2(new_n821), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n813), .B1(new_n826), .B2(new_n827), .ZN(G145));
  XOR2_X1   g403(.A(new_n717), .B(KEYINPUT105), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n492), .A2(G142), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n487), .A2(G130), .ZN(new_n831));
  OAI221_X1 g406(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n481), .C2(G118), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n829), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n628), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n772), .B(new_n513), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n763), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n753), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n835), .A2(KEYINPUT107), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT107), .B1(new_n835), .B2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n835), .A2(new_n838), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n495), .B(G160), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(new_n623), .Z(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n841), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n835), .A2(new_n838), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT106), .B(G37), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g426(.A1(new_n817), .A2(G868), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n610), .B(new_n820), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n597), .B(G299), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n854), .B(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT109), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  XNOR2_X1  g437(.A(G166), .B(KEYINPUT108), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n691), .ZN(new_n864));
  XNOR2_X1  g439(.A(G290), .B(new_n583), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n864), .B(new_n865), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n861), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n859), .A2(new_n860), .A3(new_n867), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n852), .B1(new_n870), .B2(G868), .ZN(G295));
  AOI21_X1  g446(.A(new_n852), .B1(new_n870), .B2(G868), .ZN(G331));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n873));
  INV_X1    g448(.A(new_n849), .ZN(new_n874));
  INV_X1    g449(.A(new_n866), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n818), .A2(G301), .A3(new_n819), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(G301), .B1(new_n818), .B2(new_n819), .ZN(new_n878));
  OAI21_X1  g453(.A(G286), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(G168), .A3(new_n876), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n879), .A2(new_n881), .A3(new_n858), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n855), .B1(new_n879), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n881), .A3(new_n858), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n879), .A2(new_n881), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n866), .B(new_n885), .C1(new_n886), .C2(new_n855), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n874), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT110), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n884), .B2(new_n887), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n873), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n888), .A2(KEYINPUT43), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n892), .A2(KEYINPUT43), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT44), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(G397));
  INV_X1    g474(.A(G1384), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n507), .B2(new_n511), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(KEYINPUT111), .B(G40), .Z(new_n905));
  NAND3_X1  g480(.A1(new_n475), .A2(new_n483), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT112), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n475), .A2(new_n483), .A3(KEYINPUT112), .A4(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G2067), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n772), .B(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G1996), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n762), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n717), .B(new_n720), .Z(new_n918));
  OAI21_X1  g493(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n919), .A2(KEYINPUT126), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(KEYINPUT126), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n911), .A2(G1986), .A3(G290), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT48), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n911), .B1(new_n914), .B2(new_n763), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n912), .A2(new_n915), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n929), .B(KEYINPUT47), .Z(new_n930));
  NAND2_X1  g505(.A1(new_n718), .A2(new_n720), .ZN(new_n931));
  OAI22_X1  g506(.A1(new_n917), .A2(new_n931), .B1(G2067), .B2(new_n772), .ZN(new_n932));
  AOI211_X1 g507(.A(new_n924), .B(new_n930), .C1(new_n912), .C2(new_n932), .ZN(new_n933));
  OR2_X1    g508(.A1(G305), .A2(G1981), .ZN(new_n934));
  NAND2_X1  g509(.A1(G305), .A2(G1981), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n934), .A2(KEYINPUT49), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT49), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  INV_X1    g512(.A(G8), .ZN(new_n938));
  INV_X1    g513(.A(new_n901), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n910), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n936), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n691), .A2(G1976), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT52), .B1(new_n943), .B2(new_n940), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT115), .B1(new_n691), .B2(G1976), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n945), .B(new_n940), .C1(new_n943), .C2(KEYINPUT52), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G303), .A2(G8), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n910), .A2(new_n903), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n939), .A2(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(KEYINPUT113), .B(G1971), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n901), .A2(KEYINPUT50), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n901), .A2(KEYINPUT50), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n910), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT114), .B(G2090), .Z(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n949), .A2(G8), .A3(new_n952), .A4(new_n964), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n942), .A2(G1976), .A3(G288), .ZN(new_n966));
  INV_X1    g541(.A(new_n934), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n940), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT117), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n964), .A2(G8), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n951), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(G8), .A3(new_n952), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n949), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n953), .A2(KEYINPUT116), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n910), .A2(new_n903), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n954), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1966), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n960), .A2(G2084), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(G8), .A3(G168), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n974), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n970), .B1(new_n985), .B2(KEYINPUT63), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n972), .A2(new_n949), .A3(new_n973), .ZN(new_n987));
  INV_X1    g562(.A(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT63), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n969), .B1(new_n986), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n981), .A2(G168), .A3(new_n982), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(G8), .ZN(new_n994));
  AOI21_X1  g569(.A(G168), .B1(new_n981), .B2(new_n982), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT51), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n997), .A3(G8), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n955), .B2(G2078), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n960), .A2(KEYINPUT120), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT120), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n958), .A2(new_n1006), .A3(new_n910), .A4(new_n959), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1003), .A2(G2078), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI221_X1 g585(.A(new_n1004), .B1(new_n1008), .B2(G1961), .C1(new_n979), .C2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G171), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n974), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1000), .A2(new_n1002), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n989), .A2(new_n970), .A3(new_n990), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n992), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT56), .B(G2072), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n953), .A2(new_n954), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(G1956), .B2(new_n961), .ZN(new_n1019));
  XNOR2_X1  g594(.A(G299), .B(KEYINPUT57), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI211_X1 g596(.A(KEYINPUT118), .B(new_n901), .C1(new_n908), .C2(new_n909), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n910), .B2(new_n939), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n913), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT119), .ZN(new_n1026));
  INV_X1    g601(.A(G1348), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1005), .A2(new_n1027), .A3(new_n1007), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(new_n913), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1026), .A2(KEYINPUT121), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n600), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1021), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1020), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n1018), .C1(G1956), .C2(new_n961), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1036), .B1(new_n1035), .B2(KEYINPUT60), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT60), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1042), .B(new_n600), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1035), .A2(KEYINPUT60), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(new_n1044), .A3(new_n600), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1033), .A2(new_n1042), .A3(new_n1034), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1039), .A2(new_n1021), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT61), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1039), .A2(new_n1021), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n1022), .A2(new_n1024), .A3(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(KEYINPUT122), .C1(G1996), .C2(new_n955), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT122), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n955), .A2(G1996), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1022), .A2(new_n1024), .A3(new_n1058), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1056), .B1(new_n1065), .B2(new_n551), .ZN(new_n1066));
  AOI211_X1 g641(.A(KEYINPUT59), .B(new_n816), .C1(new_n1060), .C2(new_n1064), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1055), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT123), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1055), .B(new_n1070), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1040), .B1(new_n1050), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  INV_X1    g649(.A(G40), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n484), .A2(new_n1075), .A3(new_n1010), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n954), .A2(new_n903), .A3(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1004), .B(new_n1077), .C1(new_n1008), .C2(G1961), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G171), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(KEYINPUT54), .C1(new_n1011), .C2(G171), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n987), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1078), .A2(G171), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT54), .B1(new_n1082), .B2(new_n1012), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1074), .B1(new_n1084), .B2(new_n999), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1011), .A2(G171), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1078), .B2(G171), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n974), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1082), .A2(new_n1012), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1087), .ZN(new_n1091));
  AND4_X1   g666(.A1(new_n1074), .A2(new_n1089), .A3(new_n999), .A4(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1085), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1016), .B1(new_n1073), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n917), .A2(new_n918), .ZN(new_n1095));
  XOR2_X1   g670(.A(G290), .B(G1986), .Z(new_n1096));
  AOI21_X1  g671(.A(new_n911), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n933), .B1(new_n1094), .B2(new_n1097), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g673(.A(G319), .B1(new_n651), .B2(new_n652), .ZN(new_n1100));
  NOR2_X1   g674(.A1(G227), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g675(.A1(new_n689), .A2(new_n1101), .ZN(new_n1102));
  XOR2_X1   g676(.A(new_n1102), .B(KEYINPUT127), .Z(new_n1103));
  OAI211_X1 g677(.A(new_n1103), .B(new_n850), .C1(new_n893), .C2(new_n894), .ZN(G225));
  INV_X1    g678(.A(G225), .ZN(G308));
endmodule


