//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n209), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT64), .Z(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n207), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n227), .B(new_n233), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n224), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n231), .ZN(new_n255));
  NAND3_X1  g0055(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(G274), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT68), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(new_n260), .ZN(new_n265));
  INV_X1    g0065(.A(new_n260), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n257), .A2(new_n266), .A3(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n262), .B1(new_n268), .B2(G226), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT69), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT69), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G222), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n217), .B2(new_n279), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n272), .A2(new_n278), .A3(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT70), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT70), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n272), .A2(new_n278), .A3(new_n285), .A4(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n282), .B1(G223), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n255), .A2(new_n252), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n269), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n290), .A2(G179), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n231), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n207), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n296), .A2(new_n298), .B1(G150), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n203), .A2(G20), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n294), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(new_n293), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n206), .A2(G20), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(G50), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G50), .B2(new_n303), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(new_n290), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n291), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n309), .B(KEYINPUT9), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(G190), .B(new_n269), .C1(new_n288), .C2(new_n289), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT73), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n318), .A2(new_n319), .B1(new_n290), .B2(G200), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(KEYINPUT73), .A3(new_n317), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT72), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT10), .B1(new_n316), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n290), .A2(G200), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n315), .A2(KEYINPUT72), .ZN(new_n326));
  AND4_X1   g0126(.A1(new_n317), .A2(new_n324), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n313), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n305), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n296), .A2(new_n306), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n329), .A2(new_n330), .B1(new_n296), .B2(new_n303), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n270), .A2(new_n271), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT7), .B1(new_n332), .B2(new_n207), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n277), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(G68), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G58), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n211), .ZN(new_n338));
  OAI21_X1  g0138(.A(G20), .B1(new_n338), .B2(new_n201), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n299), .A2(G159), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n336), .A2(KEYINPUT16), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT78), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n275), .A2(new_n207), .A3(new_n277), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n334), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n341), .B1(new_n348), .B2(G68), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT78), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT16), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n294), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(G20), .B1(new_n272), .B2(new_n278), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n334), .B1(new_n353), .B2(KEYINPUT7), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G68), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n342), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n331), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n274), .A2(new_n213), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n275), .A2(new_n277), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(G223), .A3(new_n280), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT79), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G226), .A2(G1698), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n280), .A2(G223), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n361), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n289), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n257), .A2(new_n266), .A3(G232), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n261), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(G169), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n289), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n332), .A2(new_n366), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n374), .A2(KEYINPUT79), .B1(new_n274), .B2(new_n213), .ZN(new_n375));
  INV_X1    g0175(.A(new_n368), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n371), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(G179), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT18), .B1(new_n359), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n331), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n350), .B1(new_n349), .B2(KEYINPUT16), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n211), .B1(new_n347), .B2(new_n334), .ZN(new_n385));
  NOR4_X1   g0185(.A1(new_n385), .A2(KEYINPUT78), .A3(new_n341), .A4(new_n357), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n293), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT16), .B1(new_n355), .B2(new_n342), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n380), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n382), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G200), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n369), .B2(new_n371), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n377), .A2(new_n395), .A3(new_n378), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n383), .B(new_n397), .C1(new_n387), .C2(new_n388), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n352), .A2(new_n358), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n383), .A4(new_n397), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n212), .B1(new_n284), .B2(new_n286), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n272), .A2(new_n278), .A3(G232), .A4(new_n280), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n279), .B2(new_n219), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n373), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n262), .B1(new_n268), .B2(G244), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(KEYINPUT71), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT71), .B1(new_n407), .B2(new_n408), .ZN(new_n411));
  OAI21_X1  g0211(.A(G190), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n407), .A2(new_n408), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT71), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(G200), .A3(new_n409), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n296), .A2(new_n299), .B1(G20), .B2(G77), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT15), .B(G87), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n418), .A2(new_n297), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n294), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n305), .A2(G77), .A3(new_n306), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(G77), .B2(new_n303), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n412), .A2(new_n416), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G179), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n410), .B2(new_n411), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n415), .A2(new_n310), .A3(new_n409), .ZN(new_n427));
  INV_X1    g0227(.A(new_n423), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n392), .A2(new_n403), .A3(new_n424), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT77), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n297), .A2(new_n217), .B1(new_n207), .B2(G68), .ZN(new_n432));
  INV_X1    g0232(.A(new_n299), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n432), .A2(KEYINPUT75), .B1(new_n202), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n432), .A2(KEYINPUT75), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n293), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT11), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n305), .A2(G68), .A3(new_n306), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT12), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n304), .B2(new_n211), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n303), .A2(KEYINPUT12), .A3(G68), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n436), .A2(new_n437), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n438), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n272), .A2(new_n278), .A3(G232), .A4(G1698), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n272), .A2(new_n278), .A3(G226), .A4(new_n280), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G97), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n373), .ZN(new_n453));
  INV_X1    g0253(.A(new_n267), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT68), .B1(new_n257), .B2(new_n266), .ZN(new_n455));
  OAI21_X1  g0255(.A(G238), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n261), .A2(KEYINPUT74), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT74), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n257), .A2(new_n458), .A3(G274), .A4(new_n260), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n453), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT13), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n268), .A2(G238), .B1(new_n457), .B2(new_n459), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT13), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n453), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n465), .A3(G190), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n448), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n393), .B1(new_n462), .B2(new_n465), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n431), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n468), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(KEYINPUT77), .A3(new_n466), .A4(new_n448), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n462), .A2(new_n465), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT14), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(G169), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n462), .A2(new_n465), .A3(G179), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n474), .B1(new_n473), .B2(G169), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n447), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n328), .A2(new_n430), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT25), .B1(new_n304), .B2(new_n219), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n219), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n274), .A2(G1), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n304), .A2(new_n293), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n483), .A2(new_n484), .B1(new_n486), .B2(G107), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT84), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n213), .A2(KEYINPUT22), .A3(G20), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n272), .A2(new_n278), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n207), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT22), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n219), .A2(KEYINPUT23), .A3(G20), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT23), .B1(new_n219), .B2(G20), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT83), .B(KEYINPUT24), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n500), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n493), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n488), .B1(new_n504), .B2(new_n293), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n493), .B2(new_n498), .ZN(new_n506));
  AOI211_X1 g0306(.A(new_n500), .B(new_n497), .C1(new_n490), .C2(new_n492), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n488), .B(new_n293), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n487), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n259), .A2(G1), .ZN(new_n511));
  NAND2_X1  g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n257), .A2(new_n515), .A3(G264), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT86), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n257), .A2(new_n515), .A3(KEYINPUT86), .A4(G264), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n514), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n512), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n257), .A2(new_n523), .A3(G274), .A4(new_n511), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n214), .A2(new_n280), .ZN(new_n525));
  INV_X1    g0325(.A(G257), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G1698), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n525), .B(new_n527), .C1(new_n270), .C2(new_n271), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT85), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G294), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n373), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n524), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(G169), .B1(new_n521), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n534), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT88), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n518), .A2(new_n539), .A3(new_n519), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n518), .B2(new_n519), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n538), .B(G179), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(KEYINPUT87), .B(G169), .C1(new_n521), .C2(new_n534), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n537), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n510), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n487), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n293), .B1(new_n506), .B2(new_n507), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n549), .B2(new_n508), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT89), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n538), .A2(new_n551), .A3(new_n395), .A4(new_n520), .ZN(new_n552));
  INV_X1    g0352(.A(new_n533), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(new_n373), .A3(new_n531), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n554), .A2(new_n520), .A3(new_n395), .A4(new_n524), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT89), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n520), .A2(KEYINPUT88), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n534), .B1(new_n557), .B2(new_n540), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n552), .B(new_n556), .C1(new_n558), .C2(G200), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n546), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g0361(.A(KEYINPUT82), .B(G303), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n272), .B2(new_n278), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n220), .A2(G1698), .ZN(new_n564));
  OAI221_X1 g0364(.A(new_n564), .B1(G257), .B2(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n373), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n257), .A2(new_n515), .A3(G270), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n524), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n486), .A2(G116), .ZN(new_n571));
  INV_X1    g0371(.A(G116), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n304), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(G20), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n293), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G283), .ZN(new_n576));
  INV_X1    g0376(.A(G97), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n576), .B(new_n207), .C1(G33), .C2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT20), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  AND4_X1   g0379(.A1(KEYINPUT20), .A2(new_n578), .A3(new_n293), .A4(new_n574), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n571), .B(new_n573), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n570), .A2(new_n581), .A3(KEYINPUT21), .A4(G169), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(G179), .A3(new_n567), .A4(new_n569), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n214), .B1(new_n259), .B2(G1), .ZN(new_n585));
  INV_X1    g0385(.A(G274), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n206), .A2(new_n586), .A3(G45), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n257), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G238), .A2(G1698), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n218), .B2(G1698), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n361), .B1(G33), .B2(G116), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n593), .B2(new_n289), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(new_n395), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n212), .A2(new_n280), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n218), .A2(G1698), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n270), .C2(new_n271), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G116), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n373), .B1(new_n589), .B2(new_n257), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n393), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n361), .A2(new_n207), .A3(G68), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n207), .B1(new_n451), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(G97), .A2(G107), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n213), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n605), .B1(new_n297), .B2(new_n577), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n293), .B1(new_n304), .B2(new_n418), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n486), .A2(G87), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g0414(.A(new_n418), .B(KEYINPUT81), .Z(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n486), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n264), .A2(new_n588), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n289), .B1(new_n598), .B2(new_n599), .ZN(new_n619));
  OAI21_X1  g0419(.A(G169), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n590), .B(G179), .C1(new_n593), .C2(new_n289), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n603), .A2(new_n614), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n581), .B1(new_n570), .B2(G200), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n395), .B2(new_n570), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n570), .A2(G169), .A3(new_n581), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n584), .A2(new_n623), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n303), .A2(G97), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n486), .B2(G97), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT6), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G97), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n632), .A2(G97), .A3(G107), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n219), .A2(KEYINPUT80), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n219), .A2(KEYINPUT80), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n634), .A2(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(KEYINPUT80), .B(G107), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n607), .A2(KEYINPUT6), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n640), .A3(new_n633), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n641), .A3(G20), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n299), .A2(G77), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(G107), .B2(new_n354), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n631), .B1(new_n645), .B2(new_n294), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT4), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n218), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n272), .A2(new_n278), .A3(new_n280), .A4(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n272), .A2(new_n278), .A3(G250), .A4(G1698), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n280), .A2(G244), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n332), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n649), .A2(new_n650), .A3(new_n576), .A4(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(new_n373), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n257), .A2(new_n515), .A3(G257), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n524), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n310), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n653), .B2(new_n373), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n425), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n646), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n354), .A2(G107), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n293), .B1(new_n661), .B2(new_n644), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n658), .A2(G200), .ZN(new_n663));
  AOI211_X1 g0463(.A(G190), .B(new_n656), .C1(new_n653), .C2(new_n373), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n662), .B(new_n631), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n629), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n481), .A2(new_n561), .A3(new_n667), .ZN(G372));
  INV_X1    g0468(.A(new_n479), .ZN(new_n669));
  INV_X1    g0469(.A(new_n429), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n669), .B1(new_n472), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n403), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n392), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n322), .A2(new_n327), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n312), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n481), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT90), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT90), .B1(new_n620), .B2(new_n621), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n617), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n603), .A2(new_n614), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n646), .A2(new_n657), .A3(new_n659), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n617), .A2(new_n622), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT26), .B1(new_n660), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n685), .A2(new_n680), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n660), .A2(new_n665), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n680), .A2(new_n681), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n550), .B2(new_n559), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n628), .A2(new_n583), .A3(new_n582), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n510), .B2(new_n545), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n690), .B(new_n692), .C1(new_n694), .C2(KEYINPUT91), .ZN(new_n695));
  INV_X1    g0495(.A(new_n693), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n546), .A2(KEYINPUT91), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n689), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n676), .B1(new_n677), .B2(new_n699), .ZN(G369));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n581), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n693), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n696), .A2(new_n625), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n701), .B(new_n709), .C1(new_n710), .C2(new_n708), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n701), .B2(new_n709), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n707), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n561), .B1(new_n550), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n546), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n510), .A2(new_n545), .A3(new_n715), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n696), .A2(new_n707), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n561), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(G399));
  NAND3_X1  g0522(.A1(new_n225), .A2(KEYINPUT93), .A3(new_n258), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT93), .B1(new_n225), .B2(new_n258), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n608), .A2(G116), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n726), .A2(new_n206), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n229), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n726), .ZN(new_n731));
  XNOR2_X1  g0531(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n694), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n690), .A3(new_n692), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n684), .B1(new_n682), .B2(new_n683), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n660), .A2(new_n687), .A3(KEYINPUT26), .ZN(new_n737));
  INV_X1    g0537(.A(new_n680), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n707), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n699), .A2(new_n707), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n742), .B2(KEYINPUT29), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n567), .A2(new_n569), .A3(G179), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n601), .B1(new_n532), .B2(new_n533), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n557), .A2(new_n540), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n746), .A2(KEYINPUT30), .A3(new_n747), .A4(new_n658), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT96), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n570), .A2(new_n425), .A3(new_n594), .ZN(new_n750));
  OR3_X1    g0550(.A1(new_n558), .A2(new_n750), .A3(new_n658), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n746), .A2(new_n747), .A3(new_n658), .ZN(new_n752));
  XOR2_X1   g0552(.A(KEYINPUT95), .B(KEYINPUT30), .Z(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n749), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n748), .A2(KEYINPUT96), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n707), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g0559(.A(KEYINPUT31), .B(new_n707), .C1(new_n755), .C2(new_n756), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n667), .A2(new_n546), .A3(new_n560), .A4(new_n715), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G330), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n743), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n733), .B1(new_n764), .B2(G1), .ZN(G364));
  AND2_X1   g0565(.A1(new_n207), .A2(G13), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n206), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n726), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n714), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n712), .A2(new_n713), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT101), .Z(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n712), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n279), .A2(G355), .A3(new_n225), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G116), .B2(new_n225), .ZN(new_n780));
  INV_X1    g0580(.A(new_n225), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n361), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n230), .B2(new_n259), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n247), .A2(new_n259), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n780), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n231), .B1(G20), .B2(new_n310), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n775), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n769), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n395), .A2(G179), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n207), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n207), .A2(G190), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(new_n425), .A3(new_n393), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n794), .A2(G294), .B1(new_n797), .B2(G329), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n207), .A2(new_n425), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(new_n395), .A3(G200), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(new_n802), .B2(KEYINPUT100), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(KEYINPUT100), .B2(new_n802), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n799), .A2(G190), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n393), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n279), .B1(G326), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(G200), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n795), .A2(G179), .A3(new_n393), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n809), .A2(G322), .B1(new_n811), .B2(G311), .ZN(new_n812));
  AOI21_X1  g0612(.A(KEYINPUT98), .B1(new_n425), .B2(G200), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n207), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n425), .A2(KEYINPUT98), .A3(G200), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(G190), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n395), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G283), .A2(new_n817), .B1(new_n818), .B2(G303), .ZN(new_n819));
  AND4_X1   g0619(.A1(new_n798), .A2(new_n808), .A3(new_n812), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(G87), .ZN(new_n821));
  INV_X1    g0621(.A(new_n817), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n279), .C1(new_n822), .C2(new_n219), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT99), .Z(new_n824));
  XOR2_X1   g0624(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n825));
  NAND3_X1  g0625(.A1(new_n797), .A2(G159), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n809), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n211), .B2(new_n800), .C1(new_n827), .C2(new_n337), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n806), .A2(G50), .B1(new_n811), .B2(G77), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n577), .B2(new_n793), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n825), .B1(new_n797), .B2(G159), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n820), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n791), .B1(new_n834), .B2(new_n788), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n778), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n772), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  NOR2_X1   g0638(.A1(new_n788), .A2(new_n773), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n769), .B1(G77), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n806), .A2(G137), .B1(new_n811), .B2(G159), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n842), .B1(new_n843), .B2(new_n827), .C1(new_n844), .C2(new_n800), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT34), .Z(new_n846));
  NAND2_X1  g0646(.A1(new_n818), .A2(G50), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n817), .A2(G68), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n797), .A2(G132), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n332), .B1(new_n794), .B2(G58), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(G294), .ZN(new_n852));
  INV_X1    g0652(.A(G311), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n827), .A2(new_n852), .B1(new_n796), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G303), .B2(new_n806), .ZN(new_n855));
  INV_X1    g0655(.A(new_n800), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n279), .B1(G283), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n794), .A2(G97), .B1(new_n811), .B2(G116), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n818), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n213), .A2(new_n822), .B1(new_n860), .B2(new_n219), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n846), .A2(new_n851), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n841), .B1(new_n862), .B2(new_n788), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT102), .ZN(new_n864));
  AND4_X1   g0664(.A1(new_n428), .A2(new_n426), .A3(new_n427), .A4(new_n715), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n423), .A2(new_n715), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT103), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n424), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n865), .B1(new_n429), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n864), .B1(new_n774), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n742), .A2(new_n869), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n698), .A2(new_n715), .A3(new_n869), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n763), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n769), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n871), .A2(new_n763), .A3(new_n873), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n870), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT104), .Z(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(G384));
  AND2_X1   g0680(.A1(new_n638), .A2(new_n641), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT35), .ZN(new_n883));
  OAI211_X1 g0683(.A(G116), .B(new_n232), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n883), .B2(new_n882), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT36), .ZN(new_n886));
  OR3_X1    g0686(.A1(new_n229), .A2(new_n217), .A3(new_n338), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n202), .A2(G68), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n206), .B(G13), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n357), .B1(new_n385), .B2(new_n341), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n331), .B1(new_n352), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n398), .B1(new_n892), .B2(new_n381), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n705), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n389), .A2(new_n380), .ZN(new_n896));
  INV_X1    g0696(.A(new_n705), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n389), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n896), .A2(new_n898), .A3(new_n899), .A4(new_n398), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n382), .A2(new_n391), .A3(new_n400), .A4(new_n402), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n902), .A2(KEYINPUT106), .A3(new_n894), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT106), .B1(new_n902), .B2(new_n894), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(KEYINPUT38), .B(new_n901), .C1(new_n903), .C2(new_n904), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n447), .A2(new_n707), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n472), .B2(new_n479), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n472), .A2(new_n479), .A3(new_n910), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT105), .ZN(new_n915));
  INV_X1    g0715(.A(new_n865), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n872), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n915), .B1(new_n872), .B2(new_n916), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n909), .B(new_n914), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n392), .A2(new_n897), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT107), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n398), .B1(new_n359), .B2(new_n381), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n359), .A2(new_n705), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT37), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(KEYINPUT108), .A3(new_n900), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n902), .A2(new_n925), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT108), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(KEYINPUT37), .C1(new_n924), .C2(new_n925), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n906), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n908), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n669), .A2(new_n715), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n919), .A2(KEYINPUT107), .A3(new_n920), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n923), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n481), .B(new_n741), .C1(KEYINPUT29), .C2(new_n742), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n676), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n762), .A2(new_n869), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n472), .A2(new_n479), .A3(new_n910), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n946), .A2(new_n911), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT40), .B1(new_n909), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n932), .A2(new_n908), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n914), .A2(KEYINPUT40), .A3(new_n762), .A4(new_n869), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n481), .A2(new_n762), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n953), .B1(new_n949), .B2(new_n952), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(G330), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n944), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n206), .B2(new_n766), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n944), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n890), .B1(new_n958), .B2(new_n959), .ZN(G367));
  NOR2_X1   g0760(.A1(new_n614), .A2(new_n715), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n738), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(KEYINPUT109), .C1(new_n691), .C2(new_n961), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(KEYINPUT109), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n777), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n822), .A2(new_n577), .ZN(new_n966));
  INV_X1    g0766(.A(new_n806), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n853), .A2(new_n967), .B1(new_n827), .B2(new_n562), .ZN(new_n968));
  INV_X1    g0768(.A(G283), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n332), .B1(new_n810), .B2(new_n969), .C1(new_n852), .C2(new_n800), .ZN(new_n970));
  INV_X1    g0770(.A(G317), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n793), .A2(new_n219), .B1(new_n796), .B2(new_n971), .ZN(new_n972));
  OR4_X1    g0772(.A1(new_n966), .A2(new_n968), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n818), .A2(G116), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT46), .Z(new_n975));
  OAI22_X1  g0775(.A1(new_n827), .A2(new_n844), .B1(new_n967), .B2(new_n843), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G137), .B2(new_n797), .ZN(new_n977));
  INV_X1    g0777(.A(new_n279), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G159), .B2(new_n856), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n794), .A2(G68), .B1(new_n811), .B2(G50), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n337), .A2(new_n860), .B1(new_n822), .B2(new_n217), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n973), .A2(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n788), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n789), .B1(new_n225), .B2(new_n418), .C1(new_n783), .C2(new_n243), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n965), .A2(new_n769), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n646), .A2(new_n707), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n690), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n683), .A2(new_n707), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n561), .A3(new_n720), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT42), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n660), .B1(new_n989), .B2(new_n546), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n715), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(KEYINPUT42), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT111), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n964), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT110), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT112), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n998), .B(new_n1003), .C1(new_n999), .C2(new_n964), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n718), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n991), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n1002), .B2(new_n1001), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1007), .A2(new_n1011), .A3(new_n1008), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n721), .A2(new_n719), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n991), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT44), .Z(new_n1017));
  NOR2_X1   g0817(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(new_n1005), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n721), .B1(new_n717), .B2(new_n720), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(new_n714), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n764), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n764), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n726), .B(KEYINPUT41), .Z(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n768), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n987), .B1(new_n1013), .B2(new_n1029), .ZN(G387));
  OR2_X1    g0830(.A1(new_n717), .A2(new_n776), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n782), .B1(new_n240), .B2(new_n259), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n279), .A2(new_n225), .A3(new_n728), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n295), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT50), .B1(new_n295), .B2(G50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n727), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1034), .A2(new_n1038), .B1(new_n219), .B2(new_n781), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n769), .B1(new_n1039), .B2(new_n790), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n615), .A2(new_n794), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n202), .B2(new_n827), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT113), .ZN(new_n1043));
  INV_X1    g0843(.A(G159), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n967), .A2(new_n1044), .B1(new_n796), .B2(new_n844), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n810), .A2(new_n211), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n361), .B1(new_n800), .B2(new_n295), .ZN(new_n1047));
  NOR4_X1   g0847(.A1(new_n966), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1043), .B(new_n1048), .C1(new_n217), .C2(new_n860), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n800), .A2(new_n853), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n827), .A2(new_n971), .B1(new_n562), .B2(new_n810), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(G322), .C2(new_n806), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT48), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(KEYINPUT48), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n818), .A2(G294), .B1(G283), .B2(new_n794), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT114), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT49), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n361), .B1(new_n797), .B2(G326), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n572), .C2(new_n822), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1057), .A2(KEYINPUT49), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1049), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1040), .B1(new_n1062), .B2(new_n788), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1031), .A2(new_n1063), .B1(new_n1023), .B2(new_n768), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1024), .A2(new_n726), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n764), .A2(new_n1023), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(G393));
  NAND2_X1  g0867(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1025), .A2(new_n726), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT115), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n767), .B1(new_n1021), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1021), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1015), .A2(new_n775), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n332), .B1(new_n797), .B2(G143), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n822), .B2(new_n213), .C1(new_n211), .C2(new_n860), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT116), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G150), .A2(new_n806), .B1(new_n809), .B2(G159), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT51), .Z(new_n1078));
  NAND2_X1  g0878(.A1(new_n811), .A2(new_n296), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G77), .A2(new_n794), .B1(new_n856), .B2(G50), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G311), .A2(new_n809), .B1(new_n806), .B2(G317), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT52), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G107), .A2(new_n817), .B1(new_n818), .B2(G283), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n562), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n279), .B1(new_n1085), .B2(new_n856), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n794), .A2(G116), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n811), .A2(G294), .B1(new_n797), .B2(G322), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1076), .A2(new_n1081), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n788), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n789), .B1(new_n577), .B2(new_n225), .C1(new_n783), .C2(new_n250), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1073), .A2(new_n1091), .A3(new_n769), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1069), .A2(new_n1072), .A3(new_n1093), .ZN(G390));
  NAND3_X1  g0894(.A1(new_n762), .A2(G330), .A3(new_n869), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1095), .A2(new_n947), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1098), .A2(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n865), .B1(new_n740), .B2(new_n869), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n937), .B1(new_n1100), .B2(new_n947), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(new_n950), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1097), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n935), .A2(new_n936), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n872), .A2(new_n916), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n872), .A2(new_n915), .A3(new_n916), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n947), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1104), .B1(new_n1108), .B2(new_n938), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1102), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n1096), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1103), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1095), .A2(new_n947), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1096), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n917), .B2(new_n918), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1096), .A2(new_n1100), .A3(new_n1113), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n481), .A2(G330), .A3(new_n762), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n942), .A2(new_n676), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT117), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1112), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n726), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1112), .B2(new_n1121), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1103), .A2(new_n1111), .A3(new_n768), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1104), .A2(new_n773), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n769), .B1(new_n296), .B2(new_n840), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n978), .B1(G137), .B2(new_n856), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1130), .A2(new_n796), .B1(new_n810), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G128), .B2(new_n806), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G159), .A2(new_n794), .B1(new_n809), .B2(G132), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1129), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n860), .A2(new_n844), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT53), .Z(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(G50), .C2(new_n817), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1138), .A2(KEYINPUT118), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(KEYINPUT118), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n967), .A2(new_n969), .B1(new_n217), .B2(new_n793), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n279), .B(new_n1141), .C1(G107), .C2(new_n856), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n827), .A2(new_n572), .B1(new_n796), .B2(new_n852), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G97), .B2(new_n811), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1142), .A2(new_n821), .A3(new_n848), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1139), .A2(new_n1140), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1128), .B1(new_n1146), .B2(new_n788), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1127), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1125), .A2(new_n1126), .A3(new_n1148), .ZN(G378));
  INV_X1    g0949(.A(KEYINPUT122), .ZN(new_n1150));
  OAI21_X1  g0950(.A(G330), .B1(new_n950), .B2(new_n951), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n949), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n902), .A2(new_n894), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT106), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n902), .A2(KEYINPUT106), .A3(new_n894), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT38), .B1(new_n1157), .B2(new_n901), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n908), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n948), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT40), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n945), .A2(new_n947), .A3(new_n1161), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n713), .B1(new_n1163), .B2(new_n933), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(KEYINPUT122), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g0965(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n309), .A2(new_n705), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT55), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n328), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n328), .A2(new_n1169), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1167), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1172), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n1166), .A3(new_n1170), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1152), .A2(new_n1165), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1176), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1178), .A2(KEYINPUT122), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n941), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n940), .A2(new_n939), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1182), .A2(new_n1177), .A3(new_n923), .A4(new_n1179), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n768), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n769), .B1(G50), .B2(new_n840), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n615), .A2(new_n811), .B1(G97), .B2(new_n856), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT119), .Z(new_n1187));
  OAI211_X1 g0987(.A(new_n258), .B(new_n332), .C1(new_n793), .C2(new_n211), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n806), .A2(G116), .B1(new_n797), .B2(G283), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n219), .B2(new_n827), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n337), .A2(new_n822), .B1(new_n860), .B2(new_n217), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1192), .A2(KEYINPUT58), .ZN(new_n1193));
  INV_X1    g0993(.A(G128), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n827), .A2(new_n1194), .B1(new_n967), .B2(new_n1130), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G137), .B2(new_n811), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G150), .A2(new_n794), .B1(new_n856), .B2(G132), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n860), .C2(new_n1131), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n797), .C2(G124), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n822), .B2(new_n1044), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT120), .Z(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1192), .A2(KEYINPUT58), .ZN(new_n1205));
  AOI21_X1  g1005(.A(G50), .B1(new_n274), .B2(new_n258), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n361), .B2(G41), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1193), .A2(new_n1204), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1185), .B1(new_n1208), .B2(new_n788), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1176), .B2(new_n774), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1184), .A2(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1103), .A2(new_n1111), .A3(new_n1117), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1120), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1214), .A2(KEYINPUT57), .A3(new_n1183), .A4(new_n1181), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n726), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1211), .B1(new_n1215), .B2(new_n1217), .ZN(G375));
  NAND2_X1  g1018(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1115), .A2(new_n1119), .A3(new_n1116), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1028), .A3(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1041), .B(new_n978), .C1(new_n572), .C2(new_n800), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n217), .A2(new_n822), .B1(new_n860), .B2(new_n577), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n811), .A2(G107), .B1(new_n797), .B2(G303), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n969), .B2(new_n827), .C1(new_n852), .C2(new_n967), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G132), .A2(new_n806), .B1(new_n809), .B2(G137), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n202), .B2(new_n793), .C1(new_n1194), .C2(new_n796), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n337), .A2(new_n822), .B1(new_n860), .B2(new_n1044), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n361), .B1(new_n810), .B2(new_n844), .C1(new_n800), .C2(new_n1131), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n788), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1232), .B(new_n769), .C1(G68), .C2(new_n840), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n947), .B2(new_n773), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1117), .B2(new_n768), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1221), .A2(new_n1235), .ZN(G381));
  OR2_X1    g1036(.A1(G375), .A2(G378), .ZN(new_n1237));
  OR4_X1    g1037(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G387), .A2(new_n1237), .A3(G381), .A4(new_n1238), .ZN(G407));
  OAI211_X1 g1039(.A(G407), .B(G213), .C1(new_n1237), .C2(G343), .ZN(G409));
  AOI21_X1  g1040(.A(new_n1027), .B1(new_n1025), .B2(new_n764), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1010), .B(new_n1012), .C1(new_n1241), .C2(new_n768), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n987), .A3(G390), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G390), .B1(new_n1242), .B2(new_n987), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(G393), .B(new_n837), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1244), .A2(new_n1245), .B1(KEYINPUT125), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1245), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1246), .B(KEYINPUT125), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n1243), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G213), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(G343), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1125), .A2(new_n1126), .A3(new_n1148), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT123), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1184), .A2(new_n1256), .A3(new_n1210), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1214), .A2(new_n1028), .A3(new_n1183), .A4(new_n1181), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1256), .B1(new_n1184), .B2(new_n1210), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1255), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1211), .C1(new_n1215), .C2(new_n1217), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1254), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1219), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1220), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1117), .A2(new_n1266), .A3(new_n1120), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(new_n1123), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n879), .A3(new_n1235), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n879), .B1(new_n1270), .B2(new_n1235), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1264), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1273), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(KEYINPUT124), .A3(new_n1271), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT62), .B1(new_n1263), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1254), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  AOI211_X1 g1082(.A(KEYINPUT126), .B(new_n1254), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1278), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1254), .A2(G2897), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1272), .A2(new_n1273), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1277), .B2(new_n1287), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1252), .B1(new_n1286), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT61), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1288), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1287), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1294), .B1(new_n1298), .B2(new_n1263), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT63), .B1(new_n1263), .B2(new_n1277), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1284), .A2(KEYINPUT63), .A3(new_n1277), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1293), .A2(new_n1303), .ZN(G405));
  NAND2_X1  g1104(.A1(new_n1262), .A2(KEYINPUT127), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G375), .A2(new_n1255), .ZN(new_n1306));
  XOR2_X1   g1106(.A(new_n1305), .B(new_n1306), .Z(new_n1307));
  NOR2_X1   g1107(.A1(new_n1307), .A2(new_n1296), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1305), .B(new_n1306), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1309), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1252), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1307), .A2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1313), .B(new_n1251), .C1(new_n1296), .C2(new_n1307), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1314), .ZN(G402));
endmodule


