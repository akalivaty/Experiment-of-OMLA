//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  OR3_X1    g003(.A1(new_n204), .A2(KEYINPUT68), .A3(KEYINPUT26), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(KEYINPUT26), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT68), .B1(new_n204), .B2(KEYINPUT26), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT27), .B(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT28), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n212), .B(KEYINPUT66), .Z(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(KEYINPUT28), .A3(new_n211), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n214), .B(KEYINPUT67), .Z(new_n215));
  OAI211_X1 g014(.A(new_n202), .B(new_n209), .C1(new_n213), .C2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(G127gat), .A2(G134gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G127gat), .A2(G134gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G113gat), .B(G120gat), .Z(new_n220));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G113gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G120gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT69), .B(G120gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G113gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(new_n221), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT70), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n231));
  OAI21_X1  g030(.A(G113gat), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n224), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT1), .B1(new_n217), .B2(new_n218), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n222), .B1(new_n229), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n204), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n203), .A2(KEYINPUT23), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n206), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT64), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n202), .A2(KEYINPUT24), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n202), .A2(KEYINPUT24), .ZN(new_n244));
  NOR2_X1   g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n243), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n241), .A2(KEYINPUT64), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT25), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n206), .B1(new_n204), .B2(new_n238), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n252), .A2(new_n239), .A3(new_n247), .A4(new_n253), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n248), .A2(new_n250), .B1(new_n254), .B2(KEYINPUT25), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n216), .A2(new_n237), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n237), .B1(new_n216), .B2(new_n255), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G227gat), .ZN(new_n260));
  INV_X1    g059(.A(G233gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT34), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT32), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n257), .A2(new_n258), .ZN(new_n266));
  INV_X1    g065(.A(new_n262), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT32), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT34), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n259), .A2(new_n262), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n268), .A2(KEYINPUT33), .ZN(new_n274));
  XOR2_X1   g073(.A(G15gat), .B(G43gat), .Z(new_n275));
  XNOR2_X1  g074(.A(G71gat), .B(G99gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n272), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n270), .A3(new_n280), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n273), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n279), .B1(new_n273), .B2(new_n281), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT36), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT36), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(new_n282), .B2(new_n283), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n289));
  NAND2_X1  g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290));
  INV_X1    g089(.A(G155gat), .ZN(new_n291));
  INV_X1    g090(.A(G162gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G141gat), .B(G148gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n290), .B(new_n293), .C1(new_n294), .C2(KEYINPUT2), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT74), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n290), .B1(new_n293), .B2(KEYINPUT2), .ZN(new_n297));
  INV_X1    g096(.A(G148gat), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n298), .A2(G141gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(G141gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(new_n299), .B2(new_n300), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n290), .A4(new_n293), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n296), .A2(new_n301), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n229), .A2(new_n236), .ZN(new_n307));
  INV_X1    g106(.A(new_n222), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT76), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310));
  AOI211_X1 g109(.A(new_n310), .B(new_n222), .C1(new_n229), .C2(new_n236), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n306), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT79), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n296), .A2(new_n301), .A3(new_n305), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n237), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT79), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n316), .B(new_n306), .C1(new_n309), .C2(new_n311), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G225gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n289), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(new_n314), .B2(new_n237), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(KEYINPUT77), .ZN(new_n325));
  INV_X1    g124(.A(new_n236), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n234), .B1(new_n233), .B2(new_n235), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n308), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT4), .B1(new_n328), .B2(new_n306), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n237), .A3(new_n323), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n325), .B1(KEYINPUT77), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n334));
  OAI22_X1  g133(.A1(new_n309), .A2(new_n311), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT75), .B1(new_n306), .B2(KEYINPUT3), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n336), .A2(new_n334), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n319), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n322), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n328), .A2(KEYINPUT4), .A3(new_n306), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT77), .B1(new_n340), .B2(new_n324), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n324), .A2(KEYINPUT77), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n334), .ZN(new_n344));
  OAI221_X1 g143(.A(new_n344), .B1(new_n333), .B2(new_n334), .C1(new_n309), .C2(new_n311), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT78), .A4(new_n319), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n321), .A2(new_n339), .A3(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(G57gat), .B(G85gat), .Z(new_n348));
  XNOR2_X1  g147(.A(G1gat), .B(G29gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT80), .B(KEYINPUT0), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT81), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n350), .B(new_n352), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n345), .A2(new_n289), .A3(new_n319), .A4(new_n331), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT6), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n354), .B1(new_n347), .B2(new_n355), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n347), .A2(KEYINPUT82), .A3(new_n354), .A4(new_n355), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(KEYINPUT6), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n216), .A2(new_n255), .ZN(new_n366));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT72), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G197gat), .B(G204gat), .Z(new_n373));
  NAND2_X1  g172(.A1(G211gat), .A2(G218gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT22), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(G211gat), .A2(G218gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n377), .B(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT71), .B(new_n379), .C1(new_n373), .C2(new_n376), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n372), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n383), .B(new_n382), .C1(new_n369), .C2(new_n371), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT73), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT73), .B1(new_n385), .B2(new_n386), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OR3_X1    g191(.A1(new_n387), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n385), .B2(new_n386), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT30), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n394), .A2(KEYINPUT30), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n365), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G228gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(new_n261), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n370), .B1(new_n306), .B2(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n402), .B(KEYINPUT85), .Z(new_n403));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n380), .B2(KEYINPUT29), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n306), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n400), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n404), .B1(new_n384), .B2(KEYINPUT29), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n306), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n400), .A3(new_n402), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OR3_X1    g210(.A1(new_n407), .A2(G22gat), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(G22gat), .B1(new_n407), .B2(new_n411), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT84), .B(G50gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT86), .B(G22gat), .C1(new_n407), .C2(new_n411), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(KEYINPUT86), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n412), .A2(new_n413), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n288), .B1(new_n398), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT37), .B1(new_n385), .B2(new_n386), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n427), .A2(KEYINPUT38), .A3(new_n392), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT37), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n394), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n431));
  AND4_X1   g230(.A1(new_n431), .A2(new_n358), .A3(new_n360), .A4(new_n361), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n347), .A2(new_n354), .A3(new_n355), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n359), .B1(new_n433), .B2(KEYINPUT82), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n434), .B2(new_n358), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n363), .B(new_n430), .C1(new_n432), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT89), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n387), .A2(new_n388), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n440), .B2(new_n392), .ZN(new_n441));
  INV_X1    g240(.A(new_n427), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n440), .A2(new_n438), .A3(new_n392), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT38), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n362), .A2(KEYINPUT88), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n434), .A2(new_n431), .A3(new_n358), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT89), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n363), .A4(new_n430), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n437), .A2(new_n445), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n319), .B1(new_n345), .B2(new_n331), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n453), .B(KEYINPUT39), .C1(new_n320), .C2(new_n318), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT39), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n353), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OR3_X1    g256(.A1(new_n457), .A2(KEYINPUT87), .A3(KEYINPUT40), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(KEYINPUT87), .B2(KEYINPUT40), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n458), .A2(new_n360), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n424), .B1(new_n460), .B2(new_n397), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n426), .B1(new_n451), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n448), .A2(new_n363), .ZN(new_n464));
  INV_X1    g263(.A(new_n397), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n425), .A2(new_n465), .A3(new_n284), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n398), .A2(KEYINPUT35), .A3(new_n425), .A4(new_n284), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT100), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT93), .B(G36gat), .Z(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G29gat), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(KEYINPUT92), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(KEYINPUT92), .ZN(new_n476));
  OR3_X1    g275(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n473), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT15), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT94), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G43gat), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT95), .B1(new_n484), .B2(G50gat), .ZN(new_n485));
  OR3_X1    g284(.A1(new_n480), .A2(KEYINPUT15), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n477), .A2(KEYINPUT96), .ZN(new_n487));
  OR4_X1    g286(.A1(KEYINPUT96), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n474), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n480), .B1(KEYINPUT15), .B2(new_n485), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n486), .A2(new_n489), .A3(new_n473), .A4(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT97), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT16), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(G1gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(G1gat), .B2(new_n494), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G8gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n492), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n481), .B(KEYINPUT94), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT17), .B1(new_n483), .B2(new_n492), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n500), .B1(new_n506), .B2(new_n499), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT18), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n501), .A2(new_n502), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n498), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n493), .A2(new_n499), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT99), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(new_n508), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  OR3_X1    g317(.A1(new_n493), .A2(KEYINPUT99), .A3(new_n499), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n507), .A2(KEYINPUT18), .A3(new_n508), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n511), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523));
  INV_X1    g322(.A(G197gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XOR2_X1   g324(.A(KEYINPUT11), .B(G169gat), .Z(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n527), .B(KEYINPUT12), .Z(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n522), .A2(KEYINPUT91), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n522), .B2(KEYINPUT91), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n471), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n528), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT100), .A3(new_n530), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n470), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G127gat), .B(G155gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G211gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  INV_X1    g341(.A(G71gat), .ZN(new_n543));
  INV_X1    g342(.A(G78gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT102), .B(G64gat), .ZN(new_n548));
  INV_X1    g347(.A(G57gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT103), .Z(new_n551));
  AND2_X1   g350(.A1(new_n549), .A2(G64gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT101), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n542), .B(new_n545), .C1(new_n555), .C2(new_n546), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n499), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(G183gat), .ZN(new_n560));
  INV_X1    g359(.A(G183gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n561), .A3(new_n499), .ZN(new_n562));
  INV_X1    g361(.A(G231gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(new_n261), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n558), .B2(new_n499), .ZN(new_n566));
  AOI211_X1 g365(.A(G183gat), .B(new_n498), .C1(new_n557), .C2(KEYINPUT21), .ZN(new_n567));
  OAI22_X1  g366(.A1(new_n566), .A2(new_n567), .B1(new_n563), .B2(new_n261), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n541), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n557), .A2(KEYINPUT21), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT104), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n571), .B(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n565), .A2(new_n568), .A3(new_n541), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n574), .ZN(new_n577));
  INV_X1    g376(.A(new_n575), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(new_n569), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT107), .ZN(new_n581));
  INV_X1    g380(.A(G85gat), .ZN(new_n582));
  INV_X1    g381(.A(G92gat), .ZN(new_n583));
  OR3_X1    g382(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT7), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT7), .B1(new_n582), .B2(new_n583), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n584), .A2(new_n585), .B1(KEYINPUT8), .B2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT106), .B(G92gat), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(G85gat), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G99gat), .B(G106gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n506), .A2(new_n593), .B1(KEYINPUT41), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n512), .A2(new_n592), .ZN(new_n597));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n598), .B1(new_n596), .B2(new_n597), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n581), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n597), .ZN(new_n603));
  INV_X1    g402(.A(new_n598), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(KEYINPUT107), .A3(new_n599), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n595), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT105), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n602), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n605), .A2(KEYINPUT107), .A3(new_n599), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n580), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n615), .A2(KEYINPUT108), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(KEYINPUT108), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n557), .A2(new_n592), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n553), .A2(new_n556), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n593), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT109), .Z(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n619), .A2(new_n627), .A3(new_n621), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n557), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n625), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n618), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n538), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n365), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g443(.A1(new_n641), .A2(new_n465), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT16), .B(G8gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(KEYINPUT42), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(KEYINPUT110), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT110), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n641), .B2(new_n465), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n649), .B1(new_n653), .B2(G8gat), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n646), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(G1325gat));
  INV_X1    g455(.A(G15gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n641), .A2(new_n657), .A3(new_n288), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n284), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n657), .B2(new_n659), .ZN(G1326gat));
  NOR2_X1   g459(.A1(new_n641), .A2(new_n425), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G22gat), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  AND3_X1   g463(.A1(new_n611), .A2(KEYINPUT114), .A3(new_n613), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT114), .B1(new_n611), .B2(new_n613), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n668), .B(new_n669), .C1(new_n462), .C2(new_n469), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n470), .A2(new_n614), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n535), .A2(new_n530), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n580), .A2(new_n639), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676), .B2(new_n364), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  NOR4_X1   g477(.A1(new_n470), .A2(new_n614), .A3(new_n537), .A4(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(G29gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n365), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(KEYINPUT112), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(KEYINPUT112), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n683), .B1(new_n682), .B2(new_n684), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n677), .B1(new_n685), .B2(new_n686), .ZN(G1328gat));
  INV_X1    g486(.A(new_n537), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n688), .A3(new_n675), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(new_n472), .A3(new_n465), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT46), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n472), .B1(new_n676), .B2(new_n465), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1329gat));
  INV_X1    g492(.A(new_n284), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n689), .A2(G43gat), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n288), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n673), .A2(new_n696), .A3(new_n674), .A4(new_n675), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(G43gat), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g498(.A1(new_n425), .A2(G50gat), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n689), .A2(KEYINPUT115), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n689), .A2(KEYINPUT115), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G50gat), .B1(new_n676), .B2(new_n425), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n703), .B2(new_n704), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(G1331gat));
  NOR2_X1   g507(.A1(new_n470), .A2(new_n674), .ZN(new_n709));
  INV_X1    g508(.A(new_n639), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n618), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n364), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n549), .ZN(G1332gat));
  NOR2_X1   g513(.A1(new_n712), .A2(new_n465), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  AND2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n715), .B2(new_n716), .ZN(G1333gat));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT116), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n712), .B2(new_n694), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n709), .A2(KEYINPUT116), .A3(new_n284), .A4(new_n711), .ZN(new_n723));
  AOI21_X1  g522(.A(G71gat), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G71gat), .B1(new_n712), .B2(new_n288), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n720), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n726), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n724), .A2(KEYINPUT50), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n727), .A2(new_n729), .ZN(G1334gat));
  NOR2_X1   g529(.A1(new_n712), .A2(new_n425), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(new_n544), .ZN(G1335gat));
  NOR3_X1   g531(.A1(new_n674), .A2(new_n580), .A3(new_n710), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n673), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(new_n582), .A3(new_n364), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n674), .A2(new_n580), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n671), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n671), .A2(KEYINPUT51), .A3(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n365), .A3(new_n639), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n735), .B1(new_n742), .B2(new_n582), .ZN(G1336gat));
  OAI21_X1  g542(.A(new_n589), .B1(new_n734), .B2(new_n465), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n397), .A2(new_n583), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n710), .B(new_n746), .C1(new_n739), .C2(new_n740), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT52), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n741), .A2(new_n639), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n749), .B(new_n744), .C1(new_n750), .C2(new_n746), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(G1337gat));
  NAND2_X1  g551(.A1(new_n451), .A2(new_n461), .ZN(new_n753));
  INV_X1    g552(.A(new_n426), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n469), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n614), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n672), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n670), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n696), .B(new_n733), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n673), .A2(KEYINPUT117), .A3(new_n696), .A4(new_n733), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(G99gat), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n694), .A2(G99gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n741), .A2(new_n639), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT118), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n765), .A2(new_n770), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1338gat));
  AND2_X1   g571(.A1(new_n673), .A2(new_n733), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n424), .ZN(new_n774));
  INV_X1    g573(.A(G106gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n424), .A2(new_n775), .A3(new_n639), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT119), .Z(new_n777));
  AOI22_X1  g576(.A1(new_n774), .A2(G106gat), .B1(new_n741), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  INV_X1    g578(.A(new_n741), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n776), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n775), .B1(new_n773), .B2(new_n424), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n778), .A2(new_n779), .B1(new_n781), .B2(new_n782), .ZN(G1339gat));
  INV_X1    g582(.A(new_n674), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n616), .A2(new_n617), .A3(new_n710), .A4(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n628), .A2(new_n629), .A3(new_n624), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n636), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n633), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n630), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT55), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n788), .A2(new_n794), .A3(new_n791), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n793), .A2(new_n795), .B1(new_n626), .B2(new_n634), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n674), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT120), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n515), .A2(new_n519), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n517), .ZN(new_n800));
  AOI211_X1 g599(.A(KEYINPUT120), .B(new_n518), .C1(new_n515), .C2(new_n519), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n507), .A2(new_n508), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OAI221_X1 g602(.A(new_n639), .B1(new_n522), .B2(new_n529), .C1(new_n527), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n797), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n667), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n803), .A2(new_n527), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n522), .A2(new_n529), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n809), .B(new_n796), .C1(new_n665), .C2(new_n666), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n580), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n786), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n364), .ZN(new_n813));
  INV_X1    g612(.A(new_n466), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n537), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n674), .A2(new_n223), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n815), .B2(new_n817), .ZN(G1340gat));
  NOR2_X1   g617(.A1(new_n815), .A2(new_n710), .ZN(new_n819));
  MUX2_X1   g618(.A(G120gat), .B(new_n226), .S(new_n819), .Z(G1341gat));
  INV_X1    g619(.A(new_n815), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n580), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n758), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(G134gat), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT56), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(G134gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1343gat));
  INV_X1    g627(.A(new_n580), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n533), .A2(new_n536), .A3(new_n796), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n758), .B1(new_n830), .B2(new_n804), .ZN(new_n831));
  INV_X1    g630(.A(new_n810), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n785), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n425), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT121), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n424), .B1(new_n786), .B2(new_n811), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n835), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n834), .A2(new_n841), .A3(new_n836), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n696), .A2(new_n364), .A3(new_n397), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n674), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(G141gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n845), .B2(G141gat), .ZN(new_n848));
  INV_X1    g647(.A(new_n839), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n844), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(G141gat), .A3(new_n537), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n847), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  INV_X1    g652(.A(G141gat), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n843), .A2(new_n844), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n688), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n851), .A2(KEYINPUT58), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n852), .A2(new_n853), .B1(new_n856), .B2(new_n857), .ZN(G1344gat));
  INV_X1    g657(.A(new_n850), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n298), .A3(new_n639), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n839), .A2(KEYINPUT57), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n424), .A2(new_n835), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n640), .A2(new_n537), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n758), .A2(new_n796), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n758), .A2(new_n796), .A3(KEYINPUT124), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n867), .A2(new_n809), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n829), .B1(new_n869), .B2(new_n831), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n863), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT123), .B1(new_n862), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n836), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n812), .A2(KEYINPUT123), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n872), .A2(new_n639), .A3(new_n844), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n298), .B1(new_n876), .B2(KEYINPUT125), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n864), .A2(new_n870), .ZN(new_n878));
  OAI22_X1  g677(.A1(new_n878), .A2(new_n863), .B1(new_n849), .B2(new_n835), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n874), .B1(new_n879), .B2(KEYINPUT123), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n639), .A4(new_n844), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n861), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT59), .B(new_n298), .C1(new_n855), .C2(new_n639), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n860), .B1(new_n883), .B2(new_n884), .ZN(G1345gat));
  AOI21_X1  g684(.A(G155gat), .B1(new_n859), .B2(new_n580), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n829), .A2(new_n291), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n855), .B2(new_n887), .ZN(G1346gat));
  NAND3_X1  g687(.A1(new_n859), .A2(new_n292), .A3(new_n758), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n855), .A2(new_n668), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n292), .ZN(G1347gat));
  NOR3_X1   g690(.A1(new_n812), .A2(new_n424), .A3(new_n694), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n365), .A2(new_n465), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G169gat), .B1(new_n894), .B2(new_n537), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n784), .A2(G169gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(G1348gat));
  INV_X1    g696(.A(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n639), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n580), .A3(new_n210), .ZN(new_n901));
  NAND2_X1  g700(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n902));
  OAI21_X1  g701(.A(G183gat), .B1(new_n894), .B2(new_n829), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n904), .B(new_n905), .Z(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n894), .B2(new_n614), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT61), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n898), .A2(new_n211), .A3(new_n668), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1351gat));
  AND2_X1   g709(.A1(new_n288), .A2(new_n893), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n849), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(G197gat), .B1(new_n913), .B2(new_n674), .ZN(new_n914));
  INV_X1    g713(.A(new_n880), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n911), .B(KEYINPUT127), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n537), .A2(new_n524), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(G1352gat));
  NAND2_X1  g719(.A1(new_n880), .A2(new_n639), .ZN(new_n921));
  OAI21_X1  g720(.A(G204gat), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n912), .A2(G204gat), .A3(new_n710), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT62), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1353gat));
  OR3_X1    g724(.A1(new_n912), .A2(G211gat), .A3(new_n829), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n880), .A2(new_n580), .A3(new_n911), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1354gat));
  AOI21_X1  g729(.A(G218gat), .B1(new_n913), .B2(new_n668), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n758), .A2(G218gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n918), .B2(new_n932), .ZN(G1355gat));
endmodule


