

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741;

  XOR2_X1 U365 ( .A(KEYINPUT38), .B(n587), .Z(n645) );
  NAND2_X1 U366 ( .A1(n565), .A2(n474), .ZN(n456) );
  XNOR2_X1 U367 ( .A(n343), .B(KEYINPUT69), .ZN(n502) );
  INV_X2 U368 ( .A(G131), .ZN(n343) );
  AND2_X2 U369 ( .A1(n448), .A2(n362), .ZN(n447) );
  AND2_X2 U370 ( .A1(n738), .A2(KEYINPUT68), .ZN(n425) );
  XNOR2_X2 U371 ( .A(n570), .B(n455), .ZN(n564) );
  INV_X2 U372 ( .A(G143), .ZN(n459) );
  XNOR2_X2 U373 ( .A(n505), .B(n344), .ZN(n606) );
  XNOR2_X2 U374 ( .A(n706), .B(n358), .ZN(n344) );
  XNOR2_X2 U375 ( .A(n524), .B(n360), .ZN(n505) );
  XNOR2_X2 U376 ( .A(G116), .B(G119), .ZN(n419) );
  XNOR2_X2 U377 ( .A(n415), .B(G113), .ZN(n420) );
  NOR2_X1 U378 ( .A1(n735), .A2(n736), .ZN(n593) );
  XNOR2_X1 U379 ( .A(n432), .B(n430), .ZN(n657) );
  BUF_X1 U380 ( .A(G143), .Z(n405) );
  AND2_X1 U381 ( .A1(n394), .A2(n395), .ZN(n345) );
  INV_X2 U382 ( .A(KEYINPUT3), .ZN(n415) );
  XNOR2_X2 U383 ( .A(n531), .B(KEYINPUT80), .ZN(n536) );
  INV_X2 U384 ( .A(G953), .ZN(n730) );
  AND2_X1 U385 ( .A1(n346), .A2(n391), .ZN(n724) );
  NOR2_X1 U386 ( .A1(n345), .A2(n347), .ZN(n346) );
  NAND2_X1 U387 ( .A1(n356), .A2(n634), .ZN(n573) );
  NOR2_X1 U388 ( .A1(n543), .A2(n542), .ZN(n627) );
  OR2_X1 U389 ( .A1(n597), .A2(G902), .ZN(n355) );
  INV_X1 U390 ( .A(G475), .ZN(n354) );
  INV_X1 U391 ( .A(KEYINPUT76), .ZN(n350) );
  AND2_X1 U392 ( .A1(n396), .A2(n427), .ZN(n394) );
  OR2_X1 U393 ( .A1(n395), .A2(n427), .ZN(n349) );
  INV_X1 U394 ( .A(n642), .ZN(n348) );
  XNOR2_X1 U395 ( .A(n351), .B(n350), .ZN(n585) );
  XNOR2_X1 U396 ( .A(n377), .B(n376), .ZN(n740) );
  XNOR2_X1 U397 ( .A(n397), .B(n592), .ZN(n735) );
  NAND2_X1 U398 ( .A1(n575), .A2(KEYINPUT47), .ZN(n352) );
  AND2_X1 U399 ( .A1(n373), .A2(n365), .ZN(n375) );
  OR2_X1 U400 ( .A1(n677), .A2(n591), .ZN(n397) );
  XNOR2_X1 U401 ( .A(n378), .B(n374), .ZN(n373) );
  INV_X1 U402 ( .A(n627), .ZN(n637) );
  OR2_X1 U403 ( .A1(n385), .A2(n382), .ZN(n570) );
  XNOR2_X1 U404 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U405 ( .A(n355), .B(n353), .ZN(n542) );
  XNOR2_X1 U406 ( .A(n441), .B(n439), .ZN(n597) );
  XNOR2_X1 U407 ( .A(n359), .B(n476), .ZN(n358) );
  XNOR2_X1 U408 ( .A(n704), .B(KEYINPUT71), .ZN(n360) );
  XNOR2_X1 U409 ( .A(n465), .B(n466), .ZN(n359) );
  XNOR2_X1 U410 ( .A(n409), .B(G104), .ZN(n704) );
  XNOR2_X1 U411 ( .A(n485), .B(n354), .ZN(n353) );
  XNOR2_X1 U412 ( .A(G122), .B(KEYINPUT16), .ZN(n464) );
  XNOR2_X1 U413 ( .A(G146), .B(G125), .ZN(n476) );
  NAND2_X1 U414 ( .A1(n349), .A2(n348), .ZN(n347) );
  NAND2_X1 U415 ( .A1(n352), .A2(n737), .ZN(n351) );
  INV_X1 U416 ( .A(n594), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n627), .B(KEYINPUT98), .ZN(n594) );
  INV_X1 U418 ( .A(n573), .ZN(n649) );
  XNOR2_X2 U419 ( .A(n520), .B(n464), .ZN(n706) );
  XNOR2_X2 U420 ( .A(n420), .B(n419), .ZN(n520) );
  XNOR2_X2 U421 ( .A(n723), .B(n463), .ZN(n524) );
  XNOR2_X2 U422 ( .A(n399), .B(n462), .ZN(n723) );
  NAND2_X1 U423 ( .A1(n713), .A2(n724), .ZN(n403) );
  XNOR2_X1 U424 ( .A(n404), .B(n371), .ZN(n713) );
  XNOR2_X1 U425 ( .A(n578), .B(KEYINPUT6), .ZN(n555) );
  XNOR2_X1 U426 ( .A(n593), .B(KEYINPUT46), .ZN(n395) );
  XNOR2_X1 U427 ( .A(G140), .B(KEYINPUT10), .ZN(n477) );
  NAND2_X1 U428 ( .A1(G214), .A2(n467), .ZN(n644) );
  AND2_X1 U429 ( .A1(n657), .A2(n532), .ZN(n655) );
  NAND2_X1 U430 ( .A1(n387), .A2(n386), .ZN(n385) );
  NAND2_X1 U431 ( .A1(G469), .A2(G902), .ZN(n386) );
  XNOR2_X1 U432 ( .A(G478), .B(n496), .ZN(n543) );
  AND2_X1 U433 ( .A1(n586), .A2(n585), .ZN(n396) );
  XNOR2_X1 U434 ( .A(KEYINPUT67), .B(G101), .ZN(n463) );
  XNOR2_X1 U435 ( .A(n422), .B(n519), .ZN(n421) );
  XNOR2_X1 U436 ( .A(n522), .B(n518), .ZN(n422) );
  XNOR2_X1 U437 ( .A(G137), .B(KEYINPUT72), .ZN(n518) );
  XNOR2_X1 U438 ( .A(n502), .B(G134), .ZN(n720) );
  XNOR2_X1 U439 ( .A(n720), .B(n390), .ZN(n525) );
  INV_X1 U440 ( .A(G146), .ZN(n390) );
  XNOR2_X1 U441 ( .A(n527), .B(n526), .ZN(n578) );
  AND2_X1 U442 ( .A1(n392), .A2(n641), .ZN(n391) );
  NAND2_X1 U443 ( .A1(n549), .A2(n364), .ZN(n404) );
  XNOR2_X1 U444 ( .A(n510), .B(n429), .ZN(n428) );
  XNOR2_X1 U445 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n429) );
  XNOR2_X1 U446 ( .A(G134), .B(KEYINPUT95), .ZN(n488) );
  XNOR2_X1 U447 ( .A(n507), .B(n483), .ZN(n441) );
  XNOR2_X1 U448 ( .A(n482), .B(n440), .ZN(n439) );
  XNOR2_X1 U449 ( .A(n398), .B(n369), .ZN(n677) );
  NOR2_X1 U450 ( .A1(n648), .A2(n647), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n589), .B(n590), .ZN(n595) );
  NAND2_X1 U452 ( .A1(n556), .A2(n644), .ZN(n560) );
  XNOR2_X1 U453 ( .A(n436), .B(KEYINPUT100), .ZN(n556) );
  NOR2_X1 U454 ( .A1(n634), .A2(n437), .ZN(n436) );
  BUF_X1 U455 ( .A(n578), .Z(n661) );
  XNOR2_X1 U456 ( .A(n517), .B(n431), .ZN(n430) );
  OR2_X1 U457 ( .A1(n698), .A2(G902), .ZN(n432) );
  INV_X1 U458 ( .A(KEYINPUT25), .ZN(n431) );
  INV_X1 U459 ( .A(KEYINPUT1), .ZN(n455) );
  INV_X1 U460 ( .A(KEYINPUT22), .ZN(n374) );
  NOR2_X1 U461 ( .A1(n647), .A2(n413), .ZN(n412) );
  NOR2_X1 U462 ( .A1(G953), .A2(G237), .ZN(n521) );
  XNOR2_X1 U463 ( .A(n407), .B(KEYINPUT15), .ZN(n498) );
  XNOR2_X1 U464 ( .A(KEYINPUT84), .B(G902), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n501), .B(n500), .ZN(n658) );
  OR2_X1 U466 ( .A1(G902), .A2(G237), .ZN(n467) );
  NAND2_X1 U467 ( .A1(n506), .A2(n384), .ZN(n383) );
  INV_X1 U468 ( .A(G902), .ZN(n384) );
  INV_X1 U469 ( .A(KEYINPUT44), .ZN(n410) );
  XOR2_X1 U470 ( .A(KEYINPUT96), .B(G122), .Z(n487) );
  XNOR2_X1 U471 ( .A(G107), .B(G116), .ZN(n486) );
  XOR2_X1 U472 ( .A(KEYINPUT7), .B(KEYINPUT97), .Z(n489) );
  XNOR2_X1 U473 ( .A(n502), .B(n484), .ZN(n440) );
  XNOR2_X1 U474 ( .A(n405), .B(G104), .ZN(n484) );
  NAND2_X1 U475 ( .A1(n424), .A2(n361), .ZN(n450) );
  INV_X1 U476 ( .A(n532), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n421), .B(n418), .ZN(n523) );
  INV_X1 U478 ( .A(n520), .ZN(n418) );
  XNOR2_X1 U479 ( .A(G107), .B(G110), .ZN(n409) );
  XNOR2_X1 U480 ( .A(n504), .B(n505), .ZN(n685) );
  XNOR2_X1 U481 ( .A(n525), .B(n388), .ZN(n504) );
  XNOR2_X1 U482 ( .A(n389), .B(n508), .ZN(n388) );
  XNOR2_X1 U483 ( .A(n503), .B(G140), .ZN(n389) );
  NAND2_X1 U484 ( .A1(n446), .A2(n444), .ZN(n443) );
  NOR2_X1 U485 ( .A1(n445), .A2(n453), .ZN(n444) );
  NOR2_X1 U486 ( .A1(n582), .A2(n581), .ZN(n588) );
  XNOR2_X1 U487 ( .A(n579), .B(n381), .ZN(n380) );
  INV_X1 U488 ( .A(KEYINPUT30), .ZN(n381) );
  XNOR2_X1 U489 ( .A(n515), .B(n719), .ZN(n698) );
  XNOR2_X1 U490 ( .A(n511), .B(n428), .ZN(n514) );
  XNOR2_X1 U491 ( .A(n495), .B(n408), .ZN(n692) );
  XNOR2_X1 U492 ( .A(n599), .B(n598), .ZN(n600) );
  INV_X1 U493 ( .A(KEYINPUT75), .ZN(n402) );
  XNOR2_X1 U494 ( .A(n435), .B(n433), .ZN(n736) );
  XNOR2_X1 U495 ( .A(n434), .B(KEYINPUT40), .ZN(n433) );
  INV_X1 U496 ( .A(KEYINPUT104), .ZN(n434) );
  NOR2_X1 U497 ( .A1(n560), .A2(n577), .ZN(n562) );
  NOR2_X1 U498 ( .A1(n666), .A2(n401), .ZN(n541) );
  INV_X1 U499 ( .A(KEYINPUT99), .ZN(n376) );
  AND2_X1 U500 ( .A1(n373), .A2(n366), .ZN(n377) );
  NAND2_X1 U501 ( .A1(n543), .A2(n542), .ZN(n634) );
  INV_X1 U502 ( .A(n661), .ZN(n400) );
  NOR2_X1 U503 ( .A1(n555), .A2(n454), .ZN(n361) );
  OR2_X1 U504 ( .A1(n452), .A2(KEYINPUT34), .ZN(n362) );
  AND2_X1 U505 ( .A1(n547), .A2(n619), .ZN(n363) );
  AND2_X1 U506 ( .A1(n548), .A2(n363), .ZN(n364) );
  AND2_X1 U507 ( .A1(n555), .A2(n530), .ZN(n365) );
  NAND2_X1 U508 ( .A1(n555), .A2(n454), .ZN(n451) );
  NOR2_X1 U509 ( .A1(n654), .A2(n528), .ZN(n366) );
  AND2_X1 U510 ( .A1(n403), .A2(n402), .ZN(n367) );
  AND2_X1 U511 ( .A1(n450), .A2(n451), .ZN(n368) );
  INV_X1 U512 ( .A(n564), .ZN(n654) );
  XOR2_X1 U513 ( .A(KEYINPUT41), .B(KEYINPUT105), .Z(n369) );
  XOR2_X1 U514 ( .A(n475), .B(KEYINPUT0), .Z(n370) );
  INV_X1 U515 ( .A(KEYINPUT34), .ZN(n453) );
  XOR2_X1 U516 ( .A(KEYINPUT45), .B(KEYINPUT77), .Z(n371) );
  XOR2_X1 U517 ( .A(KEYINPUT78), .B(KEYINPUT35), .Z(n372) );
  AND2_X1 U518 ( .A1(n373), .A2(n564), .ZN(n545) );
  XNOR2_X1 U519 ( .A(n403), .B(KEYINPUT2), .ZN(n417) );
  XNOR2_X2 U520 ( .A(n375), .B(KEYINPUT32), .ZN(n739) );
  NAND2_X1 U521 ( .A1(n414), .A2(n412), .ZN(n378) );
  XNOR2_X1 U522 ( .A(n379), .B(n523), .ZN(n613) );
  XNOR2_X1 U523 ( .A(n524), .B(n525), .ZN(n379) );
  NAND2_X1 U524 ( .A1(n380), .A2(n580), .ZN(n581) );
  NOR2_X1 U525 ( .A1(n685), .A2(n383), .ZN(n382) );
  NAND2_X1 U526 ( .A1(n685), .A2(G469), .ZN(n387) );
  NAND2_X1 U527 ( .A1(n393), .A2(KEYINPUT48), .ZN(n392) );
  INV_X1 U528 ( .A(n396), .ZN(n393) );
  XNOR2_X1 U529 ( .A(n399), .B(KEYINPUT9), .ZN(n408) );
  NAND2_X2 U530 ( .A1(n461), .A2(n460), .ZN(n399) );
  AND2_X1 U531 ( .A1(n414), .A2(n451), .ZN(n423) );
  AND2_X1 U532 ( .A1(n414), .A2(n400), .ZN(n538) );
  INV_X1 U533 ( .A(n414), .ZN(n401) );
  XNOR2_X2 U534 ( .A(n456), .B(n370), .ZN(n414) );
  XNOR2_X2 U535 ( .A(n406), .B(KEYINPUT19), .ZN(n565) );
  NAND2_X1 U536 ( .A1(n559), .A2(n644), .ZN(n406) );
  NAND2_X1 U537 ( .A1(n595), .A2(n631), .ZN(n435) );
  NAND2_X1 U538 ( .A1(n450), .A2(n423), .ZN(n449) );
  XNOR2_X1 U539 ( .A(n411), .B(n410), .ZN(n549) );
  XNOR2_X2 U540 ( .A(n468), .B(n457), .ZN(n559) );
  NAND2_X1 U541 ( .A1(n536), .A2(n425), .ZN(n411) );
  NOR2_X2 U542 ( .A1(n740), .A2(n739), .ZN(n531) );
  XNOR2_X2 U543 ( .A(n416), .B(KEYINPUT65), .ZN(n691) );
  NAND2_X1 U544 ( .A1(n417), .A2(n596), .ZN(n416) );
  INV_X1 U545 ( .A(n540), .ZN(n424) );
  XNOR2_X2 U546 ( .A(n426), .B(n372), .ZN(n738) );
  NAND2_X1 U547 ( .A1(n535), .A2(n534), .ZN(n426) );
  INV_X1 U548 ( .A(KEYINPUT48), .ZN(n427) );
  INV_X1 U549 ( .A(n634), .ZN(n631) );
  NAND2_X1 U550 ( .A1(n438), .A2(n566), .ZN(n437) );
  INV_X1 U551 ( .A(n555), .ZN(n438) );
  NAND2_X1 U552 ( .A1(n447), .A2(n443), .ZN(n535) );
  INV_X1 U553 ( .A(n452), .ZN(n445) );
  INV_X1 U554 ( .A(n449), .ZN(n446) );
  NAND2_X1 U555 ( .A1(n449), .A2(n453), .ZN(n448) );
  NAND2_X1 U556 ( .A1(n368), .A2(n452), .ZN(n678) );
  NAND2_X1 U557 ( .A1(n540), .A2(n454), .ZN(n452) );
  INV_X1 U558 ( .A(KEYINPUT33), .ZN(n454) );
  NAND2_X1 U559 ( .A1(n603), .A2(n695), .ZN(n605) );
  XNOR2_X1 U560 ( .A(n601), .B(n600), .ZN(n603) );
  BUF_X1 U561 ( .A(n691), .Z(n699) );
  AND2_X1 U562 ( .A1(G210), .A2(n467), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n613), .B(n614), .ZN(n615) );
  XNOR2_X1 U564 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U565 ( .A(n694), .B(n693), .ZN(n696) );
  INV_X1 U566 ( .A(KEYINPUT60), .ZN(n604) );
  INV_X1 U567 ( .A(G128), .ZN(n458) );
  NAND2_X1 U568 ( .A1(n458), .A2(G143), .ZN(n461) );
  NAND2_X1 U569 ( .A1(n459), .A2(G128), .ZN(n460) );
  XNOR2_X2 U570 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n462) );
  NAND2_X1 U571 ( .A1(G224), .A2(n730), .ZN(n465) );
  XNOR2_X1 U572 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n466) );
  INV_X1 U573 ( .A(n498), .ZN(n596) );
  OR2_X2 U574 ( .A1(n606), .A2(n596), .ZN(n468) );
  NAND2_X1 U575 ( .A1(G237), .A2(G234), .ZN(n469) );
  XNOR2_X1 U576 ( .A(n469), .B(KEYINPUT14), .ZN(n471) );
  NAND2_X1 U577 ( .A1(G952), .A2(n471), .ZN(n675) );
  NOR2_X1 U578 ( .A1(n675), .A2(G953), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n470), .B(KEYINPUT85), .ZN(n553) );
  NAND2_X1 U580 ( .A1(G902), .A2(n471), .ZN(n550) );
  INV_X1 U581 ( .A(n550), .ZN(n472) );
  NOR2_X1 U582 ( .A1(G898), .A2(n730), .ZN(n707) );
  NAND2_X1 U583 ( .A1(n472), .A2(n707), .ZN(n473) );
  NAND2_X1 U584 ( .A1(n553), .A2(n473), .ZN(n474) );
  INV_X1 U585 ( .A(KEYINPUT81), .ZN(n475) );
  XNOR2_X1 U586 ( .A(KEYINPUT94), .B(KEYINPUT13), .ZN(n485) );
  XNOR2_X1 U587 ( .A(n477), .B(n476), .ZN(n507) );
  XOR2_X1 U588 ( .A(KEYINPUT93), .B(KEYINPUT11), .Z(n479) );
  XNOR2_X1 U589 ( .A(G122), .B(G113), .ZN(n478) );
  XNOR2_X1 U590 ( .A(n479), .B(n478), .ZN(n483) );
  XOR2_X1 U591 ( .A(KEYINPUT92), .B(KEYINPUT12), .Z(n481) );
  NAND2_X1 U592 ( .A1(n521), .A2(G214), .ZN(n480) );
  XNOR2_X1 U593 ( .A(n481), .B(n480), .ZN(n482) );
  INV_X1 U594 ( .A(n542), .ZN(n497) );
  XNOR2_X1 U595 ( .A(n487), .B(n486), .ZN(n491) );
  XNOR2_X1 U596 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U597 ( .A(n491), .B(n490), .Z(n494) );
  NAND2_X1 U598 ( .A1(G234), .A2(n730), .ZN(n492) );
  XOR2_X1 U599 ( .A(KEYINPUT8), .B(n492), .Z(n512) );
  NAND2_X1 U600 ( .A1(G217), .A2(n512), .ZN(n493) );
  XNOR2_X1 U601 ( .A(n494), .B(n493), .ZN(n495) );
  NOR2_X1 U602 ( .A1(n692), .A2(G902), .ZN(n496) );
  NAND2_X1 U603 ( .A1(n497), .A2(n543), .ZN(n647) );
  XOR2_X1 U604 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n501) );
  NAND2_X1 U605 ( .A1(G234), .A2(n498), .ZN(n499) );
  XNOR2_X1 U606 ( .A(KEYINPUT20), .B(n499), .ZN(n516) );
  NAND2_X1 U607 ( .A1(G221), .A2(n516), .ZN(n500) );
  XOR2_X1 U608 ( .A(KEYINPUT89), .B(n658), .Z(n532) );
  INV_X1 U609 ( .A(G469), .ZN(n506) );
  XOR2_X1 U610 ( .A(KEYINPUT70), .B(G137), .Z(n508) );
  NAND2_X1 U611 ( .A1(G227), .A2(n730), .ZN(n503) );
  XNOR2_X1 U612 ( .A(n508), .B(n507), .ZN(n719) );
  XNOR2_X1 U613 ( .A(G128), .B(G110), .ZN(n509) );
  XNOR2_X1 U614 ( .A(n509), .B(KEYINPUT87), .ZN(n511) );
  XNOR2_X1 U615 ( .A(G119), .B(KEYINPUT86), .ZN(n510) );
  NAND2_X1 U616 ( .A1(G221), .A2(n512), .ZN(n513) );
  XNOR2_X1 U617 ( .A(n514), .B(n513), .ZN(n515) );
  NAND2_X1 U618 ( .A1(n516), .A2(G217), .ZN(n517) );
  XOR2_X1 U619 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n519) );
  NAND2_X1 U620 ( .A1(n521), .A2(G210), .ZN(n522) );
  NOR2_X1 U621 ( .A1(G902), .A2(n613), .ZN(n527) );
  XNOR2_X1 U622 ( .A(KEYINPUT91), .B(G472), .ZN(n526) );
  OR2_X1 U623 ( .A1(n657), .A2(n661), .ZN(n528) );
  INV_X1 U624 ( .A(n657), .ZN(n529) );
  AND2_X1 U625 ( .A1(n529), .A2(n654), .ZN(n530) );
  NAND2_X1 U626 ( .A1(n655), .A2(n654), .ZN(n540) );
  INV_X1 U627 ( .A(n543), .ZN(n533) );
  NAND2_X1 U628 ( .A1(n533), .A2(n542), .ZN(n576) );
  XNOR2_X1 U629 ( .A(n576), .B(KEYINPUT73), .ZN(n534) );
  NOR2_X1 U630 ( .A1(n738), .A2(KEYINPUT68), .ZN(n537) );
  NAND2_X1 U631 ( .A1(n537), .A2(n536), .ZN(n548) );
  NAND2_X1 U632 ( .A1(n570), .A2(n655), .ZN(n582) );
  INV_X1 U633 ( .A(n582), .ZN(n539) );
  NAND2_X1 U634 ( .A1(n539), .A2(n538), .ZN(n622) );
  NAND2_X1 U635 ( .A1(n661), .A2(n424), .ZN(n666) );
  XNOR2_X1 U636 ( .A(KEYINPUT31), .B(n541), .ZN(n636) );
  NAND2_X1 U637 ( .A1(n622), .A2(n636), .ZN(n544) );
  NAND2_X1 U638 ( .A1(n544), .A2(n573), .ZN(n547) );
  AND2_X1 U639 ( .A1(n555), .A2(n545), .ZN(n546) );
  NAND2_X1 U640 ( .A1(n546), .A2(n657), .ZN(n619) );
  BUF_X2 U641 ( .A(n559), .Z(n587) );
  NOR2_X1 U642 ( .A1(G900), .A2(n550), .ZN(n551) );
  NAND2_X1 U643 ( .A1(G953), .A2(n551), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n553), .A2(n552), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n658), .A2(n580), .ZN(n554) );
  NOR2_X1 U646 ( .A1(n657), .A2(n554), .ZN(n566) );
  NOR2_X1 U647 ( .A1(n654), .A2(n560), .ZN(n557) );
  XNOR2_X1 U648 ( .A(n557), .B(KEYINPUT43), .ZN(n558) );
  NOR2_X1 U649 ( .A1(n587), .A2(n558), .ZN(n642) );
  INV_X1 U650 ( .A(n587), .ZN(n577) );
  XNOR2_X1 U651 ( .A(KEYINPUT107), .B(KEYINPUT36), .ZN(n561) );
  XNOR2_X1 U652 ( .A(n562), .B(n561), .ZN(n563) );
  NOR2_X1 U653 ( .A1(n564), .A2(n563), .ZN(n639) );
  INV_X1 U654 ( .A(n565), .ZN(n572) );
  NAND2_X1 U655 ( .A1(n661), .A2(n566), .ZN(n569) );
  XNOR2_X1 U656 ( .A(KEYINPUT28), .B(KEYINPUT103), .ZN(n567) );
  XNOR2_X1 U657 ( .A(n567), .B(KEYINPUT102), .ZN(n568) );
  XNOR2_X1 U658 ( .A(n569), .B(n568), .ZN(n571) );
  NAND2_X1 U659 ( .A1(n571), .A2(n570), .ZN(n591) );
  NOR2_X1 U660 ( .A1(n572), .A2(n591), .ZN(n632) );
  NAND2_X1 U661 ( .A1(n632), .A2(n573), .ZN(n575) );
  NOR2_X1 U662 ( .A1(KEYINPUT47), .A2(n575), .ZN(n574) );
  NOR2_X1 U663 ( .A1(n639), .A2(n574), .ZN(n586) );
  NOR2_X1 U664 ( .A1(n577), .A2(n576), .ZN(n583) );
  NAND2_X1 U665 ( .A1(n578), .A2(n644), .ZN(n579) );
  NAND2_X1 U666 ( .A1(n583), .A2(n588), .ZN(n584) );
  XOR2_X1 U667 ( .A(KEYINPUT101), .B(n584), .Z(n737) );
  XOR2_X1 U668 ( .A(KEYINPUT79), .B(KEYINPUT39), .Z(n590) );
  NAND2_X1 U669 ( .A1(n645), .A2(n588), .ZN(n589) );
  XOR2_X1 U670 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n592) );
  NAND2_X1 U671 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n641) );
  NAND2_X1 U673 ( .A1(n691), .A2(G475), .ZN(n601) );
  XOR2_X1 U674 ( .A(n597), .B(KEYINPUT82), .Z(n599) );
  XOR2_X1 U675 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n598) );
  NOR2_X1 U676 ( .A1(G952), .A2(n730), .ZN(n602) );
  XOR2_X1 U677 ( .A(KEYINPUT83), .B(n602), .Z(n703) );
  INV_X1 U678 ( .A(n703), .ZN(n695) );
  XNOR2_X1 U679 ( .A(n605), .B(n604), .ZN(G60) );
  NAND2_X1 U680 ( .A1(n691), .A2(G210), .ZN(n610) );
  XNOR2_X1 U681 ( .A(KEYINPUT55), .B(KEYINPUT74), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n606), .B(KEYINPUT54), .ZN(n607) );
  XNOR2_X1 U683 ( .A(n610), .B(n609), .ZN(n611) );
  AND2_X2 U684 ( .A1(n611), .A2(n695), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n612), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U686 ( .A1(n691), .A2(G472), .ZN(n616) );
  INV_X1 U687 ( .A(KEYINPUT62), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n617), .A2(n695), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U690 ( .A(G101), .B(n619), .ZN(G3) );
  NOR2_X1 U691 ( .A1(n634), .A2(n622), .ZN(n620) );
  XOR2_X1 U692 ( .A(KEYINPUT108), .B(n620), .Z(n621) );
  XNOR2_X1 U693 ( .A(G104), .B(n621), .ZN(G6) );
  NOR2_X1 U694 ( .A1(n622), .A2(n637), .ZN(n626) );
  XOR2_X1 U695 ( .A(KEYINPUT26), .B(KEYINPUT109), .Z(n624) );
  XNOR2_X1 U696 ( .A(G107), .B(KEYINPUT27), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n626), .B(n625), .ZN(G9) );
  XOR2_X1 U699 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n629) );
  NAND2_X1 U700 ( .A1(n632), .A2(n627), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(n630) );
  XOR2_X1 U702 ( .A(G128), .B(n630), .Z(G30) );
  NAND2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n633), .B(G146), .ZN(G48) );
  NOR2_X1 U705 ( .A1(n634), .A2(n636), .ZN(n635) );
  XOR2_X1 U706 ( .A(G113), .B(n635), .Z(G15) );
  NOR2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U708 ( .A(G116), .B(n638), .Z(G18) );
  XNOR2_X1 U709 ( .A(n639), .B(G125), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n640), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U711 ( .A(G134), .B(n641), .ZN(G36) );
  XOR2_X1 U712 ( .A(G140), .B(n642), .Z(n643) );
  XNOR2_X1 U713 ( .A(KEYINPUT112), .B(n643), .ZN(G42) );
  NOR2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n652) );
  NOR2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U717 ( .A(KEYINPUT115), .B(n650), .Z(n651) );
  NOR2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U719 ( .A1(n653), .A2(n678), .ZN(n671) );
  XNOR2_X1 U720 ( .A(KEYINPUT114), .B(KEYINPUT51), .ZN(n668) );
  NOR2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U722 ( .A(KEYINPUT50), .B(n656), .Z(n664) );
  NOR2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n660) );
  XNOR2_X1 U724 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n659) );
  XNOR2_X1 U725 ( .A(n660), .B(n659), .ZN(n662) );
  NOR2_X1 U726 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U727 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U728 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U729 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U730 ( .A1(n669), .A2(n677), .ZN(n670) );
  NOR2_X1 U731 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U732 ( .A(n672), .B(KEYINPUT116), .ZN(n673) );
  XNOR2_X1 U733 ( .A(KEYINPUT52), .B(n673), .ZN(n674) );
  NOR2_X1 U734 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U735 ( .A(n676), .B(KEYINPUT117), .ZN(n680) );
  OR2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U737 ( .A1(n680), .A2(n679), .ZN(n682) );
  XNOR2_X1 U738 ( .A(KEYINPUT2), .B(n367), .ZN(n681) );
  NOR2_X1 U739 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U740 ( .A1(n730), .A2(n683), .ZN(n684) );
  XOR2_X1 U741 ( .A(KEYINPUT53), .B(n684), .Z(G75) );
  XOR2_X1 U742 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n687) );
  XNOR2_X1 U743 ( .A(n685), .B(KEYINPUT118), .ZN(n686) );
  XNOR2_X1 U744 ( .A(n687), .B(n686), .ZN(n689) );
  NAND2_X1 U745 ( .A1(n699), .A2(G469), .ZN(n688) );
  XNOR2_X1 U746 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U747 ( .A1(n703), .A2(n690), .ZN(G54) );
  NAND2_X1 U748 ( .A1(G478), .A2(n691), .ZN(n694) );
  INV_X1 U749 ( .A(n692), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U751 ( .A(n697), .B(KEYINPUT119), .ZN(G63) );
  XNOR2_X1 U752 ( .A(n698), .B(KEYINPUT120), .ZN(n701) );
  NAND2_X1 U753 ( .A1(G217), .A2(n699), .ZN(n700) );
  XNOR2_X1 U754 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n703), .A2(n702), .ZN(G66) );
  XOR2_X1 U756 ( .A(n704), .B(G101), .Z(n705) );
  XNOR2_X1 U757 ( .A(n706), .B(n705), .ZN(n708) );
  NOR2_X1 U758 ( .A1(n708), .A2(n707), .ZN(n718) );
  XOR2_X1 U759 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n710) );
  NAND2_X1 U760 ( .A1(G224), .A2(G953), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U762 ( .A1(G898), .A2(n711), .ZN(n712) );
  XNOR2_X1 U763 ( .A(KEYINPUT122), .B(n712), .ZN(n716) );
  NAND2_X1 U764 ( .A1(n713), .A2(n730), .ZN(n714) );
  XOR2_X1 U765 ( .A(KEYINPUT123), .B(n714), .Z(n715) );
  NAND2_X1 U766 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(G69) );
  XNOR2_X1 U768 ( .A(n719), .B(KEYINPUT124), .ZN(n721) );
  XNOR2_X1 U769 ( .A(n720), .B(n721), .ZN(n722) );
  XOR2_X1 U770 ( .A(n723), .B(n722), .Z(n726) );
  XNOR2_X1 U771 ( .A(n724), .B(n726), .ZN(n725) );
  NOR2_X1 U772 ( .A1(G953), .A2(n725), .ZN(n733) );
  XNOR2_X1 U773 ( .A(G227), .B(n726), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n727), .A2(G900), .ZN(n728) );
  XNOR2_X1 U775 ( .A(KEYINPUT125), .B(n728), .ZN(n729) );
  NOR2_X1 U776 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U777 ( .A(n731), .B(KEYINPUT126), .ZN(n732) );
  NOR2_X1 U778 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U779 ( .A(KEYINPUT127), .B(n734), .ZN(G72) );
  XOR2_X1 U780 ( .A(G137), .B(n735), .Z(G39) );
  XOR2_X1 U781 ( .A(G131), .B(n736), .Z(G33) );
  XNOR2_X1 U782 ( .A(n737), .B(n405), .ZN(G45) );
  XNOR2_X1 U783 ( .A(n738), .B(G122), .ZN(G24) );
  XOR2_X1 U784 ( .A(n739), .B(G119), .Z(G21) );
  XOR2_X1 U785 ( .A(G110), .B(n740), .Z(n741) );
  XNOR2_X1 U786 ( .A(KEYINPUT110), .B(n741), .ZN(G12) );
endmodule

