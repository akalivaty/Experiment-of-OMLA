//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1272, new_n1273;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G125), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n469), .B2(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n463), .A2(G137), .A3(new_n465), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n463), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n465), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n467), .A2(new_n468), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(G136), .B2(new_n488), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT68), .Z(G162));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n465), .B2(G114), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G102), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(new_n465), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n492), .A2(new_n494), .A3(G2104), .A4(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n467), .B2(new_n468), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n501), .B(new_n504), .C1(new_n468), .C2(new_n467), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(G164));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n513), .A2(new_n514), .B1(new_n507), .B2(new_n508), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(new_n512), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI221_X1 g094(.A(new_n510), .B1(new_n511), .B2(new_n515), .C1(new_n518), .C2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n509), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n513), .A2(new_n514), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n509), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n526), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT70), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n534), .A2(new_n537), .A3(G651), .ZN(new_n538));
  INV_X1    g113(.A(new_n515), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n507), .A2(new_n508), .ZN(new_n540));
  INV_X1    g115(.A(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(G90), .A2(new_n539), .B1(new_n542), .B2(G52), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n536), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(new_n517), .A2(G56), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n519), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n549), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n524), .A2(new_n552), .B1(new_n553), .B2(new_n515), .ZN(new_n554));
  NOR3_X1   g129(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g132(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n558));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n524), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n542), .A2(new_n565), .A3(G53), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n562), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n564), .A2(new_n562), .A3(new_n566), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n527), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n539), .B2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  XNOR2_X1  g150(.A(new_n544), .B(KEYINPUT74), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n515), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n509), .A2(KEYINPUT75), .A3(G87), .A4(new_n517), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n580), .A2(new_n581), .B1(G49), .B2(new_n542), .ZN(new_n582));
  NOR3_X1   g157(.A1(new_n513), .A2(new_n514), .A3(G74), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT76), .B1(new_n583), .B2(new_n519), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n585), .B(G651), .C1(new_n517), .C2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n582), .A2(new_n587), .ZN(G288));
  OAI211_X1 g163(.A(G48), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n515), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n516), .B2(new_n512), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n539), .A2(G85), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n542), .A2(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n519), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n527), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n605), .B(KEYINPUT78), .C1(new_n606), .C2(new_n527), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(G651), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n515), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n612), .A2(new_n615), .B1(G54), .B2(new_n542), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G301), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G284));
  AOI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(new_n617), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  INV_X1    g203(.A(new_n555), .ZN(new_n629));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n617), .A2(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(new_n630), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n463), .A2(new_n476), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT13), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n482), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n465), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n488), .A2(new_n644), .A3(G135), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n488), .B2(G135), .ZN(new_n646));
  OAI221_X1 g221(.A(new_n641), .B1(new_n642), .B2(new_n643), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(G2096), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n639), .A2(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(G2096), .ZN(new_n650));
  NAND4_X1  g225(.A1(new_n640), .A2(new_n648), .A3(new_n649), .A4(new_n650), .ZN(G156));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2067), .B(G2678), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT81), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n669), .B(KEYINPUT17), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n671), .C1(new_n668), .C2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n668), .A3(new_n670), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  NOR2_X1   g272(.A1(G29), .A2(G35), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G162), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT29), .ZN(new_n700));
  INV_X1    g275(.A(G2090), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT91), .B(KEYINPUT25), .ZN(new_n703));
  AND3_X1   g278(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(G115), .A2(G2104), .ZN(new_n706));
  INV_X1    g281(.A(G127), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n487), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G2105), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n488), .A2(G139), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n705), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n714));
  OAI21_X1  g289(.A(G29), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G33), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(G29), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(new_n443), .ZN(new_n718));
  NAND2_X1  g293(.A1(G160), .A2(G29), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(KEYINPUT24), .A2(G34), .ZN(new_n721));
  NOR2_X1   g296(.A1(KEYINPUT24), .A2(G34), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT93), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n476), .A2(G105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT94), .ZN(new_n728));
  INV_X1    g303(.A(G141), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n463), .A2(new_n465), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT26), .Z(new_n733));
  INV_X1    g308(.A(G129), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n481), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(new_n720), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n720), .B2(G32), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n726), .A2(G2084), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n718), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(KEYINPUT95), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(KEYINPUT95), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n702), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n738), .A2(new_n739), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n720), .A2(G27), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G164), .B2(new_n720), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2078), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n749), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1966), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT31), .B(G11), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(G28), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n720), .B1(new_n754), .B2(G28), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n753), .B1(new_n755), .B2(new_n756), .C1(new_n647), .C2(new_n720), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n745), .A2(new_n748), .A3(new_n752), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n749), .A2(G4), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n626), .B2(new_n749), .ZN(new_n760));
  INV_X1    g335(.A(G1348), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n720), .A2(G26), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT28), .Z(new_n764));
  INV_X1    g339(.A(KEYINPUT88), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n488), .A2(new_n765), .A3(G140), .ZN(new_n766));
  INV_X1    g341(.A(G140), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT88), .B1(new_n730), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G128), .ZN(new_n770));
  OAI21_X1  g345(.A(KEYINPUT89), .B1(new_n481), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n463), .A2(new_n772), .A3(G128), .A4(G2105), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT90), .Z(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n769), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n764), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2067), .ZN(new_n780));
  NOR2_X1   g355(.A1(G5), .A2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT96), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n544), .B2(new_n749), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1961), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n758), .A2(new_n762), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n749), .A2(KEYINPUT82), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n749), .A2(KEYINPUT82), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT23), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n623), .B2(new_n749), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1956), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n789), .A2(G19), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n555), .B2(new_n789), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(G1341), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(G1341), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n726), .B2(G2084), .ZN(new_n798));
  OR4_X1    g373(.A1(new_n785), .A2(new_n793), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n744), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G23), .B(G288), .S(G16), .Z(new_n802));
  XOR2_X1   g377(.A(KEYINPUT33), .B(G1976), .Z(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n788), .A2(G22), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G166), .B2(new_n788), .ZN(new_n806));
  INV_X1    g381(.A(G1971), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n749), .A2(G6), .ZN(new_n809));
  INV_X1    g384(.A(G305), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n749), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT32), .B(G1981), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT84), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n811), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n802), .A2(new_n803), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n804), .A2(new_n808), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT85), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n789), .A2(G24), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT83), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G290), .B2(new_n788), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G1986), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n720), .A2(G25), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n463), .A2(G131), .A3(new_n465), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n463), .A2(G119), .A3(G2105), .ZN(new_n828));
  OR2_X1    g403(.A1(G95), .A2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n826), .B1(new_n832), .B2(new_n720), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G1991), .Z(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n820), .A2(new_n821), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT86), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n820), .A2(new_n841), .A3(new_n821), .A4(new_n837), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT87), .Z(new_n843));
  AOI21_X1  g418(.A(new_n801), .B1(new_n840), .B2(new_n843), .ZN(G311));
  INV_X1    g419(.A(KEYINPUT86), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n839), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n842), .B(KEYINPUT87), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n800), .B1(new_n846), .B2(new_n847), .ZN(G150));
  XOR2_X1   g423(.A(KEYINPUT98), .B(G860), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AOI22_X1  g425(.A1(G93), .A2(new_n539), .B1(new_n542), .B2(G55), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n519), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n629), .A2(KEYINPUT97), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(KEYINPUT97), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(KEYINPUT97), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n555), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT38), .Z(new_n859));
  NOR2_X1   g434(.A1(new_n617), .A2(new_n627), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n850), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n853), .A2(new_n850), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT100), .B1(new_n713), .B2(new_n714), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n712), .A3(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n503), .A2(new_n505), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n497), .A2(new_n498), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n769), .A2(new_n774), .A3(new_n777), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n736), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n778), .B1(new_n878), .B2(new_n877), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n882), .B1(new_n881), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n873), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n736), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n871), .B1(new_n870), .B2(new_n712), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n881), .A2(new_n883), .A3(new_n882), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n463), .A2(G142), .A3(new_n465), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n463), .A2(G130), .A3(G2105), .ZN(new_n894));
  OR2_X1    g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n895), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(new_n831), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n832), .A2(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT101), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n832), .A2(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n831), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n901), .A2(new_n637), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n637), .B1(new_n901), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n868), .B1(new_n892), .B2(new_n909), .ZN(new_n910));
  AOI211_X1 g485(.A(KEYINPUT102), .B(new_n908), .C1(new_n886), .C2(new_n891), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT103), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n884), .A2(new_n885), .A3(new_n869), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n869), .A2(new_n872), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(new_n888), .B2(new_n890), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n909), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT102), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n892), .A2(new_n868), .A3(new_n909), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n892), .A2(new_n909), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n912), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n647), .B(new_n479), .ZN(new_n924));
  XNOR2_X1  g499(.A(G162), .B(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n917), .A2(new_n919), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n921), .A2(new_n926), .ZN(new_n929));
  AOI21_X1  g504(.A(G37), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n927), .A2(KEYINPUT104), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT104), .B1(new_n927), .B2(new_n930), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n921), .B1(new_n928), .B2(KEYINPUT103), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n925), .B1(new_n936), .B2(new_n920), .ZN(new_n937));
  INV_X1    g512(.A(new_n930), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n927), .A2(KEYINPUT104), .A3(new_n930), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT40), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n934), .A2(new_n941), .ZN(G395));
  XNOR2_X1  g517(.A(G290), .B(KEYINPUT105), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(G288), .ZN(new_n944));
  XOR2_X1   g519(.A(G303), .B(G305), .Z(new_n945));
  XNOR2_X1  g520(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n947), .A2(KEYINPUT106), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(KEYINPUT106), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n950));
  OR3_X1    g525(.A1(new_n946), .A2(new_n950), .A3(KEYINPUT42), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n946), .B2(KEYINPUT42), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n948), .A2(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n858), .B(new_n632), .ZN(new_n954));
  XNOR2_X1  g529(.A(G299), .B(new_n617), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT41), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(G299), .B(new_n626), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT41), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n955), .B2(new_n954), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n953), .A2(KEYINPUT108), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n961), .A2(KEYINPUT108), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n961), .A2(KEYINPUT108), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n953), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n853), .A2(new_n630), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n967), .ZN(G331));
  NOR2_X1   g544(.A1(G301), .A2(G286), .ZN(new_n970));
  NOR2_X1   g545(.A1(G171), .A2(G168), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n858), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n854), .B(new_n857), .C1(new_n970), .C2(new_n971), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n958), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n973), .A2(new_n957), .A3(new_n959), .A4(new_n974), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n946), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G37), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n946), .B1(new_n976), .B2(new_n977), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n984), .B(new_n946), .C1(new_n976), .C2(new_n977), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n980), .B(new_n981), .C1(new_n983), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n978), .A2(new_n979), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT43), .B1(new_n987), .B2(new_n982), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n981), .B1(new_n987), .B2(new_n982), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n980), .B1(new_n983), .B2(new_n985), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(new_n981), .ZN(new_n992));
  MUX2_X1   g567(.A(new_n989), .B(new_n992), .S(KEYINPUT44), .Z(G397));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT110), .B1(new_n879), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n505), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n504), .B1(new_n463), .B2(new_n501), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n498), .B(new_n497), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT99), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(KEYINPUT110), .A3(new_n994), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n474), .A2(G40), .A3(new_n477), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n470), .A2(new_n471), .ZN(new_n1006));
  AOI211_X1 g581(.A(KEYINPUT67), .B(new_n465), .C1(new_n469), .C2(new_n461), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n995), .A2(new_n1003), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(G1986), .A3(G290), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G290), .A2(G1986), .ZN(new_n1011));
  XOR2_X1   g586(.A(new_n1011), .B(KEYINPUT111), .Z(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT112), .ZN(new_n1015));
  OR3_X1    g590(.A1(new_n995), .A2(new_n1003), .A3(new_n1008), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(G1996), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n736), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1009), .B(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g594(.A(G2067), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n880), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n778), .A2(G2067), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1996), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n736), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n831), .A2(new_n835), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n832), .A2(new_n834), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1019), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1015), .A2(new_n1018), .A3(new_n1026), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G2084), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1004), .B1(new_n466), .B2(new_n472), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n998), .A2(new_n1034), .A3(new_n994), .ZN(new_n1035));
  AND4_X1   g610(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT45), .B1(new_n998), .B2(new_n994), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT117), .B1(new_n1037), .B2(new_n1008), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1384), .B1(new_n874), .B2(new_n875), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1033), .B(new_n1039), .C1(KEYINPUT45), .C2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1002), .A2(G1384), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n998), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1966), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1036), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G286), .A2(G8), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT51), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1047), .B(new_n1051), .C1(new_n1046), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n1052), .B(new_n1051), .C1(new_n1046), .C2(G168), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1048), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT124), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n999), .A2(new_n1000), .A3(new_n1042), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1002), .B1(G164), .B2(G1384), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1058), .A2(new_n444), .A3(new_n1033), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  INV_X1    g636(.A(G1961), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1060), .A2(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1061), .A2(G2078), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1038), .A2(new_n1041), .A3(new_n1043), .A4(new_n1065), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n1057), .B(G301), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1063), .A2(new_n1062), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT124), .B1(new_n1070), .B2(new_n619), .ZN(new_n1071));
  NOR4_X1   g646(.A1(new_n1004), .A2(new_n470), .A3(new_n1061), .A4(G2078), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1058), .B(new_n1072), .C1(new_n995), .C2(new_n1003), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1073), .A2(new_n1064), .A3(G301), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1067), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1056), .B1(new_n1075), .B2(KEYINPUT54), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n510), .B1(new_n511), .B2(new_n515), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n518), .A2(new_n519), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT55), .B(G8), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1042), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n877), .A2(new_n878), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1033), .B1(new_n1040), .B2(KEYINPUT45), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n807), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1032), .A2(new_n701), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1052), .B(new_n1082), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n998), .A2(new_n994), .ZN(new_n1089));
  OAI21_X1  g664(.A(G8), .B1(new_n1008), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(G61), .B1(new_n513), .B2(new_n514), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n519), .B1(new_n1091), .B2(new_n595), .ZN(new_n1092));
  OAI21_X1  g667(.A(G1981), .B1(new_n591), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n509), .A2(G86), .A3(new_n517), .ZN(new_n1094));
  INV_X1    g669(.A(G1981), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n597), .A2(new_n1094), .A3(new_n1095), .A4(new_n589), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT49), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n1096), .A3(KEYINPUT49), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1093), .A2(new_n1096), .A3(new_n1101), .A4(KEYINPUT49), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1052), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n580), .A2(new_n581), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n542), .A2(G49), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1106), .A2(new_n587), .A3(G1976), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT114), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n582), .A2(KEYINPUT114), .A3(G1976), .A4(new_n587), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1105), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT52), .ZN(new_n1113));
  INV_X1    g688(.A(G1976), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT52), .B1(G288), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1115), .A2(new_n1110), .A3(new_n1105), .A4(new_n1111), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1104), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1088), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1034), .B1(new_n998), .B2(new_n994), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT116), .B1(new_n1120), .B2(new_n1008), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1033), .B(new_n1122), .C1(new_n1034), .C2(new_n1040), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(new_n701), .A3(new_n1123), .A4(new_n1035), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1086), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1082), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1118), .A2(new_n1119), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1082), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1037), .A2(new_n1008), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1971), .B1(new_n1130), .B2(new_n1058), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1087), .ZN(new_n1132));
  OAI211_X1 g707(.A(G8), .B(new_n1129), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(new_n1113), .A3(new_n1116), .A4(new_n1104), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1129), .B1(new_n1125), .B2(G8), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT125), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1064), .A2(G301), .A3(new_n1066), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1073), .A2(new_n1064), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT54), .B(new_n1137), .C1(new_n1138), .C2(new_n544), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1128), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT126), .B1(new_n1076), .B2(new_n1140), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1128), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1070), .A2(new_n619), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1057), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1070), .A2(KEYINPUT124), .A3(new_n619), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1073), .A2(new_n1064), .A3(G301), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1142), .A2(new_n1143), .A3(new_n1056), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1121), .A2(new_n1035), .A3(new_n1123), .ZN(new_n1152));
  INV_X1    g727(.A(G1956), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT56), .B(G2072), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1130), .A2(new_n1058), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n569), .ZN(new_n1158));
  OAI211_X1 g733(.A(KEYINPUT57), .B(new_n574), .C1(new_n1158), .C2(new_n567), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n564), .A2(new_n566), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT57), .B1(new_n1160), .B2(new_n574), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n570), .A2(new_n1162), .A3(KEYINPUT57), .A4(new_n574), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1157), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1154), .A2(new_n1164), .A3(new_n1165), .A4(new_n1156), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT61), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1058), .A2(new_n1024), .A3(new_n1033), .A4(new_n1059), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT58), .B(G1341), .Z(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1008), .B2(new_n1089), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT59), .B1(new_n1173), .B2(new_n555), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1175), .B(new_n629), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1063), .A2(new_n761), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1033), .A2(new_n1020), .A3(new_n1040), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(KEYINPUT60), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n611), .B2(new_n616), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT60), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1063), .A2(new_n761), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1179), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n617), .A2(KEYINPUT122), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1188), .A2(new_n1182), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1189), .A2(new_n1178), .A3(KEYINPUT60), .A4(new_n1179), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1183), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1177), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1169), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT121), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1167), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1157), .A2(KEYINPUT121), .A3(new_n1166), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1195), .A2(KEYINPUT61), .A3(new_n1196), .A4(new_n1168), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n626), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1195), .A2(new_n1198), .A3(new_n1196), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1193), .A2(new_n1197), .B1(new_n1199), .B2(new_n1168), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1141), .A2(new_n1151), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1117), .A2(new_n1133), .ZN(new_n1203));
  NOR2_X1   g778(.A1(G288), .A2(G1976), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1104), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1090), .B1(new_n1205), .B2(new_n1096), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1046), .A2(new_n1052), .A3(G286), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1208), .A2(KEYINPUT63), .A3(new_n1133), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(G8), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1211), .A2(new_n1082), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1117), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT119), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1129), .B1(new_n1210), .B2(G8), .ZN(new_n1216));
  OAI21_X1  g791(.A(KEYINPUT119), .B1(new_n1216), .B2(new_n1117), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1209), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g793(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1219), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1220), .B1(new_n1221), .B2(new_n1208), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1207), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1052), .B1(new_n1046), .B2(G168), .ZN(new_n1224));
  INV_X1    g799(.A(new_n1051), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1226), .A2(new_n1053), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1227), .A2(new_n1228), .A3(new_n1048), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1228), .B1(new_n1227), .B2(new_n1048), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1128), .A2(new_n1231), .A3(new_n1136), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1223), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g809(.A(new_n1030), .B1(new_n1202), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1026), .A2(new_n1018), .A3(new_n1027), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1236), .A2(new_n1021), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1237), .A2(new_n1019), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n1013), .B(KEYINPUT48), .ZN(new_n1239));
  NAND4_X1  g814(.A1(new_n1029), .A2(new_n1026), .A3(new_n1239), .A4(new_n1018), .ZN(new_n1240));
  XOR2_X1   g815(.A(new_n1017), .B(KEYINPUT46), .Z(new_n1241));
  INV_X1    g816(.A(KEYINPUT47), .ZN(new_n1242));
  INV_X1    g817(.A(new_n1023), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1019), .B1(new_n882), .B2(new_n1243), .ZN(new_n1244));
  AND3_X1   g819(.A1(new_n1241), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g820(.A(new_n1242), .B1(new_n1241), .B2(new_n1244), .ZN(new_n1246));
  OAI211_X1 g821(.A(new_n1238), .B(new_n1240), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g822(.A(KEYINPUT127), .B1(new_n1235), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g823(.A(KEYINPUT127), .ZN(new_n1249));
  INV_X1    g824(.A(new_n1247), .ZN(new_n1250));
  AND3_X1   g825(.A1(new_n1128), .A2(new_n1231), .A3(new_n1136), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1056), .A2(KEYINPUT62), .ZN(new_n1252));
  NAND3_X1  g827(.A1(new_n1251), .A2(new_n1252), .A3(new_n1229), .ZN(new_n1253));
  INV_X1    g828(.A(new_n1207), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1255));
  INV_X1    g830(.A(new_n1209), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1118), .A2(new_n1127), .ZN(new_n1258));
  INV_X1    g833(.A(new_n1208), .ZN(new_n1259));
  OAI21_X1  g834(.A(new_n1219), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g835(.A(new_n1254), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g836(.A1(new_n1253), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g837(.A(new_n1119), .B1(new_n1118), .B2(new_n1127), .ZN(new_n1263));
  NOR3_X1   g838(.A1(new_n1134), .A2(new_n1135), .A3(KEYINPUT125), .ZN(new_n1264));
  NOR2_X1   g839(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g840(.A1(new_n1265), .A2(new_n1139), .A3(new_n1150), .A4(new_n1056), .ZN(new_n1266));
  AOI21_X1  g841(.A(new_n1200), .B1(new_n1266), .B2(KEYINPUT126), .ZN(new_n1267));
  AOI21_X1  g842(.A(new_n1262), .B1(new_n1267), .B2(new_n1151), .ZN(new_n1268));
  OAI211_X1 g843(.A(new_n1249), .B(new_n1250), .C1(new_n1268), .C2(new_n1030), .ZN(new_n1269));
  NAND2_X1  g844(.A1(new_n1248), .A2(new_n1269), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g845(.A(G319), .ZN(new_n1272));
  NOR4_X1   g846(.A1(G229), .A2(new_n1272), .A3(G401), .A4(G227), .ZN(new_n1273));
  OAI211_X1 g847(.A(new_n989), .B(new_n1273), .C1(new_n931), .C2(new_n932), .ZN(G225));
  INV_X1    g848(.A(G225), .ZN(G308));
endmodule


