//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n592, new_n593, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n637, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT69), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n469), .A2(new_n470), .B1(new_n478), .B2(G2105), .ZN(G160));
  INV_X1    g054(.A(new_n465), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT71), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n475), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n482), .B(new_n485), .C1(G124), .C2(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(G126), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n463), .B2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT72), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n475), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OAI211_X1 g071(.A(KEYINPUT73), .B(new_n495), .C1(new_n465), .C2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(KEYINPUT73), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n475), .A2(new_n499), .A3(new_n461), .A4(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n494), .A2(new_n497), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT74), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT76), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n510), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n521), .B1(new_n508), .B2(new_n509), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OAI211_X1 g098(.A(G88), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n526));
  INV_X1    g101(.A(new_n523), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n515), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT75), .A3(G50), .ZN(new_n529));
  OAI211_X1 g104(.A(G50), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n525), .B1(new_n529), .B2(new_n532), .ZN(G166));
  XOR2_X1   g108(.A(KEYINPUT77), .B(G51), .Z(new_n534));
  NAND2_X1  g109(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n537), .A2(new_n538), .B1(new_n520), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n520), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n526), .B2(new_n527), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G89), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n543), .A2(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n528), .A2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n542), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(new_n510), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n542), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(new_n510), .ZN(new_n558));
  OAI211_X1 g133(.A(G43), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n559));
  OAI211_X1 g134(.A(G81), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT78), .ZN(new_n561));
  AOI21_X1  g136(.A(KEYINPUT78), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g140(.A(KEYINPUT79), .B(new_n558), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  OAI211_X1 g148(.A(G53), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n575), .A2(new_n576), .B1(G91), .B2(new_n543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  INV_X1    g153(.A(new_n517), .ZN(new_n579));
  NOR2_X1   g154(.A1(KEYINPUT5), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT80), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n516), .A2(new_n582), .A3(new_n517), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n578), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(G78), .A2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT81), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n588), .B(G651), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n577), .A2(new_n590), .ZN(G299));
  NAND2_X1  g166(.A1(new_n529), .A2(new_n532), .ZN(new_n592));
  INV_X1    g167(.A(new_n525), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G303));
  NAND2_X1  g169(.A1(new_n543), .A2(G87), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n528), .A2(G49), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(new_n543), .A2(G86), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n528), .A2(G48), .ZN(new_n602));
  INV_X1    g177(.A(G61), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n516), .B2(new_n517), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT82), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G73), .A2(G543), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n604), .B2(KEYINPUT82), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n510), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n543), .A2(KEYINPUT83), .A3(G86), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n601), .A2(new_n602), .A3(new_n609), .A4(new_n610), .ZN(G305));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n542), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n510), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT84), .ZN(new_n616));
  AOI22_X1  g191(.A1(G85), .A2(new_n543), .B1(new_n528), .B2(G47), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(G290));
  NAND2_X1  g193(.A1(G301), .A2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n543), .A2(G92), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT85), .B(KEYINPUT10), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT86), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n620), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n581), .A2(new_n583), .ZN(new_n625));
  INV_X1    g200(.A(G66), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n627), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n619), .B1(new_n630), .B2(G868), .ZN(G284));
  OAI21_X1  g206(.A(new_n619), .B1(new_n630), .B2(G868), .ZN(G321));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(G299), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(G168), .ZN(G297));
  OAI21_X1  g210(.A(new_n634), .B1(new_n633), .B2(G168), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n630), .B1(new_n637), .B2(G860), .ZN(G148));
  NAND2_X1  g213(.A1(new_n567), .A2(new_n633), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n629), .A2(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g217(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  INV_X1    g220(.A(G2100), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  OR2_X1    g223(.A1(G99), .A2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n649), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n650));
  INV_X1    g225(.A(G135), .ZN(new_n651));
  INV_X1    g226(.A(G123), .ZN(new_n652));
  OAI221_X1 g227(.A(new_n650), .B1(new_n465), .B2(new_n651), .C1(new_n486), .C2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n647), .A2(new_n648), .A3(new_n655), .ZN(G156));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT87), .Z(G401));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n646), .ZN(new_n680));
  XOR2_X1   g255(.A(G2072), .B(G2078), .Z(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n676), .B2(KEYINPUT18), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(new_n654), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n688), .A2(new_n689), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(new_n695), .B(new_n694), .S(new_n687), .Z(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1981), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT89), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(KEYINPUT24), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(G34), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(G34), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G160), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G29), .ZN(new_n710));
  INV_X1    g285(.A(G2084), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT99), .ZN(new_n714));
  INV_X1    g289(.A(G141), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n465), .ZN(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT26), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(KEYINPUT26), .ZN(new_n719));
  INV_X1    g294(.A(G129), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n718), .B(new_n719), .C1(new_n486), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT100), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  OR2_X1    g299(.A1(G29), .A2(G32), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n724), .A2(KEYINPUT101), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(KEYINPUT101), .B2(new_n724), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT27), .B(G1996), .Z(new_n728));
  AOI21_X1  g303(.A(new_n712), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G21), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G168), .B2(new_n730), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(G1966), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n729), .B1(KEYINPUT104), .B2(new_n733), .C1(new_n728), .C2(new_n727), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n736), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT105), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n733), .A2(KEYINPUT104), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G1348), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n630), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G4), .B2(G16), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n740), .B1(new_n741), .B2(new_n743), .C1(new_n735), .C2(new_n739), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n736), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n736), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT29), .Z(new_n748));
  INV_X1    g323(.A(G2090), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G171), .A2(new_n730), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G5), .B2(new_n730), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n752), .A2(new_n753), .B1(new_n732), .B2(G1966), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n750), .B(new_n754), .C1(new_n753), .C2(new_n752), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n736), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n480), .A2(G140), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT96), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n760));
  INV_X1    g335(.A(G116), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT97), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n487), .A2(G128), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n759), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT98), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n757), .B1(new_n767), .B2(new_n736), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2067), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n743), .A2(new_n741), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n736), .A2(G33), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT25), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n475), .A2(G127), .ZN(new_n774));
  NAND2_X1  g349(.A1(G115), .A2(G2104), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n461), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n773), .B(new_n776), .C1(G139), .C2(new_n480), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n771), .B1(new_n777), .B2(new_n736), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G2072), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(G2072), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n653), .A2(new_n736), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT103), .B(G28), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n782), .B2(KEYINPUT30), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(KEYINPUT30), .B2(new_n782), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT102), .B(KEYINPUT31), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G11), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n770), .B(new_n788), .C1(new_n748), .C2(new_n749), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n755), .A2(new_n769), .A3(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT92), .B(G16), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G20), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT23), .Z(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1956), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n745), .A2(new_n790), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n791), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(G19), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n568), .B2(new_n797), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G1341), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n791), .A2(G22), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT94), .Z(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G303), .B2(new_n797), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT95), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n730), .A2(G23), .ZN(new_n808));
  INV_X1    g383(.A(G288), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n730), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT33), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1976), .ZN(new_n812));
  MUX2_X1   g387(.A(G6), .B(G305), .S(G16), .Z(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n807), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n818));
  MUX2_X1   g393(.A(G24), .B(G290), .S(new_n797), .Z(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT93), .B(G1986), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n736), .A2(G25), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n480), .A2(G131), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT90), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n826));
  INV_X1    g401(.A(G107), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(G2105), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n487), .B2(G119), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n824), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n825), .B1(new_n824), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n822), .B1(new_n832), .B2(new_n736), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT35), .B(G1991), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n821), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n817), .A2(new_n818), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT36), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n817), .A2(new_n839), .A3(new_n818), .A4(new_n836), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n801), .B1(new_n838), .B2(new_n840), .ZN(G311));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n840), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n842), .A2(new_n800), .A3(new_n796), .ZN(G150));
  NAND2_X1  g418(.A1(new_n630), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n543), .A2(G93), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n528), .A2(G55), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n542), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n510), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n846), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n565), .A2(new_n566), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n563), .A2(new_n846), .A3(new_n847), .A4(new_n851), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT106), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n853), .A2(new_n857), .A3(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n845), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n845), .A2(new_n859), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n861), .B1(new_n860), .B2(new_n862), .ZN(new_n866));
  OR3_X1    g441(.A1(new_n865), .A2(KEYINPUT107), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT107), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n852), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(G145));
  INV_X1    g448(.A(new_n722), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n777), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n723), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n777), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n494), .A2(new_n503), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n497), .A2(KEYINPUT109), .A3(new_n501), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT109), .B1(new_n497), .B2(new_n501), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n480), .A2(G142), .ZN(new_n884));
  INV_X1    g459(.A(G130), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n461), .A2(G118), .ZN(new_n886));
  OAI21_X1  g461(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n887));
  OAI221_X1 g462(.A(new_n884), .B1(new_n885), .B2(new_n486), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n644), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n830), .B2(new_n831), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n832), .A2(new_n889), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n766), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n766), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n883), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  INV_X1    g472(.A(new_n883), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n878), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(G160), .B(new_n653), .Z(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(G162), .Z(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n896), .A2(new_n899), .A3(new_n878), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n903), .B1(new_n907), .B2(new_n900), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g486(.A1(new_n859), .A2(new_n640), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n856), .B(new_n858), .C1(G559), .C2(new_n629), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n623), .A2(new_n590), .A3(new_n577), .A4(new_n628), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n623), .A2(new_n628), .B1(new_n577), .B2(new_n590), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n629), .A2(G299), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(KEYINPUT41), .A3(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n913), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n919), .A2(KEYINPUT110), .A3(new_n915), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT110), .B1(new_n919), .B2(new_n915), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n912), .B2(new_n913), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT42), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n927), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n930), .A3(new_n922), .ZN(new_n931));
  XNOR2_X1  g506(.A(G290), .B(new_n809), .ZN(new_n932));
  XNOR2_X1  g507(.A(G305), .B(G303), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n928), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n928), .B2(new_n931), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n852), .A2(new_n633), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G295));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n938), .ZN(G331));
  OR2_X1    g515(.A1(G301), .A2(KEYINPUT111), .ZN(new_n941));
  NAND2_X1  g516(.A1(G301), .A2(KEYINPUT111), .ZN(new_n942));
  NAND3_X1  g517(.A1(G168), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(G286), .A2(KEYINPUT111), .A3(G301), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n853), .A2(new_n857), .A3(new_n854), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n857), .B1(new_n853), .B2(new_n854), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n944), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n856), .A2(new_n858), .A3(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n948), .A2(new_n950), .A3(new_n926), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n921), .B1(new_n948), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n934), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n921), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n946), .A2(new_n945), .A3(new_n947), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n949), .B1(new_n856), .B2(new_n858), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n934), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n916), .A2(new_n917), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n948), .A2(new_n950), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n953), .A2(new_n961), .A3(new_n909), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT112), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n953), .A2(new_n961), .A3(new_n964), .A4(new_n909), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(KEYINPUT43), .A3(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n948), .A2(new_n950), .A3(new_n959), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n934), .B1(new_n967), .B2(new_n952), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n968), .A2(new_n961), .A3(new_n969), .A4(new_n909), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n970), .A2(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n961), .A2(new_n909), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n969), .B1(new_n974), .B2(new_n968), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n972), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT45), .B1(new_n883), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G40), .ZN(new_n981));
  AOI221_X4 g556(.A(new_n981), .B1(new_n478), .B2(G2105), .C1(new_n469), .C2(new_n470), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n766), .B(G2067), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n874), .A2(G1996), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n876), .B2(G1996), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n832), .B(new_n834), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(G290), .B(G1986), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n984), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n504), .B2(new_n979), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT114), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n996));
  NAND3_X1  g571(.A1(new_n883), .A2(new_n979), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n995), .A2(new_n711), .A3(new_n982), .A4(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G1384), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n504), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n497), .A2(new_n501), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n497), .A2(KEYINPUT109), .A3(new_n501), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n1006), .B2(new_n880), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1001), .B(new_n982), .C1(new_n1007), .C2(KEYINPUT45), .ZN(new_n1008));
  INV_X1    g583(.A(G1966), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n998), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT118), .B(G8), .Z(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G168), .A2(new_n1012), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(KEYINPUT51), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n998), .B2(new_n1010), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT51), .B1(new_n1019), .B2(new_n1015), .ZN(new_n1020));
  AOI211_X1 g595(.A(G168), .B(new_n1012), .C1(new_n998), .C2(new_n1010), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT116), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G166), .A2(new_n1018), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT55), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n1026), .B2(KEYINPUT55), .ZN(new_n1030));
  NOR4_X1   g605(.A1(G166), .A2(KEYINPUT115), .A3(new_n1024), .A4(new_n1018), .ZN(new_n1031));
  OAI22_X1  g606(.A1(new_n1025), .A2(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT117), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n995), .A2(new_n749), .A3(new_n982), .A4(new_n997), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n883), .A2(new_n1000), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n999), .B1(G164), .B2(G1384), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n982), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n805), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1018), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT115), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1031), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1023), .A2(KEYINPUT116), .A3(new_n1024), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1027), .B1(new_n1026), .B2(KEYINPUT55), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1033), .A2(new_n1039), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1038), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n996), .B1(new_n883), .B2(new_n979), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n504), .A2(new_n993), .A3(new_n979), .ZN(new_n1051));
  NAND3_X1  g626(.A1(G160), .A2(new_n1051), .A3(G40), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1050), .A2(new_n1052), .A3(G2090), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1013), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  NOR2_X1   g631(.A1(G305), .A2(G1981), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n609), .A2(new_n602), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n599), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1056), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(new_n1058), .A3(new_n601), .A4(new_n610), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1059), .A2(new_n599), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT49), .B(new_n1062), .C1(new_n1063), .C2(new_n1058), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1012), .B1(new_n1007), .B2(new_n982), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1976), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT52), .B1(G288), .B2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1065), .B(new_n1068), .C1(new_n1067), .C2(G288), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n883), .A2(new_n979), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G160), .A2(G40), .ZN(new_n1071));
  OAI221_X1 g646(.A(new_n1013), .B1(new_n1067), .B2(G288), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1066), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1048), .A2(new_n1055), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n994), .A2(KEYINPUT114), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n1078), .B(new_n993), .C1(new_n504), .C2(new_n979), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n997), .B(new_n982), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT122), .B(G1961), .Z(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1035), .A2(new_n982), .A3(new_n1036), .A4(new_n735), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1070), .A2(new_n999), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n735), .A2(KEYINPUT53), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n982), .A3(new_n1001), .A4(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1082), .A2(G301), .A3(new_n1085), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT54), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1086), .A2(new_n982), .A3(new_n1035), .A4(new_n1088), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1082), .A2(new_n1085), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G301), .B1(new_n1093), .B2(KEYINPUT126), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1082), .A2(new_n1095), .A3(new_n1085), .A4(new_n1092), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1091), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1022), .A2(new_n1076), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1956), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT56), .B(G2072), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1035), .A2(new_n982), .A3(new_n1036), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n577), .A2(new_n590), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1100), .A2(new_n1102), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G2067), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1080), .A2(new_n741), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n629), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1100), .A2(new_n1103), .A3(new_n1105), .A4(new_n1102), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT61), .B1(new_n1106), .B2(KEYINPUT121), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1111), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1116), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n1111), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  INV_X1    g695(.A(G1996), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1035), .A2(new_n982), .A3(new_n1036), .A4(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1122), .A2(KEYINPUT120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1007), .A2(new_n982), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  AOI22_X1  g700(.A1(new_n1122), .A2(KEYINPUT120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1120), .B1(new_n1127), .B2(new_n568), .ZN(new_n1128));
  AOI211_X1 g703(.A(KEYINPUT59), .B(new_n567), .C1(new_n1123), .C2(new_n1126), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1118), .B(new_n1119), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1080), .A2(new_n741), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1108), .A2(new_n1107), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1131), .A2(new_n629), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT60), .B1(new_n1110), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1109), .A2(new_n1135), .A3(new_n630), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1112), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1082), .A2(G301), .A3(new_n1085), .A4(new_n1092), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1001), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n980), .A2(new_n1071), .A3(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1142), .A2(new_n1088), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1143));
  AOI21_X1  g718(.A(G301), .B1(new_n1143), .B2(new_n1082), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1139), .B2(KEYINPUT124), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT125), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1150));
  OAI21_X1  g725(.A(G171), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(KEYINPUT124), .A3(new_n1139), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1146), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1148), .A2(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1098), .A2(new_n1138), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1065), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n809), .A2(new_n1067), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT119), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1057), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n1048), .A2(new_n1074), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g738(.A(G286), .B(new_n1012), .C1(new_n998), .C2(new_n1010), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1048), .A2(new_n1055), .A3(new_n1075), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT63), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1014), .A2(new_n1166), .A3(G286), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1039), .A2(new_n1032), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1168), .A2(new_n1048), .A3(new_n1075), .A4(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1163), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1022), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1076), .A2(new_n1151), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1017), .B(KEYINPUT62), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n992), .B1(new_n1157), .B2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n988), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n767), .A2(new_n1107), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n983), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OR3_X1    g757(.A1(new_n983), .A2(G1986), .A3(G290), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n990), .A2(new_n984), .B1(KEYINPUT48), .B2(new_n1184), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1184), .A2(KEYINPUT48), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1182), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n984), .B1(new_n985), .B2(new_n874), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n984), .A2(new_n1121), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT46), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT47), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1188), .A2(KEYINPUT47), .A3(new_n1190), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1193), .A2(KEYINPUT127), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1187), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT127), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1178), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(G319), .ZN(new_n1201));
  NOR4_X1   g775(.A1(G229), .A2(new_n1201), .A3(new_n671), .A4(G227), .ZN(new_n1202));
  OAI211_X1 g776(.A(new_n910), .B(new_n1202), .C1(new_n975), .C2(new_n976), .ZN(G225));
  INV_X1    g777(.A(G225), .ZN(G308));
endmodule


