//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT64), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  OAI22_X1  g047(.A1(new_n462), .A2(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n473), .A2(new_n476), .ZN(G160));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  OR3_X1    g053(.A1(new_n469), .A2(KEYINPUT65), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n464), .A2(new_n466), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n468), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT65), .B1(new_n469), .B2(new_n478), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n479), .A2(new_n482), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT4), .B1(new_n469), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n480), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(new_n491), .A3(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n481), .A2(G126), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(KEYINPUT6), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT66), .A3(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT67), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT68), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  AND2_X1   g091(.A1(G75), .A2(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n515), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n505), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n507), .A2(new_n522), .A3(G50), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n510), .A2(new_n518), .A3(new_n521), .A4(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  AND2_X1   g100(.A1(new_n503), .A2(new_n504), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(G89), .A3(new_n515), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n503), .A2(G51), .A3(G543), .A4(new_n504), .ZN(new_n528));
  AND3_X1   g103(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT5), .B1(KEYINPUT68), .B2(G543), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT69), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n513), .A2(new_n532), .A3(new_n514), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  AND4_X1   g112(.A1(new_n527), .A2(new_n528), .A3(new_n535), .A4(new_n537), .ZN(G168));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n531), .B2(new_n533), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(G651), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n503), .A2(new_n515), .A3(G90), .A4(new_n504), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n503), .A2(G52), .A3(G543), .A4(new_n504), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n546), .B1(new_n544), .B2(new_n545), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n507), .A2(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n526), .A2(new_n515), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n534), .A2(G56), .ZN(new_n555));
  AND2_X1   g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n499), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  AOI22_X1  g140(.A1(new_n507), .A2(G53), .B1(KEYINPUT71), .B2(KEYINPUT9), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  AND4_X1   g142(.A1(KEYINPUT71), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n515), .B2(G91), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n567), .A2(new_n499), .B1(new_n569), .B2(new_n505), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n549), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g148(.A(KEYINPUT72), .B(new_n543), .C1(new_n547), .C2(new_n548), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G301));
  NAND4_X1  g150(.A1(new_n527), .A2(new_n528), .A3(new_n535), .A4(new_n537), .ZN(G286));
  NAND2_X1  g151(.A1(new_n520), .A2(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n507), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n507), .A2(G48), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n520), .A2(G86), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n515), .A2(G61), .ZN(new_n583));
  AND2_X1   g158(.A1(G73), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(KEYINPUT73), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(KEYINPUT73), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n588), .A2(G651), .A3(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(G47), .A2(new_n507), .B1(new_n520), .B2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n553), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n519), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(G54), .A2(new_n507), .B1(new_n597), .B2(G651), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT10), .B1(new_n553), .B2(new_n593), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G301), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G284));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  XNOR2_X1  g183(.A(G280), .B(KEYINPUT74), .ZN(G297));
  INV_X1    g184(.A(new_n600), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  NOR2_X1   g187(.A1(new_n600), .A2(G559), .ZN(new_n613));
  OR3_X1    g188(.A1(new_n613), .A2(KEYINPUT75), .A3(new_n601), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT75), .B1(new_n613), .B2(new_n601), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n614), .B(new_n615), .C1(G868), .C2(new_n559), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XOR2_X1   g192(.A(new_n470), .B(KEYINPUT64), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n467), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n621), .A2(KEYINPUT77), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT76), .B(G2100), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n481), .A2(G123), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n490), .A2(G135), .ZN(new_n627));
  OR2_X1    g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n628), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n621), .A2(KEYINPUT77), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n624), .B(new_n632), .C1(new_n625), .C2(new_n631), .ZN(G156));
  XOR2_X1   g208(.A(KEYINPUT15), .B(G2435), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT78), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT14), .ZN(new_n639));
  XOR2_X1   g214(.A(G2443), .B(G2446), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G14), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT79), .Z(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT80), .Z(new_n655));
  XOR2_X1   g230(.A(new_n653), .B(KEYINPUT17), .Z(new_n656));
  OAI21_X1  g231(.A(new_n655), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n653), .A3(new_n649), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n651), .A3(new_n649), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2096), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(KEYINPUT81), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(KEYINPUT81), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n665), .A2(new_n666), .ZN(new_n675));
  AOI22_X1  g250(.A1(new_n673), .A2(new_n674), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n671), .A2(new_n667), .A3(new_n675), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n676), .B(new_n677), .C1(new_n674), .C2(new_n673), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  INV_X1    g256(.A(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n680), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G22), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n686), .A2(G16), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G303), .B2(G16), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n687), .B(new_n688), .S(KEYINPUT85), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1971), .ZN(new_n690));
  NOR2_X1   g265(.A1(G16), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(G16), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G6), .ZN(new_n697));
  INV_X1    g272(.A(G305), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT84), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n690), .A2(new_n695), .A3(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT34), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n481), .A2(G119), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n490), .A2(G131), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n468), .A2(G107), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n706), .B(new_n707), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT82), .ZN(new_n711));
  MUX2_X1   g286(.A(G25), .B(new_n711), .S(G29), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G24), .ZN(new_n715));
  INV_X1    g290(.A(G290), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G16), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT83), .B(G1986), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n704), .A2(new_n705), .A3(new_n714), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT36), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(G26), .ZN(new_n723));
  AOI22_X1  g298(.A1(G128), .A2(new_n481), .B1(new_n490), .B2(G140), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n725));
  NOR2_X1   g300(.A1(G104), .A2(G2105), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT86), .Z(new_n727));
  OAI21_X1  g302(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n723), .B1(new_n728), .B2(G29), .ZN(new_n729));
  MUX2_X1   g304(.A(new_n723), .B(new_n729), .S(KEYINPUT28), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2067), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n559), .A2(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G16), .B2(G19), .ZN(new_n733));
  INV_X1    g308(.A(G1341), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(G171), .A2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G5), .B2(G16), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(G29), .A2(G32), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n618), .A2(G105), .B1(G129), .B2(new_n481), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n490), .A2(G141), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT26), .Z(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(new_n722), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G2084), .ZN(new_n749));
  AND2_X1   g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  NOR2_X1   g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n750), .A2(new_n751), .A3(G29), .ZN(new_n752));
  INV_X1    g327(.A(G160), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G29), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n748), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT89), .Z(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G21), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G168), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1966), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n490), .A2(G139), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n761), .B(new_n762), .C1(new_n763), .C2(new_n468), .ZN(new_n764));
  MUX2_X1   g339(.A(G33), .B(new_n764), .S(G29), .Z(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G2072), .Z(new_n766));
  AND2_X1   g341(.A1(KEYINPUT30), .A2(G28), .ZN(new_n767));
  NOR2_X1   g342(.A1(KEYINPUT30), .A2(G28), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n722), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n769), .B(new_n770), .C1(new_n630), .C2(new_n722), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT88), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n766), .B(new_n772), .C1(new_n733), .C2(new_n734), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n722), .A2(G35), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G162), .B2(new_n722), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT29), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n759), .B(new_n773), .C1(G2090), .C2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n696), .A2(KEYINPUT23), .A3(G20), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT23), .ZN(new_n779));
  INV_X1    g354(.A(G20), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(G16), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n778), .B(new_n781), .C1(new_n607), .C2(new_n696), .ZN(new_n782));
  INV_X1    g357(.A(G1956), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G2090), .B2(new_n776), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n746), .A2(new_n747), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT87), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n749), .B2(new_n754), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n696), .A2(G4), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n610), .B2(new_n696), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1348), .ZN(new_n791));
  NOR2_X1   g366(.A1(G164), .A2(new_n722), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G27), .B2(new_n722), .ZN(new_n793));
  INV_X1    g368(.A(G2078), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n793), .A2(new_n794), .B1(new_n737), .B2(new_n738), .ZN(new_n795));
  NOR4_X1   g370(.A1(new_n785), .A2(new_n788), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n756), .A2(new_n777), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n721), .A2(new_n731), .A3(new_n735), .A4(new_n797), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n793), .A2(new_n794), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(G311));
  INV_X1    g375(.A(G311), .ZN(G150));
  AND2_X1   g376(.A1(new_n534), .A2(G67), .ZN(new_n802));
  NAND2_X1  g377(.A1(G80), .A2(G543), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(G651), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT90), .B(G55), .ZN(new_n806));
  AOI22_X1  g381(.A1(G93), .A2(new_n520), .B1(new_n507), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT92), .B(G860), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n610), .A2(G559), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT39), .ZN(new_n814));
  INV_X1    g389(.A(new_n558), .ZN(new_n815));
  AOI22_X1  g390(.A1(G43), .A2(new_n507), .B1(new_n520), .B2(G81), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n808), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n805), .B(new_n807), .C1(new_n554), .C2(new_n558), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n814), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n812), .B1(new_n822), .B2(new_n809), .ZN(G145));
  XNOR2_X1  g398(.A(G160), .B(new_n630), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G162), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n489), .A2(new_n492), .B1(G126), .B2(new_n481), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(new_n495), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n728), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n745), .B(new_n764), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n481), .A2(G130), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n490), .A2(G142), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n468), .A2(G118), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n620), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n711), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n830), .A2(new_n837), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n838), .B1(new_n841), .B2(KEYINPUT95), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n839), .B(KEYINPUT94), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n825), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  INV_X1    g422(.A(new_n825), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n841), .A2(new_n848), .A3(new_n838), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g426(.A1(new_n808), .A2(new_n601), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n692), .A2(new_n698), .ZN(new_n853));
  NAND2_X1  g428(.A1(G288), .A2(G305), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n716), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(G290), .A2(new_n854), .A3(new_n853), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n856), .A2(G166), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(G166), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT96), .Z(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT97), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n600), .B(G299), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT41), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n819), .B(new_n613), .ZN(new_n869));
  MUX2_X1   g444(.A(new_n867), .B(new_n868), .S(new_n869), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n865), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n852), .B1(new_n871), .B2(new_n601), .ZN(G295));
  OAI21_X1  g447(.A(new_n852), .B1(new_n871), .B2(new_n601), .ZN(G331));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n817), .A2(new_n818), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n549), .B2(G168), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(G301), .B2(G168), .ZN(new_n880));
  AOI211_X1 g455(.A(new_n878), .B(G286), .C1(new_n573), .C2(new_n574), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n544), .A2(new_n545), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT70), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT72), .B1(new_n886), .B2(new_n543), .ZN(new_n887));
  INV_X1    g462(.A(new_n574), .ZN(new_n888));
  OAI211_X1 g463(.A(KEYINPUT99), .B(G168), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G286), .B1(new_n573), .B2(new_n574), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n889), .B(new_n819), .C1(new_n890), .C2(new_n879), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n876), .B1(new_n882), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n891), .A2(new_n876), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n875), .B1(new_n894), .B2(new_n868), .ZN(new_n895));
  NOR4_X1   g470(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT101), .A4(new_n866), .ZN(new_n896));
  INV_X1    g471(.A(new_n891), .ZN(new_n897));
  OAI21_X1  g472(.A(G168), .B1(new_n887), .B2(new_n888), .ZN(new_n898));
  INV_X1    g473(.A(new_n879), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n819), .B1(new_n900), .B2(new_n889), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n866), .B(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n895), .A2(new_n896), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n847), .B1(new_n906), .B2(new_n860), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT102), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT100), .B1(new_n897), .B2(new_n901), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n891), .A2(new_n876), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n868), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT101), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n894), .A2(new_n875), .A3(new_n868), .ZN(new_n913));
  INV_X1    g488(.A(new_n905), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n860), .A4(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(KEYINPUT98), .B(KEYINPUT43), .Z(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n918), .B(new_n847), .C1(new_n906), .C2(new_n860), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n908), .A2(new_n915), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n860), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n897), .A2(new_n901), .A3(new_n866), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n921), .B(new_n922), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n847), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n867), .B1(new_n892), .B2(new_n893), .ZN(new_n927));
  INV_X1    g502(.A(new_n924), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n860), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(new_n922), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n915), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n874), .B1(new_n920), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n931), .A2(new_n935), .A3(new_n915), .A4(new_n917), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n929), .B2(new_n922), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT103), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n937), .A2(new_n939), .A3(new_n915), .A4(new_n917), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT104), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n908), .A2(new_n915), .A3(new_n919), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n916), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n934), .B1(new_n944), .B2(new_n874), .ZN(G397));
  NOR2_X1   g520(.A1(G290), .A2(G1986), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n948));
  NAND2_X1  g523(.A1(G290), .A2(G1986), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n826), .B2(new_n495), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n951), .A2(KEYINPUT105), .ZN(new_n952));
  XOR2_X1   g527(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(KEYINPUT105), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G160), .A2(G40), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n950), .B(new_n958), .C1(new_n948), .C2(new_n949), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT108), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n745), .B(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G2067), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n728), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n711), .B(new_n713), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n958), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT109), .ZN(new_n969));
  INV_X1    g544(.A(G1976), .ZN(new_n970));
  AND2_X1   g545(.A1(G160), .A2(G40), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n951), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G8), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n698), .A2(new_n682), .ZN(new_n975));
  NAND2_X1  g550(.A1(G305), .A2(G1981), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT49), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n977), .A2(KEYINPUT111), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT111), .B1(new_n977), .B2(new_n978), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n974), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n975), .A2(KEYINPUT49), .A3(new_n976), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT112), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n970), .B(new_n692), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n984), .A2(new_n975), .ZN(new_n985));
  NAND2_X1  g560(.A1(G303), .A2(G8), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT55), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n957), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n954), .B1(G164), .B2(G1384), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(KEYINPUT110), .A3(new_n990), .ZN(new_n994));
  AOI21_X1  g569(.A(G1971), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n951), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n998), .A3(new_n971), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G2090), .ZN(new_n1000));
  OAI211_X1 g575(.A(G8), .B(new_n988), .C1(new_n995), .C2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G288), .A2(new_n970), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT52), .B1(new_n973), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(G288), .B2(new_n970), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n974), .B(new_n1004), .C1(new_n970), .C2(G288), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1003), .B(new_n1005), .C1(new_n981), .C2(new_n983), .ZN(new_n1006));
  OAI22_X1  g581(.A1(new_n985), .A2(new_n973), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(G8), .B1(new_n995), .B2(new_n1000), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n987), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1006), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n1001), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n999), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n749), .ZN(new_n1014));
  INV_X1    g589(.A(G1966), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n971), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n1016));
  AOI211_X1 g591(.A(G1384), .B(new_n954), .C1(new_n826), .C2(new_n495), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n1015), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1014), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(G8), .A3(G168), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT114), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1012), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT63), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(KEYINPUT115), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1012), .B(new_n1024), .C1(new_n1028), .C2(KEYINPUT63), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1007), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(G2072), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n989), .A2(new_n990), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT117), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n989), .A2(new_n1035), .A3(new_n990), .A4(new_n1032), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n1038));
  XNOR2_X1  g613(.A(G299), .B(KEYINPUT57), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n999), .A2(new_n783), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(new_n1041), .A3(new_n1036), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT118), .B1(new_n1043), .B2(new_n1039), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g620(.A1(new_n1013), .A2(G1348), .B1(G2067), .B2(new_n972), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1046), .A2(new_n610), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1043), .A2(new_n1039), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(KEYINPUT119), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1043), .A2(new_n1053), .A3(new_n1039), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1052), .A2(new_n1042), .A3(new_n1044), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1051), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1046), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1037), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1059), .A2(KEYINPUT61), .A3(new_n1049), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1055), .A2(new_n1051), .A3(new_n1056), .ZN(new_n1062));
  INV_X1    g637(.A(new_n972), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT58), .B(G1341), .ZN(new_n1064));
  OAI22_X1  g639(.A1(new_n991), .A2(G1996), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n559), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT59), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1046), .A2(new_n610), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT60), .B1(new_n1047), .B2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1062), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1050), .B1(new_n1061), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1011), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1009), .A2(new_n1010), .A3(KEYINPUT124), .A4(new_n1001), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1014), .A2(new_n1019), .A3(G168), .A4(new_n1021), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT121), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1022), .A2(G8), .A3(G286), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1077), .A2(new_n1083), .A3(new_n1078), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n993), .A2(new_n794), .A3(new_n994), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n999), .A2(new_n738), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1088), .A2(G2078), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n956), .A2(new_n989), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT123), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n956), .A2(new_n1097), .A3(new_n989), .A4(new_n1094), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1092), .A2(G301), .A3(new_n1093), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT122), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1094), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1102), .A2(new_n1093), .A3(new_n1089), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n603), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1100), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1092), .A2(G301), .A3(new_n1093), .A4(new_n1104), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1102), .A2(new_n1093), .A3(new_n1089), .A4(new_n1099), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G171), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1107), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1075), .B(new_n1085), .C1(new_n1108), .C2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1030), .B1(new_n1071), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1106), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1081), .A2(new_n1117), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT125), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1115), .A2(new_n1116), .A3(new_n1121), .A4(new_n1118), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n969), .B1(new_n1114), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT46), .ZN(new_n1125));
  INV_X1    g700(.A(new_n958), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(G1996), .ZN(new_n1127));
  INV_X1    g702(.A(new_n964), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n958), .B1(new_n745), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n958), .A2(KEYINPUT46), .A3(new_n961), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT47), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n958), .A2(new_n946), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT127), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT48), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1135), .A2(new_n967), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n713), .B(new_n711), .C1(new_n958), .C2(new_n965), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n728), .A2(G2067), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT126), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1132), .B(new_n1136), .C1(new_n958), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1124), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g717(.A1(G229), .A2(new_n460), .ZN(new_n1144));
  INV_X1    g718(.A(new_n1144), .ZN(new_n1145));
  AOI21_X1  g719(.A(G227), .B1(new_n646), .B2(G14), .ZN(new_n1146));
  NAND2_X1  g720(.A1(new_n850), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g721(.A1(new_n943), .A2(new_n916), .ZN(new_n1148));
  AND2_X1   g722(.A1(new_n936), .A2(new_n941), .ZN(new_n1149));
  AOI211_X1 g723(.A(new_n1145), .B(new_n1147), .C1(new_n1148), .C2(new_n1149), .ZN(G308));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  INV_X1    g725(.A(new_n1147), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n1151), .A2(new_n1144), .A3(new_n1152), .ZN(G225));
endmodule


