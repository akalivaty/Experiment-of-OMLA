//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n466));
  OAI211_X1 g041(.A(new_n462), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT66), .B(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n469), .A2(new_n473), .ZN(G160));
  OAI221_X1 g049(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n462), .A2(new_n464), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT67), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n475), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n478), .A2(new_n480), .ZN(new_n486));
  INV_X1    g061(.A(new_n470), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT68), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n486), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n485), .B1(new_n492), .B2(G124), .ZN(G162));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n476), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n460), .A2(G102), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n479), .A2(new_n470), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n499), .B1(new_n467), .B2(new_n500), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n497), .A2(new_n498), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n511), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n506), .A2(new_n512), .B1(new_n513), .B2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND2_X1  g094(.A1(new_n511), .A2(new_n516), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT70), .B(G89), .ZN(new_n521));
  AND3_X1   g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n520), .A2(new_n521), .B1(KEYINPUT7), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n511), .A2(G63), .ZN(new_n524));
  NAND3_X1  g099(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n506), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n516), .A2(KEYINPUT69), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n514), .A2(new_n529), .A3(new_n515), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n528), .A2(G543), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n527), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n506), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n528), .A2(G543), .A3(new_n530), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n520), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n540), .A2(KEYINPUT71), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(KEYINPUT71), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g120(.A(KEYINPUT72), .B(new_n536), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n508), .A2(new_n510), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G651), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  OAI221_X1 g129(.A(new_n552), .B1(new_n553), .B2(new_n520), .C1(new_n537), .C2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n528), .A2(G53), .A3(G543), .A4(new_n530), .ZN(new_n563));
  NOR2_X1   g138(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(new_n520), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n563), .A2(new_n564), .B1(new_n565), .B2(G91), .ZN(new_n566));
  XOR2_X1   g141(.A(KEYINPUT73), .B(KEYINPUT9), .Z(new_n567));
  NAND3_X1  g142(.A1(new_n531), .A2(G53), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n549), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT74), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n571), .A2(new_n574), .A3(G651), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n566), .A2(new_n568), .A3(new_n573), .A4(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  OAI21_X1  g152(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n511), .A2(G87), .A3(new_n516), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n528), .A2(G49), .A3(G543), .A4(new_n530), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  AND2_X1   g158(.A1(new_n516), .A2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n549), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(G543), .A2(new_n584), .B1(new_n587), .B2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n565), .A2(G86), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n549), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n565), .A2(G85), .B1(new_n593), .B2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n531), .A2(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n531), .A2(KEYINPUT75), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT75), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n537), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(G54), .A3(new_n600), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n511), .A2(G92), .A3(new_n516), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(new_n506), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n601), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT76), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n597), .B1(G868), .B2(new_n607), .ZN(G284));
  XOR2_X1   g183(.A(G284), .B(KEYINPUT77), .Z(G321));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g185(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n607), .B1(new_n612), .B2(G860), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT79), .Z(G148));
  OAI21_X1  g189(.A(KEYINPUT80), .B1(new_n556), .B2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n612), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  MUX2_X1   g192(.A(KEYINPUT80), .B(new_n615), .S(new_n617), .Z(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g194(.A(G123), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n489), .B2(new_n491), .ZN(new_n621));
  OAI221_X1 g196(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n622));
  INV_X1    g197(.A(G135), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n483), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2096), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n479), .A2(new_n460), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2100), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n626), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2435), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2438), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2443), .B(G2446), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2451), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT83), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n647), .A2(G14), .A3(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n651), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n653), .A2(new_n654), .ZN(new_n660));
  AOI21_X1  g235(.A(KEYINPUT18), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n658), .B(new_n661), .Z(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  INV_X1    g246(.A(new_n668), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n671), .B1(new_n664), .B2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT22), .B(G1981), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  INV_X1    g259(.A(G34), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n685), .A2(KEYINPUT24), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(KEYINPUT24), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G160), .B2(new_n684), .ZN(new_n689));
  INV_X1    g264(.A(G2084), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(G28), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(G28), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n694), .A3(new_n684), .ZN(new_n695));
  INV_X1    g270(.A(G2072), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G29), .B2(G33), .ZN(new_n698));
  OR3_X1    g273(.A1(new_n697), .A2(G29), .A3(G33), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n482), .A2(G139), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(new_n470), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n698), .B(new_n699), .C1(new_n706), .C2(new_n684), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n691), .B(new_n695), .C1(new_n696), .C2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G27), .A2(G29), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G164), .B2(G29), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n708), .B1(G2078), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G5), .A2(G16), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G171), .B2(G16), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G1961), .Z(new_n715));
  NAND2_X1  g290(.A1(G299), .A2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n717), .A2(KEYINPUT23), .A3(G20), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n719));
  INV_X1    g294(.A(G20), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G16), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n716), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT98), .B(G1956), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n715), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n482), .A2(G131), .ZN(new_n726));
  OAI221_X1 g301(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n492), .B2(G119), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(new_n684), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G25), .B2(new_n684), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT35), .B(G1991), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n732), .B(new_n730), .C1(G25), .C2(new_n684), .ZN(new_n735));
  MUX2_X1   g310(.A(G24), .B(G290), .S(G16), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1986), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  OR2_X1    g313(.A1(G16), .A2(G23), .ZN(new_n739));
  AOI21_X1  g314(.A(KEYINPUT87), .B1(new_n581), .B2(new_n582), .ZN(new_n740));
  INV_X1    g315(.A(new_n582), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n741), .A2(new_n580), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n739), .B1(new_n744), .B2(new_n717), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT33), .B(G1976), .Z(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n717), .A2(G22), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G166), .B2(new_n717), .ZN(new_n750));
  INV_X1    g325(.A(G1971), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n746), .B(new_n739), .C1(new_n744), .C2(new_n717), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n748), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT32), .B(G1981), .Z(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n717), .A2(G6), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G305), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n758), .A2(new_n759), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n758), .A2(new_n759), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n764), .A2(new_n755), .A3(new_n760), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n754), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(KEYINPUT34), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(KEYINPUT34), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n738), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(KEYINPUT88), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n738), .B1(KEYINPUT88), .B2(new_n771), .C1(new_n768), .C2(new_n769), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n712), .B(new_n725), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT31), .B(G11), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n707), .A2(new_n696), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n710), .A2(G2078), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n717), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n717), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1966), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n780), .B(new_n783), .C1(G29), .C2(new_n625), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n775), .A2(new_n776), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n460), .A2(G105), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT26), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n482), .B2(G141), .ZN(new_n789));
  AOI21_X1  g364(.A(KEYINPUT95), .B1(new_n492), .B2(G129), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n791));
  INV_X1    g366(.A(G129), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n489), .C2(new_n491), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n786), .B(new_n789), .C1(new_n790), .C2(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(KEYINPUT96), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(KEYINPUT96), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G32), .B(new_n797), .S(G29), .Z(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT27), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G1996), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(KEYINPUT27), .ZN(new_n801));
  INV_X1    g376(.A(G1996), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G35), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT97), .B1(new_n805), .B2(G29), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n805), .A2(KEYINPUT97), .A3(G29), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n806), .B(new_n807), .C1(G162), .C2(new_n684), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT29), .B(G2090), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G4), .A2(G16), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n607), .B2(G16), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1348), .Z(new_n813));
  INV_X1    g388(.A(KEYINPUT28), .ZN(new_n814));
  INV_X1    g389(.A(G26), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(G29), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(G29), .ZN(new_n817));
  OAI221_X1 g392(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT90), .Z(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n492), .B2(G128), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n482), .A2(G140), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT89), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n817), .B1(new_n823), .B2(G29), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n816), .B1(new_n824), .B2(new_n814), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(G2067), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(G2067), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n717), .A2(G19), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n556), .B2(new_n717), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(G1341), .Z(new_n830));
  NAND4_X1  g405(.A1(new_n813), .A2(new_n826), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT91), .Z(new_n832));
  NOR4_X1   g407(.A1(new_n785), .A2(new_n804), .A3(new_n810), .A4(new_n832), .ZN(G311));
  INV_X1    g408(.A(new_n785), .ZN(new_n834));
  INV_X1    g409(.A(new_n810), .ZN(new_n835));
  INV_X1    g410(.A(new_n832), .ZN(new_n836));
  INV_X1    g411(.A(new_n804), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(G150));
  AOI22_X1  g413(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT99), .B(G93), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n839), .A2(new_n506), .B1(new_n520), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n537), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n556), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n841), .A2(new_n843), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n555), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n607), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n846), .B1(new_n854), .B2(G860), .ZN(G145));
  NAND3_X1  g430(.A1(new_n820), .A2(new_n822), .A3(G164), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(G164), .B1(new_n820), .B2(new_n822), .ZN(new_n858));
  OAI21_X1  g433(.A(KEYINPUT100), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n823), .A2(new_n504), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n861), .A3(new_n856), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n797), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n706), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n859), .B(new_n862), .C1(new_n795), .C2(new_n796), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n794), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n860), .A3(new_n856), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n794), .B1(new_n857), .B2(new_n858), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n706), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(KEYINPUT101), .A3(new_n706), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n867), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(G160), .B1(new_n621), .B2(new_n624), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G162), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n621), .A2(G160), .A3(new_n624), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n479), .A2(new_n470), .A3(G137), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n479), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n461), .B(new_n882), .C1(new_n883), .C2(new_n470), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n625), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(G162), .B1(new_n885), .B2(new_n877), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n629), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  OAI221_X1 g462(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n470), .C2(G118), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n482), .A2(G142), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT102), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n492), .A2(new_n891), .A3(G130), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n492), .B2(G130), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n888), .B(new_n890), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n729), .ZN(new_n896));
  INV_X1    g471(.A(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n892), .ZN(new_n898));
  INV_X1    g473(.A(new_n729), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n888), .A4(new_n890), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(new_n902));
  INV_X1    g477(.A(new_n629), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n885), .A2(G162), .A3(new_n877), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n887), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n901), .B1(new_n887), .B2(new_n905), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n876), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n906), .A2(new_n907), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n910), .A2(new_n867), .A3(new_n874), .A4(new_n875), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n909), .A2(new_n911), .A3(KEYINPUT104), .A4(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT40), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(G395));
  OR2_X1    g496(.A1(new_n606), .A2(G299), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n606), .A2(G299), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n922), .A2(KEYINPUT41), .A3(new_n923), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT41), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n850), .B(KEYINPUT105), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(new_n616), .ZN(new_n929));
  MUX2_X1   g504(.A(new_n924), .B(new_n927), .S(new_n929), .Z(new_n930));
  NAND3_X1  g505(.A1(new_n581), .A2(KEYINPUT87), .A3(new_n582), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n742), .B1(new_n741), .B2(new_n580), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(G290), .B(G303), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G305), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n934), .A2(G305), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n937), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n935), .A3(new_n744), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n941), .B(KEYINPUT42), .Z(new_n942));
  XNOR2_X1  g517(.A(new_n930), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(G868), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g520(.A(new_n944), .B1(G868), .B2(new_n848), .ZN(G331));
  NAND3_X1  g521(.A1(G286), .A2(new_n847), .A3(new_n849), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(G286), .B1(new_n847), .B2(new_n849), .ZN(new_n949));
  OAI21_X1  g524(.A(G171), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n850), .A2(G168), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(new_n546), .A3(new_n545), .A4(new_n947), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n924), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n950), .B(new_n952), .C1(new_n926), .C2(new_n925), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n941), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n955), .A3(new_n941), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n912), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n954), .A2(new_n955), .A3(new_n941), .A4(KEYINPUT107), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n958), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n963), .B1(new_n969), .B2(new_n962), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n965), .A2(new_n967), .A3(new_n958), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT108), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n965), .A2(new_n975), .A3(new_n967), .A4(new_n958), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n966), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n960), .A2(new_n966), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT44), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n979), .ZN(G397));
  INV_X1    g555(.A(G2067), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n823), .B(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n983));
  INV_X1    g558(.A(G40), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n884), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  INV_X1    g563(.A(new_n494), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n479), .B2(G126), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n498), .B(new_n502), .C1(new_n990), .C2(new_n481), .ZN(new_n991));
  INV_X1    g566(.A(new_n503), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n982), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n998), .B(KEYINPUT111), .Z(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n794), .B2(new_n802), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n797), .B2(new_n802), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n899), .A2(new_n732), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n729), .A2(new_n733), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n996), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  OR3_X1    g581(.A1(new_n997), .A2(G1986), .A3(G290), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n996), .A2(G1986), .A3(G290), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT110), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT45), .B1(new_n504), .B2(new_n988), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT117), .B1(new_n987), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n995), .A2(new_n1015), .A3(new_n985), .A4(new_n986), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1966), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n993), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n504), .A2(KEYINPUT50), .A3(new_n988), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n987), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n690), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1012), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT114), .B(G8), .Z(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G168), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT51), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT120), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1032), .B(KEYINPUT51), .C1(new_n1026), .C2(new_n1029), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1018), .A2(new_n1019), .B1(new_n690), .B2(new_n1024), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(new_n1028), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1029), .A2(KEYINPUT51), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1034), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT121), .B(new_n1037), .C1(new_n1035), .C2(new_n1028), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1031), .A2(new_n1033), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1036), .A2(G286), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT126), .B1(new_n1043), .B2(KEYINPUT62), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT126), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT62), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1045), .B(new_n1046), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1041), .A2(new_n1046), .A3(new_n1042), .ZN(new_n1048));
  NAND3_X1  g623(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT112), .B(KEYINPUT113), .Z(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(G166), .B2(new_n1012), .ZN(new_n1054));
  NAND4_X1  g629(.A1(G303), .A2(KEYINPUT55), .A3(G8), .A4(new_n1050), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2090), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1024), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n995), .A2(new_n1017), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n1061));
  NOR4_X1   g636(.A1(new_n469), .A2(new_n473), .A3(new_n983), .A4(new_n984), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1971), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(G8), .B(new_n1056), .C1(new_n1059), .C2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(G1976), .B1(new_n740), .B2(new_n743), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT115), .ZN(new_n1067));
  INV_X1    g642(.A(new_n993), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1028), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n933), .A2(new_n1070), .A3(G1976), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT116), .B(G86), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n588), .B1(new_n520), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G1981), .ZN(new_n1075));
  INV_X1    g650(.A(G1981), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n588), .A2(new_n1076), .A3(new_n589), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1075), .A2(KEYINPUT49), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT49), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g655(.A1(KEYINPUT52), .A2(new_n1072), .B1(new_n1080), .B2(new_n1069), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1056), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1063), .A2(new_n1017), .A3(new_n995), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1024), .A2(new_n1057), .B1(new_n1083), .B2(new_n751), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1084), .B2(new_n1028), .ZN(new_n1085));
  INV_X1    g660(.A(G1976), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .A4(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1065), .A2(new_n1081), .A3(new_n1085), .A4(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1024), .A2(G1961), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1083), .B2(G2078), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1091), .A2(G2078), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1090), .B(new_n1092), .C1(new_n1093), .C2(new_n1018), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT123), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1097), .A3(G171), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1089), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1048), .A2(new_n1099), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1044), .A2(new_n1047), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1080), .A2(new_n1069), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n1088), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n1065), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n987), .A2(new_n993), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1103), .A2(new_n1086), .A3(new_n582), .A4(new_n581), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1106), .B(new_n1028), .C1(new_n1107), .C2(new_n1077), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1036), .A2(G168), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT118), .B1(new_n1089), .B2(new_n1109), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1084), .A2(new_n1012), .A3(new_n1082), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1104), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1035), .A2(G286), .A3(new_n1028), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1085), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1110), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(G8), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1116), .B1(new_n1118), .B2(new_n1082), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1112), .A2(new_n1119), .A3(new_n1114), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1105), .B(new_n1108), .C1(new_n1117), .C2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT58), .B(G1341), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1083), .A2(G1996), .B1(new_n1106), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n556), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT59), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1126), .A3(new_n556), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n1129));
  XNOR2_X1  g704(.A(G299), .B(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT56), .B(G2072), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1063), .A2(new_n1017), .A3(new_n995), .A4(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1130), .B(new_n1132), .C1(G1956), .C2(new_n1024), .ZN(new_n1133));
  XNOR2_X1  g708(.A(G299), .B(KEYINPUT57), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1135));
  AOI21_X1  g710(.A(G1956), .B1(new_n1135), .B2(new_n1063), .ZN(new_n1136));
  AND4_X1   g711(.A1(new_n1063), .A2(new_n1017), .A3(new_n995), .A4(new_n1131), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1133), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1128), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1128), .B(KEYINPUT119), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1106), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n1146), .A2(G2067), .B1(new_n1024), .B2(G1348), .ZN(new_n1147));
  OR3_X1    g722(.A1(new_n1147), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1147), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1149), .A2(new_n606), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n606), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT60), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1144), .A2(new_n1145), .A3(new_n1148), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1133), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1153), .A2(new_n1154), .A3(new_n1138), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1094), .A2(G171), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1156), .A2(KEYINPUT54), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n884), .A2(new_n984), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1093), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1060), .B(new_n1160), .C1(new_n1159), .C2(new_n1158), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1090), .A2(new_n1092), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(G171), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1089), .B1(new_n1157), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1162), .A2(G171), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1043), .A2(new_n1166), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1121), .B1(new_n1155), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1011), .B1(new_n1101), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n820), .A2(new_n822), .A3(new_n981), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n997), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1007), .B(KEYINPUT48), .Z(new_n1177));
  NOR2_X1   g752(.A1(new_n1006), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n802), .B1(KEYINPUT127), .B2(KEYINPUT46), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n982), .A2(new_n868), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n996), .A2(new_n802), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT127), .B(KEYINPUT46), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1180), .A2(new_n996), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT47), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1176), .A2(new_n1178), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1173), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g761(.A(G227), .ZN(new_n1188));
  INV_X1    g762(.A(G319), .ZN(new_n1189));
  NOR3_X1   g763(.A1(G401), .A2(new_n1189), .A3(G229), .ZN(new_n1190));
  AND4_X1   g764(.A1(new_n1188), .A2(new_n970), .A3(new_n917), .A4(new_n1190), .ZN(G308));
  NAND4_X1  g765(.A1(new_n970), .A2(new_n917), .A3(new_n1188), .A4(new_n1190), .ZN(G225));
endmodule


