// Benchmark "locked_c1355" written by ABC on Sat Dec 16 10:33:26 2023

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138, new_n139, new_n140, new_n141, new_n142, new_n143, new_n144,
    new_n145, new_n146, new_n147, new_n148, new_n149, new_n150, new_n151,
    new_n152, new_n153, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n138));
  INV_X1    g001(.A(KEYINPUT34), .ZN(new_n139));
  NAND2_X1  g002(.A1(G227gat), .A2(G233gat), .ZN(new_n140));
  INV_X1    g003(.A(new_n140), .ZN(new_n141));
  INV_X1    g004(.A(G113gat), .ZN(new_n142));
  INV_X1    g005(.A(G120gat), .ZN(new_n143));
  NAND2_X1  g006(.A1(new_n142), .A2(new_n143), .ZN(new_n144));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n145));
  NAND2_X1  g008(.A1(G113gat), .A2(G120gat), .ZN(new_n146));
  NAND3_X1  g009(.A1(new_n144), .A2(new_n145), .A3(new_n146), .ZN(new_n147));
  XNOR2_X1  g010(.A(G127gat), .B(G134gat), .ZN(new_n148));
  XNOR2_X1  g011(.A(new_n147), .B(new_n148), .ZN(new_n149));
  INV_X1    g012(.A(G190gat), .ZN(new_n150));
  AND2_X1   g013(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n151));
  NOR2_X1   g014(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n152));
  OAI21_X1  g015(.A(new_n150), .B1(new_n151), .B2(new_n152), .ZN(new_n153));
  NAND2_X1  g016(.A1(new_n153), .A2(KEYINPUT28), .ZN(new_n154));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n155));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n156));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n157));
  NAND2_X1  g020(.A1(new_n156), .A2(new_n157), .ZN(new_n158));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n159));
  OAI21_X1  g022(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n160));
  NAND3_X1  g023(.A1(new_n158), .A2(new_n159), .A3(new_n160), .ZN(new_n161));
  INV_X1    g024(.A(KEYINPUT28), .ZN(new_n162));
  OAI211_X1 g025(.A(new_n162), .B(new_n150), .C1(new_n151), .C2(new_n152), .ZN(new_n163));
  NAND4_X1  g026(.A1(new_n154), .A2(new_n155), .A3(new_n161), .A4(new_n163), .ZN(new_n164));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n165));
  INV_X1    g028(.A(G169gat), .ZN(new_n166));
  INV_X1    g029(.A(G176gat), .ZN(new_n167));
  NAND3_X1  g030(.A1(new_n165), .A2(new_n166), .A3(new_n167), .ZN(new_n168));
  NAND2_X1  g031(.A1(new_n159), .A2(KEYINPUT23), .ZN(new_n169));
  OAI21_X1  g032(.A(new_n168), .B1(new_n169), .B2(new_n156), .ZN(new_n170));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n171));
  NAND2_X1  g034(.A1(new_n155), .A2(new_n171), .ZN(new_n172));
  OR2_X1    g035(.A1(G183gat), .A2(G190gat), .ZN(new_n173));
  NAND3_X1  g036(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n174));
  NAND3_X1  g037(.A1(new_n172), .A2(new_n173), .A3(new_n174), .ZN(new_n175));
  AND3_X1   g038(.A1(new_n170), .A2(KEYINPUT25), .A3(new_n175), .ZN(new_n176));
  AOI21_X1  g039(.A(KEYINPUT25), .B1(new_n170), .B2(new_n175), .ZN(new_n177));
  OAI211_X1 g040(.A(new_n149), .B(new_n164), .C1(new_n176), .C2(new_n177), .ZN(new_n178));
  INV_X1    g041(.A(new_n178), .ZN(new_n179));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n180));
  NOR3_X1   g043(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n181));
  AOI21_X1  g044(.A(new_n165), .B1(G169gat), .B2(G176gat), .ZN(new_n182));
  INV_X1    g045(.A(new_n156), .ZN(new_n183));
  AOI21_X1  g046(.A(new_n181), .B1(new_n182), .B2(new_n183), .ZN(new_n184));
  AND3_X1   g047(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n185));
  AOI21_X1  g048(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n186));
  NOR2_X1   g049(.A1(G183gat), .A2(G190gat), .ZN(new_n187));
  NOR3_X1   g050(.A1(new_n185), .A2(new_n186), .A3(new_n187), .ZN(new_n188));
  OAI21_X1  g051(.A(new_n180), .B1(new_n184), .B2(new_n188), .ZN(new_n189));
  NAND3_X1  g052(.A1(new_n170), .A2(KEYINPUT25), .A3(new_n175), .ZN(new_n190));
  NAND2_X1  g053(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  AOI21_X1  g054(.A(new_n149), .B1(new_n191), .B2(new_n164), .ZN(new_n192));
  OAI21_X1  g055(.A(new_n141), .B1(new_n179), .B2(new_n192), .ZN(new_n193));
  INV_X1    g056(.A(KEYINPUT33), .ZN(new_n194));
  NAND2_X1  g057(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XOR2_X1   g058(.A(G15gat), .B(G43gat), .Z(new_n196));
  XNOR2_X1  g059(.A(G71gat), .B(G99gat), .ZN(new_n197));
  XNOR2_X1  g060(.A(new_n196), .B(new_n197), .ZN(new_n198));
  AOI21_X1  g061(.A(new_n139), .B1(new_n195), .B2(new_n198), .ZN(new_n199));
  OAI21_X1  g062(.A(new_n164), .B1(new_n176), .B2(new_n177), .ZN(new_n200));
  INV_X1    g063(.A(new_n148), .ZN(new_n201));
  NAND2_X1  g064(.A1(new_n201), .A2(new_n147), .ZN(new_n202));
  NAND4_X1  g065(.A1(new_n148), .A2(new_n145), .A3(new_n144), .A4(new_n146), .ZN(new_n203));
  NAND2_X1  g066(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g067(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g068(.A(new_n140), .B1(new_n205), .B2(new_n178), .ZN(new_n206));
  OAI211_X1 g069(.A(new_n139), .B(new_n198), .C1(new_n206), .C2(KEYINPUT33), .ZN(new_n207));
  INV_X1    g070(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g071(.A1(new_n205), .A2(new_n140), .A3(new_n178), .ZN(new_n209));
  INV_X1    g072(.A(KEYINPUT32), .ZN(new_n210));
  NAND2_X1  g073(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g074(.A1(new_n205), .A2(KEYINPUT32), .A3(new_n140), .A4(new_n178), .ZN(new_n212));
  NAND3_X1  g075(.A1(new_n211), .A2(new_n193), .A3(new_n212), .ZN(new_n213));
  NOR3_X1   g076(.A1(new_n199), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  AND3_X1   g077(.A1(new_n211), .A2(new_n193), .A3(new_n212), .ZN(new_n215));
  OAI21_X1  g078(.A(new_n198), .B1(new_n206), .B2(KEYINPUT33), .ZN(new_n216));
  NAND2_X1  g079(.A1(new_n216), .A2(KEYINPUT34), .ZN(new_n217));
  AOI21_X1  g080(.A(new_n215), .B1(new_n217), .B2(new_n207), .ZN(new_n218));
  OAI21_X1  g081(.A(new_n138), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g082(.A(new_n213), .B1(new_n199), .B2(new_n208), .ZN(new_n220));
  NAND3_X1  g083(.A1(new_n215), .A2(new_n217), .A3(new_n207), .ZN(new_n221));
  NAND3_X1  g084(.A1(new_n220), .A2(KEYINPUT36), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g085(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g086(.A(G22gat), .B(G50gat), .ZN(new_n224));
  NAND2_X1  g087(.A1(G228gat), .A2(G233gat), .ZN(new_n225));
  XNOR2_X1  g088(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g089(.A(new_n226), .ZN(new_n227));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n228));
  INV_X1    g091(.A(G211gat), .ZN(new_n229));
  INV_X1    g092(.A(G218gat), .ZN(new_n230));
  NOR2_X1   g093(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g094(.A(new_n228), .B1(KEYINPUT22), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n233));
  INV_X1    g096(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g097(.A(new_n232), .B(new_n234), .ZN(new_n235));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n236));
  NAND2_X1  g099(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g100(.A(new_n232), .B(new_n233), .ZN(new_n238));
  NAND2_X1  g101(.A1(new_n238), .A2(KEYINPUT29), .ZN(new_n239));
  AND2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n240));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n241));
  NOR2_X1   g104(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g105(.A(G141gat), .B(G148gat), .ZN(new_n243));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n244));
  AOI21_X1  g107(.A(new_n244), .B1(G155gat), .B2(G162gat), .ZN(new_n245));
  OAI21_X1  g108(.A(new_n242), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g109(.A(G148gat), .ZN(new_n247));
  NAND2_X1  g110(.A1(new_n247), .A2(G141gat), .ZN(new_n248));
  INV_X1    g111(.A(G141gat), .ZN(new_n249));
  NAND2_X1  g112(.A1(new_n249), .A2(G148gat), .ZN(new_n250));
  NAND2_X1  g113(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g114(.A(G155gat), .B(G162gat), .ZN(new_n252));
  INV_X1    g115(.A(G155gat), .ZN(new_n253));
  INV_X1    g116(.A(G162gat), .ZN(new_n254));
  OAI21_X1  g117(.A(KEYINPUT2), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g118(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g119(.A1(new_n246), .A2(new_n256), .ZN(new_n257));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g121(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g122(.A1(new_n246), .A2(new_n256), .A3(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g123(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g124(.A1(new_n237), .A2(new_n239), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g125(.A(G78gat), .B(G106gat), .ZN(new_n263));
  XNOR2_X1  g126(.A(new_n263), .B(KEYINPUT31), .ZN(new_n264));
  INV_X1    g127(.A(new_n264), .ZN(new_n265));
  INV_X1    g128(.A(new_n257), .ZN(new_n266));
  NAND2_X1  g129(.A1(new_n235), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g130(.A1(new_n262), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g131(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g132(.A(new_n265), .B1(new_n262), .B2(new_n267), .ZN(new_n270));
  OAI21_X1  g133(.A(new_n227), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g134(.A(new_n270), .ZN(new_n272));
  NAND3_X1  g135(.A1(new_n272), .A2(new_n226), .A3(new_n268), .ZN(new_n273));
  NAND2_X1  g136(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g137(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n276));
  NAND2_X1  g139(.A1(new_n204), .A2(new_n257), .ZN(new_n277));
  NAND4_X1  g140(.A1(new_n202), .A2(new_n246), .A3(new_n203), .A4(new_n256), .ZN(new_n278));
  AOI21_X1  g141(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g142(.A1(new_n246), .A2(new_n256), .A3(KEYINPUT3), .ZN(new_n280));
  AOI21_X1  g143(.A(KEYINPUT3), .B1(new_n246), .B2(new_n256), .ZN(new_n281));
  OAI21_X1  g144(.A(new_n204), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g145(.A1(new_n266), .A2(new_n149), .A3(KEYINPUT4), .ZN(new_n283));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n284));
  NAND2_X1  g147(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g148(.A1(new_n282), .A2(new_n276), .A3(new_n283), .A4(new_n285), .ZN(new_n286));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n287));
  AOI21_X1  g150(.A(new_n279), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI22_X1  g151(.A1(new_n261), .A2(new_n204), .B1(new_n284), .B2(new_n278), .ZN(new_n289));
  NAND4_X1  g152(.A1(new_n289), .A2(KEYINPUT5), .A3(new_n276), .A4(new_n283), .ZN(new_n290));
  NAND2_X1  g153(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n292));
  XNOR2_X1  g155(.A(new_n292), .B(KEYINPUT0), .ZN(new_n293));
  XNOR2_X1  g156(.A(new_n293), .B(G57gat), .ZN(new_n294));
  INV_X1    g157(.A(G85gat), .ZN(new_n295));
  XNOR2_X1  g158(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g159(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n298));
  XNOR2_X1  g161(.A(new_n294), .B(G85gat), .ZN(new_n299));
  NAND3_X1  g162(.A1(new_n288), .A2(new_n299), .A3(new_n290), .ZN(new_n300));
  NAND3_X1  g163(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g164(.A1(new_n288), .A2(new_n290), .ZN(new_n302));
  NAND3_X1  g165(.A1(new_n302), .A2(KEYINPUT6), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g166(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n305));
  INV_X1    g168(.A(G64gat), .ZN(new_n306));
  XNOR2_X1  g169(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g170(.A(G92gat), .ZN(new_n308));
  XNOR2_X1  g171(.A(new_n307), .B(new_n308), .ZN(new_n309));
  AND2_X1   g172(.A1(G226gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g173(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g174(.A1(new_n311), .A2(new_n236), .ZN(new_n312));
  NAND2_X1  g175(.A1(new_n200), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g176(.A(new_n164), .B(new_n311), .C1(new_n176), .C2(new_n177), .ZN(new_n314));
  AND3_X1   g177(.A1(new_n313), .A2(new_n235), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g178(.A(new_n235), .B1(new_n313), .B2(new_n314), .ZN(new_n316));
  OAI21_X1  g179(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g180(.A1(new_n191), .A2(new_n164), .B1(new_n236), .B2(new_n311), .ZN(new_n318));
  INV_X1    g181(.A(new_n314), .ZN(new_n319));
  OAI21_X1  g182(.A(new_n238), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g183(.A1(new_n313), .A2(new_n235), .A3(new_n314), .ZN(new_n321));
  INV_X1    g184(.A(new_n309), .ZN(new_n322));
  NAND3_X1  g185(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g186(.A1(new_n317), .A2(KEYINPUT30), .A3(new_n323), .ZN(new_n324));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n325));
  NAND4_X1  g188(.A1(new_n320), .A2(new_n321), .A3(new_n325), .A4(new_n322), .ZN(new_n326));
  NAND2_X1  g189(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g190(.A(new_n275), .B1(new_n304), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g191(.A1(new_n223), .A2(new_n328), .ZN(new_n329));
  INV_X1    g192(.A(new_n327), .ZN(new_n330));
  INV_X1    g193(.A(KEYINPUT40), .ZN(new_n331));
  NAND3_X1  g194(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n332));
  INV_X1    g195(.A(new_n276), .ZN(new_n333));
  NAND2_X1  g196(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g197(.A1(new_n277), .A2(new_n276), .A3(new_n278), .ZN(new_n335));
  NAND3_X1  g198(.A1(new_n334), .A2(KEYINPUT39), .A3(new_n335), .ZN(new_n336));
  INV_X1    g199(.A(KEYINPUT39), .ZN(new_n337));
  NAND3_X1  g200(.A1(new_n332), .A2(new_n337), .A3(new_n333), .ZN(new_n338));
  NAND3_X1  g201(.A1(new_n336), .A2(new_n296), .A3(new_n338), .ZN(new_n339));
  AOI22_X1  g202(.A1(new_n331), .A2(new_n339), .B1(new_n302), .B2(new_n299), .ZN(new_n340));
  OR2_X1    g203(.A1(new_n339), .A2(new_n331), .ZN(new_n341));
  NAND3_X1  g204(.A1(new_n330), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g205(.A(KEYINPUT37), .B1(new_n315), .B2(new_n316), .ZN(new_n343));
  INV_X1    g206(.A(KEYINPUT37), .ZN(new_n344));
  NAND3_X1  g207(.A1(new_n320), .A2(new_n321), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g208(.A1(new_n343), .A2(new_n309), .A3(new_n345), .ZN(new_n346));
  INV_X1    g209(.A(KEYINPUT38), .ZN(new_n347));
  NAND2_X1  g210(.A1(new_n323), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g211(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g212(.A1(new_n343), .A2(new_n345), .A3(new_n347), .A4(new_n309), .ZN(new_n350));
  NAND4_X1  g213(.A1(new_n301), .A2(new_n303), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g214(.A1(new_n342), .A2(new_n351), .A3(new_n275), .ZN(new_n352));
  NAND2_X1  g215(.A1(new_n220), .A2(new_n221), .ZN(new_n353));
  NAND4_X1  g216(.A1(new_n304), .A2(new_n353), .A3(new_n327), .A4(new_n275), .ZN(new_n354));
  NAND2_X1  g217(.A1(new_n354), .A2(KEYINPUT35), .ZN(new_n355));
  AOI21_X1  g218(.A(new_n274), .B1(new_n301), .B2(new_n303), .ZN(new_n356));
  INV_X1    g219(.A(KEYINPUT35), .ZN(new_n357));
  NAND4_X1  g220(.A1(new_n356), .A2(new_n357), .A3(new_n353), .A4(new_n327), .ZN(new_n358));
  AOI22_X1  g221(.A1(new_n329), .A2(new_n352), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g222(.A(G15gat), .B(G22gat), .ZN(new_n360));
  INV_X1    g223(.A(G1gat), .ZN(new_n361));
  NAND2_X1  g224(.A1(new_n361), .A2(KEYINPUT16), .ZN(new_n362));
  AND2_X1   g225(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g226(.A1(new_n360), .A2(G1gat), .ZN(new_n364));
  OAI21_X1  g227(.A(G8gat), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g228(.A1(new_n360), .A2(new_n362), .ZN(new_n366));
  INV_X1    g229(.A(G8gat), .ZN(new_n367));
  OAI211_X1 g230(.A(new_n366), .B(new_n367), .C1(G1gat), .C2(new_n360), .ZN(new_n368));
  AND2_X1   g231(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g232(.A(G43gat), .B(G50gat), .ZN(new_n370));
  NAND2_X1  g233(.A1(new_n370), .A2(KEYINPUT15), .ZN(new_n371));
  NAND2_X1  g234(.A1(G29gat), .A2(G36gat), .ZN(new_n372));
  NOR2_X1   g235(.A1(G29gat), .A2(G36gat), .ZN(new_n373));
  OAI21_X1  g236(.A(new_n372), .B1(new_n373), .B2(KEYINPUT14), .ZN(new_n374));
  INV_X1    g237(.A(new_n374), .ZN(new_n375));
  INV_X1    g238(.A(G43gat), .ZN(new_n376));
  INV_X1    g239(.A(G50gat), .ZN(new_n377));
  NAND2_X1  g240(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g241(.A(KEYINPUT15), .ZN(new_n379));
  NAND2_X1  g242(.A1(G43gat), .A2(G50gat), .ZN(new_n380));
  NAND3_X1  g243(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g244(.A1(new_n373), .A2(KEYINPUT14), .ZN(new_n382));
  NAND4_X1  g245(.A1(new_n371), .A2(new_n375), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  INV_X1    g246(.A(new_n382), .ZN(new_n384));
  OAI211_X1 g247(.A(KEYINPUT15), .B(new_n370), .C1(new_n384), .C2(new_n374), .ZN(new_n385));
  NAND2_X1  g248(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g250(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g251(.A1(new_n383), .A2(KEYINPUT17), .A3(new_n385), .ZN(new_n389));
  NAND3_X1  g252(.A1(new_n369), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g253(.A1(G229gat), .A2(G233gat), .ZN(new_n391));
  NAND2_X1  g254(.A1(new_n365), .A2(new_n368), .ZN(new_n392));
  NAND2_X1  g255(.A1(new_n392), .A2(new_n386), .ZN(new_n393));
  NAND3_X1  g256(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g257(.A(KEYINPUT18), .ZN(new_n395));
  NAND2_X1  g258(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g259(.A1(new_n390), .A2(KEYINPUT18), .A3(new_n391), .A4(new_n393), .ZN(new_n397));
  XNOR2_X1  g260(.A(new_n391), .B(KEYINPUT13), .ZN(new_n398));
  INV_X1    g261(.A(new_n398), .ZN(new_n399));
  INV_X1    g262(.A(new_n393), .ZN(new_n400));
  NOR2_X1   g263(.A1(new_n392), .A2(new_n386), .ZN(new_n401));
  OAI21_X1  g264(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g265(.A1(new_n396), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g266(.A(G113gat), .B(G141gat), .ZN(new_n404));
  INV_X1    g267(.A(KEYINPUT11), .ZN(new_n405));
  XNOR2_X1  g268(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g269(.A1(new_n406), .A2(G169gat), .ZN(new_n407));
  XNOR2_X1  g270(.A(new_n404), .B(KEYINPUT11), .ZN(new_n408));
  NAND2_X1  g271(.A1(new_n408), .A2(new_n166), .ZN(new_n409));
  NAND2_X1  g272(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g273(.A(G197gat), .ZN(new_n411));
  NAND2_X1  g274(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g275(.A1(new_n407), .A2(new_n409), .A3(G197gat), .ZN(new_n413));
  NAND3_X1  g276(.A1(new_n412), .A2(KEYINPUT12), .A3(new_n413), .ZN(new_n414));
  INV_X1    g277(.A(KEYINPUT12), .ZN(new_n415));
  AND3_X1   g278(.A1(new_n407), .A2(new_n409), .A3(G197gat), .ZN(new_n416));
  AOI21_X1  g279(.A(G197gat), .B1(new_n407), .B2(new_n409), .ZN(new_n417));
  OAI21_X1  g280(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g281(.A1(new_n403), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g282(.A1(new_n418), .A2(new_n414), .ZN(new_n420));
  NAND4_X1  g283(.A1(new_n396), .A2(new_n420), .A3(new_n397), .A4(new_n402), .ZN(new_n421));
  NAND2_X1  g284(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g285(.A(new_n422), .ZN(new_n423));
  INV_X1    g286(.A(KEYINPUT21), .ZN(new_n424));
  XOR2_X1   g287(.A(G71gat), .B(G78gat), .Z(new_n425));
  INV_X1    g288(.A(new_n425), .ZN(new_n426));
  XOR2_X1   g289(.A(G57gat), .B(G64gat), .Z(new_n427));
  NAND2_X1  g290(.A1(G71gat), .A2(G78gat), .ZN(new_n428));
  INV_X1    g291(.A(KEYINPUT9), .ZN(new_n429));
  NAND2_X1  g292(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g293(.A1(new_n426), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g294(.A1(new_n427), .A2(new_n430), .ZN(new_n432));
  NAND2_X1  g295(.A1(new_n432), .A2(new_n425), .ZN(new_n433));
  NAND2_X1  g296(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g297(.A(new_n369), .B1(new_n424), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n436));
  INV_X1    g299(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g300(.A(new_n435), .B(new_n437), .ZN(new_n438));
  XNOR2_X1  g301(.A(G127gat), .B(G155gat), .ZN(new_n439));
  XNOR2_X1  g302(.A(new_n439), .B(KEYINPUT19), .ZN(new_n440));
  XOR2_X1   g303(.A(new_n440), .B(KEYINPUT20), .Z(new_n441));
  INV_X1    g304(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g305(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g306(.A(new_n435), .B(new_n436), .ZN(new_n444));
  NAND2_X1  g307(.A1(new_n444), .A2(new_n441), .ZN(new_n445));
  NAND2_X1  g308(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g309(.A1(new_n434), .A2(new_n424), .ZN(new_n447));
  XNOR2_X1  g310(.A(G183gat), .B(G211gat), .ZN(new_n448));
  XOR2_X1   g311(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g312(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g313(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g314(.A1(new_n443), .A2(new_n445), .A3(new_n449), .ZN(new_n452));
  NAND2_X1  g315(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n454));
  XNOR2_X1  g317(.A(new_n454), .B(KEYINPUT7), .ZN(new_n455));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n456));
  AOI22_X1  g319(.A1(KEYINPUT8), .A2(new_n456), .B1(new_n295), .B2(new_n308), .ZN(new_n457));
  NAND2_X1  g320(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g321(.A(G99gat), .B(G106gat), .Z(new_n459));
  NAND2_X1  g322(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g323(.A(new_n459), .ZN(new_n461));
  NAND3_X1  g324(.A1(new_n461), .A2(new_n455), .A3(new_n457), .ZN(new_n462));
  AOI22_X1  g325(.A1(new_n460), .A2(new_n462), .B1(new_n431), .B2(new_n433), .ZN(new_n463));
  NAND2_X1  g326(.A1(new_n460), .A2(new_n462), .ZN(new_n464));
  NOR2_X1   g327(.A1(new_n464), .A2(new_n434), .ZN(new_n465));
  INV_X1    g328(.A(KEYINPUT10), .ZN(new_n466));
  AOI21_X1  g329(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g330(.A1(G230gat), .A2(G233gat), .ZN(new_n468));
  OAI21_X1  g331(.A(KEYINPUT10), .B1(new_n464), .B2(new_n434), .ZN(new_n469));
  NAND3_X1  g332(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g333(.A1(new_n465), .A2(new_n463), .ZN(new_n471));
  OAI21_X1  g334(.A(new_n470), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g335(.A(G120gat), .B(G148gat), .ZN(new_n473));
  XNOR2_X1  g336(.A(new_n473), .B(new_n167), .ZN(new_n474));
  INV_X1    g337(.A(G204gat), .ZN(new_n475));
  XNOR2_X1  g338(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XNOR2_X1  g339(.A(new_n472), .B(new_n476), .ZN(new_n477));
  INV_X1    g340(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n479));
  INV_X1    g342(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g343(.A1(new_n480), .A2(KEYINPUT41), .ZN(new_n481));
  XNOR2_X1  g344(.A(new_n481), .B(G218gat), .ZN(new_n482));
  INV_X1    g345(.A(new_n482), .ZN(new_n483));
  AND2_X1   g346(.A1(new_n460), .A2(new_n462), .ZN(new_n484));
  AOI22_X1  g347(.A1(new_n484), .A2(new_n386), .B1(KEYINPUT41), .B2(new_n480), .ZN(new_n485));
  NAND3_X1  g348(.A1(new_n388), .A2(new_n464), .A3(new_n389), .ZN(new_n486));
  XNOR2_X1  g349(.A(G134gat), .B(G162gat), .ZN(new_n487));
  XNOR2_X1  g350(.A(new_n487), .B(new_n150), .ZN(new_n488));
  INV_X1    g351(.A(new_n488), .ZN(new_n489));
  AND3_X1   g352(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g353(.A(new_n489), .B1(new_n485), .B2(new_n486), .ZN(new_n491));
  OAI21_X1  g354(.A(new_n483), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g355(.A1(new_n485), .A2(new_n486), .ZN(new_n493));
  NAND2_X1  g356(.A1(new_n493), .A2(new_n488), .ZN(new_n494));
  NAND3_X1  g357(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n495));
  NAND3_X1  g358(.A1(new_n494), .A2(new_n482), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g359(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g360(.A1(new_n453), .A2(new_n478), .A3(new_n497), .ZN(new_n498));
  NOR3_X1   g361(.A1(new_n359), .A2(new_n423), .A3(new_n498), .ZN(new_n499));
  INV_X1    g362(.A(new_n304), .ZN(new_n500));
  NAND2_X1  g363(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g364(.A(new_n501), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g365(.A1(new_n499), .A2(new_n330), .ZN(new_n503));
  XOR2_X1   g366(.A(KEYINPUT16), .B(G8gat), .Z(new_n504));
  NAND3_X1  g367(.A1(new_n503), .A2(KEYINPUT42), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g368(.A1(new_n499), .A2(new_n330), .A3(new_n504), .ZN(new_n506));
  INV_X1    g369(.A(KEYINPUT42), .ZN(new_n507));
  NAND2_X1  g370(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g371(.A(new_n505), .B(new_n508), .C1(new_n367), .C2(new_n503), .ZN(G1325gat));
  INV_X1    g372(.A(G15gat), .ZN(new_n510));
  NAND3_X1  g373(.A1(new_n499), .A2(new_n510), .A3(new_n353), .ZN(new_n511));
  AND2_X1   g374(.A1(new_n499), .A2(new_n223), .ZN(new_n512));
  OAI21_X1  g375(.A(new_n511), .B1(new_n512), .B2(new_n510), .ZN(G1326gat));
  NAND2_X1  g376(.A1(new_n499), .A2(new_n274), .ZN(new_n514));
  XNOR2_X1  g377(.A(KEYINPUT43), .B(G22gat), .ZN(new_n515));
  XNOR2_X1  g378(.A(new_n514), .B(new_n515), .ZN(G1327gat));
  NAND2_X1  g379(.A1(new_n355), .A2(new_n358), .ZN(new_n517));
  AND2_X1   g380(.A1(new_n219), .A2(new_n222), .ZN(new_n518));
  NAND2_X1  g381(.A1(new_n304), .A2(new_n327), .ZN(new_n519));
  NAND2_X1  g382(.A1(new_n519), .A2(new_n274), .ZN(new_n520));
  NAND3_X1  g383(.A1(new_n518), .A2(new_n520), .A3(new_n352), .ZN(new_n521));
  AOI21_X1  g384(.A(new_n497), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  INV_X1    g385(.A(G29gat), .ZN(new_n523));
  NOR3_X1   g386(.A1(new_n453), .A2(new_n423), .A3(new_n477), .ZN(new_n524));
  NAND4_X1  g387(.A1(new_n522), .A2(new_n523), .A3(new_n500), .A4(new_n524), .ZN(new_n525));
  XNOR2_X1  g388(.A(new_n525), .B(KEYINPUT45), .ZN(new_n526));
  INV_X1    g389(.A(new_n524), .ZN(new_n527));
  OAI21_X1  g390(.A(KEYINPUT44), .B1(new_n359), .B2(new_n497), .ZN(new_n528));
  NAND2_X1  g391(.A1(new_n517), .A2(new_n521), .ZN(new_n529));
  INV_X1    g392(.A(KEYINPUT44), .ZN(new_n530));
  AND2_X1   g393(.A1(new_n492), .A2(new_n496), .ZN(new_n531));
  NAND3_X1  g394(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g395(.A(new_n527), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g396(.A1(new_n533), .A2(new_n500), .ZN(new_n534));
  OAI21_X1  g397(.A(new_n526), .B1(new_n534), .B2(new_n523), .ZN(G1328gat));
  NAND2_X1  g398(.A1(new_n529), .A2(new_n531), .ZN(new_n536));
  NOR4_X1   g399(.A1(new_n536), .A2(G36gat), .A3(new_n327), .A4(new_n527), .ZN(new_n537));
  XNOR2_X1  g400(.A(new_n537), .B(KEYINPUT46), .ZN(new_n538));
  NAND2_X1  g401(.A1(new_n533), .A2(new_n330), .ZN(new_n539));
  NAND2_X1  g402(.A1(new_n539), .A2(G36gat), .ZN(new_n540));
  NAND2_X1  g403(.A1(new_n538), .A2(new_n540), .ZN(G1329gat));
  INV_X1    g404(.A(KEYINPUT47), .ZN(new_n542));
  AOI21_X1  g405(.A(new_n376), .B1(new_n533), .B2(new_n223), .ZN(new_n543));
  NOR2_X1   g406(.A1(new_n536), .A2(new_n527), .ZN(new_n544));
  INV_X1    g407(.A(new_n353), .ZN(new_n545));
  NOR2_X1   g408(.A1(new_n545), .A2(G43gat), .ZN(new_n546));
  NAND2_X1  g409(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g410(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g411(.A(new_n542), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g412(.A1(new_n522), .A2(new_n530), .ZN(new_n550));
  AOI211_X1 g413(.A(KEYINPUT44), .B(new_n497), .C1(new_n517), .C2(new_n521), .ZN(new_n551));
  OAI211_X1 g414(.A(new_n223), .B(new_n524), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g415(.A1(new_n552), .A2(G43gat), .ZN(new_n553));
  NAND3_X1  g416(.A1(new_n553), .A2(KEYINPUT47), .A3(new_n547), .ZN(new_n554));
  NAND2_X1  g417(.A1(new_n549), .A2(new_n554), .ZN(G1330gat));
  INV_X1    g418(.A(KEYINPUT48), .ZN(new_n556));
  AOI21_X1  g419(.A(new_n377), .B1(new_n533), .B2(new_n274), .ZN(new_n557));
  NOR4_X1   g420(.A1(new_n536), .A2(G50gat), .A3(new_n275), .A4(new_n527), .ZN(new_n558));
  OAI21_X1  g421(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g422(.A(new_n274), .B(new_n524), .C1(new_n550), .C2(new_n551), .ZN(new_n560));
  NAND2_X1  g423(.A1(new_n560), .A2(G50gat), .ZN(new_n561));
  INV_X1    g424(.A(new_n558), .ZN(new_n562));
  NAND3_X1  g425(.A1(new_n561), .A2(KEYINPUT48), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g426(.A1(new_n559), .A2(new_n563), .ZN(G1331gat));
  NAND3_X1  g427(.A1(new_n453), .A2(new_n423), .A3(new_n497), .ZN(new_n565));
  NOR3_X1   g428(.A1(new_n359), .A2(new_n478), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g429(.A1(new_n566), .A2(new_n500), .ZN(new_n567));
  XNOR2_X1  g430(.A(new_n567), .B(G57gat), .ZN(G1332gat));
  INV_X1    g431(.A(KEYINPUT49), .ZN(new_n569));
  OAI211_X1 g432(.A(new_n566), .B(new_n330), .C1(new_n569), .C2(new_n306), .ZN(new_n570));
  NAND2_X1  g433(.A1(new_n569), .A2(new_n306), .ZN(new_n571));
  XNOR2_X1  g434(.A(new_n570), .B(new_n571), .ZN(G1333gat));
  NAND2_X1  g435(.A1(new_n566), .A2(new_n223), .ZN(new_n573));
  NAND2_X1  g436(.A1(new_n573), .A2(G71gat), .ZN(new_n574));
  INV_X1    g437(.A(G71gat), .ZN(new_n575));
  NAND3_X1  g438(.A1(new_n566), .A2(new_n575), .A3(new_n353), .ZN(new_n576));
  NAND2_X1  g439(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g440(.A(KEYINPUT50), .ZN(new_n578));
  NAND2_X1  g441(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g442(.A1(new_n574), .A2(KEYINPUT50), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g443(.A1(new_n579), .A2(new_n580), .ZN(G1334gat));
  NAND2_X1  g444(.A1(new_n566), .A2(new_n274), .ZN(new_n582));
  XNOR2_X1  g445(.A(new_n582), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g446(.A1(new_n453), .A2(new_n422), .ZN(new_n584));
  NAND2_X1  g447(.A1(new_n584), .A2(new_n477), .ZN(new_n585));
  AOI21_X1  g448(.A(new_n585), .B1(new_n528), .B2(new_n532), .ZN(new_n586));
  AND2_X1   g449(.A1(new_n586), .A2(new_n500), .ZN(new_n587));
  NAND3_X1  g450(.A1(new_n522), .A2(KEYINPUT51), .A3(new_n584), .ZN(new_n588));
  INV_X1    g451(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g452(.A(KEYINPUT51), .B1(new_n522), .B2(new_n584), .ZN(new_n590));
  OAI211_X1 g453(.A(new_n295), .B(new_n500), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  OAI22_X1  g454(.A1(new_n587), .A2(new_n295), .B1(new_n591), .B2(new_n478), .ZN(G1336gat));
  AOI21_X1  g455(.A(new_n308), .B1(new_n586), .B2(new_n330), .ZN(new_n593));
  NOR3_X1   g456(.A1(new_n478), .A2(G92gat), .A3(new_n327), .ZN(new_n594));
  INV_X1    g457(.A(new_n594), .ZN(new_n595));
  INV_X1    g458(.A(KEYINPUT51), .ZN(new_n596));
  INV_X1    g459(.A(new_n584), .ZN(new_n597));
  OAI21_X1  g460(.A(new_n596), .B1(new_n536), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g461(.A(new_n595), .B1(new_n598), .B2(new_n588), .ZN(new_n599));
  OAI21_X1  g462(.A(KEYINPUT52), .B1(new_n593), .B2(new_n599), .ZN(new_n600));
  INV_X1    g463(.A(new_n585), .ZN(new_n601));
  OAI211_X1 g464(.A(new_n330), .B(new_n601), .C1(new_n550), .C2(new_n551), .ZN(new_n602));
  NAND2_X1  g465(.A1(new_n602), .A2(G92gat), .ZN(new_n603));
  INV_X1    g466(.A(KEYINPUT52), .ZN(new_n604));
  OAI21_X1  g467(.A(new_n594), .B1(new_n589), .B2(new_n590), .ZN(new_n605));
  NAND3_X1  g468(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g469(.A1(new_n600), .A2(new_n606), .ZN(G1337gat));
  NAND2_X1  g470(.A1(new_n586), .A2(new_n223), .ZN(new_n608));
  NAND2_X1  g471(.A1(new_n608), .A2(G99gat), .ZN(new_n609));
  NOR3_X1   g472(.A1(new_n545), .A2(new_n478), .A3(G99gat), .ZN(new_n610));
  OAI21_X1  g473(.A(new_n610), .B1(new_n589), .B2(new_n590), .ZN(new_n611));
  NAND2_X1  g474(.A1(new_n609), .A2(new_n611), .ZN(G1338gat));
  INV_X1    g475(.A(G106gat), .ZN(new_n613));
  AOI21_X1  g476(.A(new_n613), .B1(new_n586), .B2(new_n274), .ZN(new_n614));
  NOR3_X1   g477(.A1(new_n478), .A2(new_n275), .A3(G106gat), .ZN(new_n615));
  INV_X1    g478(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g479(.A(new_n616), .B1(new_n598), .B2(new_n588), .ZN(new_n617));
  OAI21_X1  g480(.A(KEYINPUT53), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  OAI211_X1 g481(.A(new_n274), .B(new_n601), .C1(new_n550), .C2(new_n551), .ZN(new_n619));
  NAND2_X1  g482(.A1(new_n619), .A2(G106gat), .ZN(new_n620));
  INV_X1    g483(.A(KEYINPUT53), .ZN(new_n621));
  OAI21_X1  g484(.A(new_n615), .B1(new_n589), .B2(new_n590), .ZN(new_n622));
  NAND3_X1  g485(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g486(.A1(new_n618), .A2(new_n623), .ZN(G1339gat));
  NOR2_X1   g487(.A1(new_n472), .A2(new_n476), .ZN(new_n625));
  NOR3_X1   g488(.A1(new_n400), .A2(new_n401), .A3(new_n399), .ZN(new_n626));
  AOI21_X1  g489(.A(new_n391), .B1(new_n390), .B2(new_n393), .ZN(new_n627));
  OAI211_X1 g490(.A(new_n413), .B(new_n412), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g491(.A1(new_n421), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g492(.A(new_n625), .B1(new_n531), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g493(.A1(new_n419), .A2(new_n421), .A3(new_n497), .ZN(new_n631));
  INV_X1    g494(.A(KEYINPUT55), .ZN(new_n632));
  AOI21_X1  g495(.A(new_n468), .B1(new_n467), .B2(new_n469), .ZN(new_n633));
  INV_X1    g496(.A(KEYINPUT54), .ZN(new_n634));
  OAI21_X1  g497(.A(new_n470), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND4_X1  g498(.A1(new_n467), .A2(KEYINPUT54), .A3(new_n468), .A4(new_n469), .ZN(new_n636));
  NAND2_X1  g499(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g500(.A(new_n632), .B1(new_n637), .B2(new_n476), .ZN(new_n638));
  INV_X1    g501(.A(new_n476), .ZN(new_n639));
  AOI211_X1 g502(.A(KEYINPUT55), .B(new_n639), .C1(new_n635), .C2(new_n636), .ZN(new_n640));
  OAI211_X1 g503(.A(new_n630), .B(new_n631), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  NAND4_X1  g504(.A1(new_n477), .A2(new_n421), .A3(new_n497), .A4(new_n628), .ZN(new_n642));
  AOI21_X1  g505(.A(new_n453), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g506(.A1(new_n498), .A2(new_n422), .ZN(new_n644));
  NOR2_X1   g507(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g508(.A1(new_n645), .A2(new_n304), .ZN(new_n646));
  NOR2_X1   g509(.A1(new_n545), .A2(new_n274), .ZN(new_n647));
  NAND3_X1  g510(.A1(new_n646), .A2(new_n327), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g511(.A1(new_n648), .A2(new_n423), .ZN(new_n649));
  XNOR2_X1  g512(.A(new_n649), .B(new_n142), .ZN(G1340gat));
  NOR2_X1   g513(.A1(new_n648), .A2(new_n478), .ZN(new_n651));
  XNOR2_X1  g514(.A(new_n651), .B(new_n143), .ZN(G1341gat));
  NAND4_X1  g515(.A1(new_n646), .A2(new_n327), .A3(new_n453), .A4(new_n647), .ZN(new_n653));
  XNOR2_X1  g516(.A(new_n653), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g517(.A1(new_n648), .A2(new_n497), .ZN(new_n655));
  NAND2_X1  g518(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n656));
  INV_X1    g519(.A(KEYINPUT56), .ZN(new_n657));
  INV_X1    g520(.A(G134gat), .ZN(new_n658));
  NAND2_X1  g521(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g522(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  OAI211_X1 g523(.A(new_n657), .B(new_n658), .C1(new_n648), .C2(new_n497), .ZN(new_n661));
  AND2_X1   g524(.A1(new_n660), .A2(new_n661), .ZN(G1343gat));
  NOR2_X1   g525(.A1(new_n223), .A2(new_n304), .ZN(new_n663));
  NAND2_X1  g526(.A1(new_n663), .A2(new_n327), .ZN(new_n664));
  OAI21_X1  g527(.A(new_n274), .B1(new_n643), .B2(new_n644), .ZN(new_n665));
  INV_X1    g528(.A(KEYINPUT57), .ZN(new_n666));
  NAND2_X1  g529(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI211_X1 g530(.A(KEYINPUT57), .B(new_n274), .C1(new_n643), .C2(new_n644), .ZN(new_n668));
  AOI21_X1  g531(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g532(.A(new_n249), .B1(new_n669), .B2(new_n422), .ZN(new_n670));
  NAND2_X1  g533(.A1(new_n641), .A2(new_n642), .ZN(new_n671));
  INV_X1    g534(.A(new_n453), .ZN(new_n672));
  NAND2_X1  g535(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g536(.A(new_n644), .ZN(new_n674));
  NAND2_X1  g537(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g538(.A1(new_n675), .A2(new_n274), .A3(new_n663), .ZN(new_n676));
  NOR4_X1   g539(.A1(new_n676), .A2(G141gat), .A3(new_n423), .A4(new_n330), .ZN(new_n677));
  OAI21_X1  g540(.A(KEYINPUT58), .B1(new_n670), .B2(new_n677), .ZN(new_n678));
  INV_X1    g541(.A(new_n676), .ZN(new_n679));
  NAND4_X1  g542(.A1(new_n679), .A2(new_n249), .A3(new_n422), .A4(new_n327), .ZN(new_n680));
  INV_X1    g543(.A(KEYINPUT58), .ZN(new_n681));
  AOI211_X1 g544(.A(new_n423), .B(new_n664), .C1(new_n667), .C2(new_n668), .ZN(new_n682));
  OAI211_X1 g545(.A(new_n680), .B(new_n681), .C1(new_n682), .C2(new_n249), .ZN(new_n683));
  NAND2_X1  g546(.A1(new_n678), .A2(new_n683), .ZN(G1344gat));
  NOR2_X1   g547(.A1(new_n676), .A2(new_n330), .ZN(new_n685));
  NAND3_X1  g548(.A1(new_n685), .A2(new_n247), .A3(new_n477), .ZN(new_n686));
  AOI211_X1 g549(.A(KEYINPUT59), .B(new_n247), .C1(new_n669), .C2(new_n477), .ZN(new_n687));
  INV_X1    g550(.A(KEYINPUT59), .ZN(new_n688));
  INV_X1    g551(.A(new_n664), .ZN(new_n689));
  AOI21_X1  g552(.A(KEYINPUT57), .B1(new_n675), .B2(new_n274), .ZN(new_n690));
  INV_X1    g553(.A(new_n668), .ZN(new_n691));
  OAI211_X1 g554(.A(new_n477), .B(new_n689), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  AOI21_X1  g555(.A(new_n688), .B1(new_n692), .B2(G148gat), .ZN(new_n693));
  OAI21_X1  g556(.A(new_n686), .B1(new_n687), .B2(new_n693), .ZN(G1345gat));
  NAND3_X1  g557(.A1(new_n685), .A2(new_n253), .A3(new_n453), .ZN(new_n695));
  AND2_X1   g558(.A1(new_n669), .A2(new_n453), .ZN(new_n696));
  OAI21_X1  g559(.A(new_n695), .B1(new_n696), .B2(new_n253), .ZN(G1346gat));
  NAND3_X1  g560(.A1(new_n685), .A2(new_n254), .A3(new_n531), .ZN(new_n698));
  AND2_X1   g561(.A1(new_n669), .A2(new_n531), .ZN(new_n699));
  OAI21_X1  g562(.A(new_n698), .B1(new_n699), .B2(new_n254), .ZN(G1347gat));
  NAND2_X1  g563(.A1(new_n356), .A2(new_n353), .ZN(new_n701));
  NOR2_X1   g564(.A1(new_n645), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g565(.A1(new_n702), .A2(new_n519), .ZN(new_n703));
  OAI21_X1  g566(.A(G169gat), .B1(new_n703), .B2(new_n423), .ZN(new_n704));
  NOR2_X1   g567(.A1(new_n423), .A2(new_n327), .ZN(new_n705));
  NAND3_X1  g568(.A1(new_n702), .A2(new_n166), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g569(.A1(new_n704), .A2(new_n706), .ZN(G1348gat));
  OAI21_X1  g570(.A(G176gat), .B1(new_n703), .B2(new_n478), .ZN(new_n708));
  NAND4_X1  g571(.A1(new_n702), .A2(new_n167), .A3(new_n330), .A4(new_n477), .ZN(new_n709));
  NAND2_X1  g572(.A1(new_n708), .A2(new_n709), .ZN(G1349gat));
  OAI21_X1  g573(.A(G183gat), .B1(new_n703), .B2(new_n672), .ZN(new_n711));
  NOR2_X1   g574(.A1(new_n672), .A2(new_n327), .ZN(new_n712));
  OAI211_X1 g575(.A(new_n702), .B(new_n712), .C1(new_n152), .C2(new_n151), .ZN(new_n713));
  NAND2_X1  g576(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g577(.A1(new_n714), .A2(KEYINPUT60), .ZN(new_n715));
  INV_X1    g578(.A(KEYINPUT60), .ZN(new_n716));
  NAND3_X1  g579(.A1(new_n711), .A2(new_n716), .A3(new_n713), .ZN(new_n717));
  NAND2_X1  g580(.A1(new_n715), .A2(new_n717), .ZN(G1350gat));
  NAND4_X1  g581(.A1(new_n702), .A2(new_n150), .A3(new_n330), .A4(new_n531), .ZN(new_n719));
  NAND3_X1  g582(.A1(new_n702), .A2(new_n519), .A3(new_n531), .ZN(new_n720));
  INV_X1    g583(.A(KEYINPUT61), .ZN(new_n721));
  NAND3_X1  g584(.A1(new_n720), .A2(new_n721), .A3(G190gat), .ZN(new_n722));
  INV_X1    g585(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g586(.A(new_n721), .B1(new_n720), .B2(G190gat), .ZN(new_n724));
  OAI21_X1  g587(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(G1351gat));
  NOR2_X1   g588(.A1(new_n223), .A2(new_n500), .ZN(new_n726));
  NAND2_X1  g589(.A1(new_n726), .A2(new_n330), .ZN(new_n727));
  AOI21_X1  g590(.A(new_n727), .B1(new_n667), .B2(new_n668), .ZN(new_n728));
  AND2_X1   g591(.A1(new_n728), .A2(new_n422), .ZN(new_n729));
  NAND3_X1  g592(.A1(new_n675), .A2(new_n274), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g593(.A1(new_n705), .A2(new_n411), .ZN(new_n731));
  OAI22_X1  g594(.A1(new_n729), .A2(new_n411), .B1(new_n730), .B2(new_n731), .ZN(G1352gat));
  NOR2_X1   g595(.A1(new_n730), .A2(new_n327), .ZN(new_n733));
  NOR2_X1   g596(.A1(new_n478), .A2(G204gat), .ZN(new_n734));
  AND3_X1   g597(.A1(new_n733), .A2(KEYINPUT62), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g598(.A(KEYINPUT62), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  AND2_X1   g599(.A1(new_n728), .A2(new_n477), .ZN(new_n737));
  OAI22_X1  g600(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n475), .ZN(G1353gat));
  NAND3_X1  g601(.A1(new_n733), .A2(new_n229), .A3(new_n453), .ZN(new_n739));
  INV_X1    g602(.A(KEYINPUT63), .ZN(new_n740));
  AOI211_X1 g603(.A(new_n740), .B(new_n229), .C1(new_n728), .C2(new_n453), .ZN(new_n741));
  INV_X1    g604(.A(new_n727), .ZN(new_n742));
  OAI211_X1 g605(.A(new_n453), .B(new_n742), .C1(new_n690), .C2(new_n691), .ZN(new_n743));
  AOI21_X1  g606(.A(KEYINPUT63), .B1(new_n743), .B2(G211gat), .ZN(new_n744));
  OAI21_X1  g607(.A(new_n739), .B1(new_n741), .B2(new_n744), .ZN(G1354gat));
  NAND3_X1  g608(.A1(new_n733), .A2(new_n230), .A3(new_n531), .ZN(new_n746));
  AND2_X1   g609(.A1(new_n728), .A2(new_n531), .ZN(new_n747));
  OAI21_X1  g610(.A(new_n746), .B1(new_n747), .B2(new_n230), .ZN(G1355gat));
endmodule


