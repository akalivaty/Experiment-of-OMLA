//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT65), .B(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  OR3_X1    g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G68), .Z(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NOR2_X1   g0044(.A1(G20), .A2(G33), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G150), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n213), .A2(G33), .ZN(new_n249));
  OAI221_X1 g0049(.A(new_n247), .B1(new_n207), .B2(new_n201), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n214), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n254), .A2(new_n207), .A3(G1), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n252), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n207), .A2(G1), .ZN(new_n257));
  INV_X1    g0057(.A(G50), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n256), .A2(new_n259), .B1(new_n258), .B2(new_n255), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G222), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(G1698), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n267), .B1(new_n202), .B2(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n274), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n276), .B1(new_n281), .B2(G226), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n273), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G179), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  AOI211_X1 g0085(.A(new_n262), .B(new_n284), .C1(new_n285), .C2(new_n283), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(G200), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT9), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n261), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n262), .A2(KEYINPUT9), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  OR3_X1    g0091(.A1(new_n289), .A2(new_n291), .A3(KEYINPUT10), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT10), .B1(new_n289), .B2(new_n291), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n286), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT71), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n268), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(new_n297), .B2(new_n269), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n268), .A2(KEYINPUT71), .A3(G223), .A4(new_n296), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n265), .A2(new_n296), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n301), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n279), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n276), .B1(new_n281), .B2(G232), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(G200), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G226), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n270), .A2(new_n307), .B1(new_n277), .B2(new_n220), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n298), .B2(new_n299), .ZN(new_n309));
  OAI211_X1 g0109(.A(G190), .B(new_n304), .C1(new_n309), .C2(new_n279), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n256), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n248), .A2(new_n257), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(KEYINPUT70), .B2(new_n313), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n314), .A2(new_n315), .B1(new_n255), .B2(new_n248), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT7), .B1(new_n268), .B2(G20), .ZN(new_n317));
  OR2_X1    g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT65), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n318), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n317), .B(G68), .C1(KEYINPUT7), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G58), .A2(G68), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT69), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT69), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G58), .A3(G68), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n328), .C1(G58), .C2(G68), .ZN(new_n329));
  AOI22_X1  g0129(.A1(G159), .A2(new_n246), .B1(new_n329), .B2(G20), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(new_n330), .A3(KEYINPUT16), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n252), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(KEYINPUT7), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n265), .A2(new_n334), .A3(new_n207), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(G68), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT16), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n316), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n311), .A2(new_n339), .A3(KEYINPUT17), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n330), .A2(new_n336), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n252), .B(new_n331), .C1(new_n341), .C2(KEYINPUT16), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n306), .A2(new_n342), .A3(new_n316), .A4(new_n310), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(G179), .B(new_n304), .C1(new_n309), .C2(new_n279), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT71), .B1(new_n266), .B2(G223), .ZN(new_n347));
  INV_X1    g0147(.A(new_n299), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n302), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n305), .B1(new_n349), .B2(new_n272), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n346), .B1(new_n350), .B2(new_n285), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n351), .A2(KEYINPUT18), .A3(new_n338), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT18), .B1(new_n351), .B2(new_n338), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n340), .B(new_n345), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n218), .A2(G20), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n249), .B2(new_n202), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT66), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n245), .B(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n258), .ZN(new_n360));
  OAI211_X1 g0160(.A(KEYINPUT11), .B(new_n252), .C1(new_n357), .C2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n254), .A2(G1), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G20), .ZN(new_n363));
  OR3_X1    g0163(.A1(new_n363), .A2(KEYINPUT12), .A3(G68), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT12), .B1(new_n363), .B2(G68), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n257), .A2(new_n218), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n364), .A2(new_n365), .B1(new_n256), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n356), .B1(new_n249), .B2(new_n202), .C1(new_n258), .C2(new_n359), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT11), .B1(new_n369), .B2(new_n252), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n230), .A2(G1698), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n268), .B(new_n373), .C1(G226), .C2(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G97), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n272), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT13), .ZN(new_n378));
  INV_X1    g0178(.A(new_n276), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n280), .B2(new_n219), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n279), .B1(new_n374), .B2(new_n375), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT13), .B1(new_n383), .B2(new_n380), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(G169), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n382), .A2(G179), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n386), .B1(new_n385), .B2(G169), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n372), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n385), .A2(G200), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n382), .A2(G190), .A3(new_n384), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n392), .A2(new_n371), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n257), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G77), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n312), .A2(new_n399), .B1(G77), .B2(new_n363), .ZN(new_n400));
  INV_X1    g0200(.A(new_n248), .ZN(new_n401));
  INV_X1    g0201(.A(new_n213), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n246), .A2(new_n401), .B1(new_n402), .B2(G77), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT15), .B(G87), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n249), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n405), .B2(new_n252), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n407));
  OR2_X1    g0207(.A1(KEYINPUT68), .A2(G107), .ZN(new_n408));
  NAND2_X1  g0208(.A1(KEYINPUT68), .A2(G107), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n265), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n407), .B(new_n411), .C1(new_n297), .C2(new_n230), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n272), .ZN(new_n413));
  INV_X1    g0213(.A(G244), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n379), .B1(new_n280), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT67), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT67), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n379), .B(new_n417), .C1(new_n280), .C2(new_n414), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n413), .A2(G190), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n406), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n413), .A2(new_n416), .A3(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G200), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n406), .ZN(new_n424));
  INV_X1    g0224(.A(G179), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n413), .A2(new_n425), .A3(new_n416), .A4(new_n418), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n421), .A2(new_n285), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n294), .A2(new_n355), .A3(new_n397), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n319), .B(new_n321), .C1(new_n263), .C2(new_n264), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT22), .B1(new_n432), .B2(new_n220), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT22), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n213), .A2(new_n268), .A3(new_n434), .A4(G87), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT24), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT23), .ZN(new_n438));
  AND2_X1   g0238(.A1(KEYINPUT68), .A2(G107), .ZN(new_n439));
  NOR2_X1   g0239(.A1(KEYINPUT68), .A2(G107), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n441), .B2(G20), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n443));
  INV_X1    g0243(.A(G107), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n213), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n436), .A2(new_n437), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n437), .B1(new_n436), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n252), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT77), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT77), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n252), .C1(new_n448), .C2(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT79), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n363), .B2(G107), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT78), .B(KEYINPUT25), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n277), .A2(G1), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n255), .A2(new_n252), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G107), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n255), .A2(KEYINPUT79), .A3(new_n444), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n456), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G294), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n468), .C1(new_n297), .C2(new_n221), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n272), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n469), .A2(new_n272), .B1(G264), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n472), .A2(new_n279), .A3(G274), .A4(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n285), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(G179), .B2(new_n476), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n469), .A2(new_n272), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(G264), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n480), .A2(G190), .A3(new_n475), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n465), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G200), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n474), .B2(new_n475), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n466), .A2(new_n479), .B1(new_n454), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n363), .A2(G116), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n460), .B2(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G283), .ZN(new_n490));
  INV_X1    g0290(.A(G97), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n213), .B(new_n490), .C1(G33), .C2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n251), .A2(new_n214), .B1(G20), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n492), .A2(KEYINPUT20), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT20), .B1(new_n492), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n489), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n268), .A2(G264), .A3(G1698), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n268), .A2(G257), .A3(new_n296), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n265), .A2(G303), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n272), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n272), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n473), .A2(G270), .B1(new_n505), .B2(new_n472), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G200), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n498), .B(new_n508), .C1(new_n290), .C2(new_n507), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n509), .B(KEYINPUT76), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n497), .A2(G179), .A3(new_n503), .A4(new_n506), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n285), .B1(new_n503), .B2(new_n506), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n497), .A3(KEYINPUT21), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT21), .B1(new_n512), .B2(new_n497), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT75), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n414), .A2(G1698), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(G238), .B2(G1698), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n521), .A2(new_n265), .B1(new_n277), .B2(new_n493), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n272), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT73), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n272), .B2(new_n504), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n279), .A2(KEYINPUT73), .A3(G274), .A4(new_n471), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n272), .A2(new_n221), .A3(new_n471), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n523), .A2(new_n527), .A3(new_n425), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT74), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n523), .A2(new_n527), .A3(new_n529), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n285), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n319), .A2(new_n321), .A3(G33), .A4(G97), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G87), .A2(G97), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n408), .A2(new_n537), .A3(new_n409), .ZN(new_n538));
  NAND3_X1  g0338(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n319), .A2(new_n321), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n213), .A2(new_n268), .A3(G68), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n536), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n252), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n404), .A2(new_n255), .ZN(new_n545));
  INV_X1    g0345(.A(new_n404), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n460), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n528), .B1(new_n522), .B2(new_n272), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT74), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n425), .A4(new_n527), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n531), .A2(new_n533), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n532), .A2(G200), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n549), .A2(G190), .A3(new_n527), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n543), .A2(new_n252), .B1(new_n255), .B2(new_n404), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n460), .A2(G87), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n519), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n552), .A2(new_n519), .A3(new_n557), .ZN(new_n560));
  OAI211_X1 g0360(.A(G244), .B(new_n296), .C1(new_n263), .C2(new_n264), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n490), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G250), .A2(G1698), .ZN(new_n565));
  NAND2_X1  g0365(.A1(KEYINPUT4), .A2(G244), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(G1698), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n268), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n272), .ZN(new_n570));
  AND2_X1   g0370(.A1(KEYINPUT5), .A2(G41), .ZN(new_n571));
  NOR2_X1   g0371(.A1(KEYINPUT5), .A2(G41), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n471), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(G257), .A3(new_n279), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n574), .A2(new_n475), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n570), .A2(new_n575), .A3(new_n290), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n279), .B1(new_n563), .B2(new_n568), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n475), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n484), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n363), .A2(G97), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n460), .B2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n333), .A2(new_n335), .A3(new_n410), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT6), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n585), .A2(G97), .A3(G107), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n491), .A2(KEYINPUT6), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n444), .A2(KEYINPUT72), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n444), .A2(KEYINPUT72), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n586), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g0390(.A(KEYINPUT72), .B(G107), .ZN(new_n591));
  INV_X1    g0391(.A(new_n587), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n491), .A2(new_n444), .A3(KEYINPUT6), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n594), .A3(new_n402), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n246), .A2(G77), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n584), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n583), .B1(new_n597), .B2(new_n252), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n580), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n570), .A2(new_n575), .A3(new_n425), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n285), .B1(new_n577), .B2(new_n578), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n598), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n559), .A2(new_n560), .A3(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n431), .A2(new_n487), .A3(new_n518), .A4(new_n605), .ZN(G372));
  NAND3_X1  g0406(.A1(new_n533), .A2(new_n548), .A3(new_n530), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n557), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n454), .B2(new_n486), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT80), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n514), .B2(new_n515), .ZN(new_n611));
  INV_X1    g0411(.A(new_n515), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(KEYINPUT80), .A3(new_n511), .A4(new_n513), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n464), .B1(new_n451), .B2(new_n453), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n478), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n604), .B(new_n609), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n603), .A2(new_n607), .A3(new_n557), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n607), .B1(new_n618), .B2(KEYINPUT26), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n559), .A2(new_n560), .A3(new_n603), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n431), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT81), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n352), .B2(new_n353), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n351), .A2(new_n338), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT18), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n351), .A2(KEYINPUT18), .A3(new_n338), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(KEYINPUT81), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT82), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n428), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n424), .A2(new_n427), .A3(KEYINPUT82), .A4(new_n426), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n395), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n391), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n343), .B(KEYINPUT17), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n625), .B(new_n630), .C1(new_n635), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n292), .A2(new_n293), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n286), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n623), .A2(new_n640), .ZN(G369));
  NAND2_X1  g0441(.A1(new_n213), .A2(new_n362), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n213), .A2(new_n644), .A3(new_n362), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n498), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT83), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n510), .B2(new_n516), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n510), .A2(new_n651), .A3(new_n516), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n650), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n614), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT84), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n654), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n656), .B1(new_n659), .B2(new_n652), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT84), .ZN(new_n661));
  INV_X1    g0461(.A(new_n657), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n466), .A2(new_n648), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n487), .A2(new_n665), .B1(new_n616), .B2(new_n648), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(G330), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n612), .A2(new_n511), .A3(new_n513), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n487), .A2(new_n669), .A3(new_n649), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n616), .A2(new_n649), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n210), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G1), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n441), .A2(new_n493), .A3(new_n537), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n678), .A2(new_n679), .B1(new_n215), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n518), .A2(new_n487), .A3(new_n605), .A4(new_n649), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n507), .A2(new_n425), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n570), .A2(new_n575), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n532), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n686), .A3(new_n474), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n684), .A2(new_n686), .A3(KEYINPUT30), .A4(new_n474), .ZN(new_n690));
  AOI21_X1  g0490(.A(G179), .B1(new_n549), .B2(new_n527), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n476), .A2(new_n507), .A3(new_n685), .A4(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n648), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT31), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n682), .B1(new_n683), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT26), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n618), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n552), .A2(new_n519), .A3(new_n557), .ZN(new_n700));
  AOI21_X1  g0500(.A(G169), .B1(new_n570), .B2(new_n575), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n577), .A2(new_n578), .A3(G179), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n597), .A2(new_n252), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n582), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n700), .A2(new_n558), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n699), .B1(new_n707), .B2(KEYINPUT26), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n516), .B1(new_n615), .B2(new_n478), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT85), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n580), .A2(new_n598), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n706), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n710), .B1(new_n706), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(new_n714), .A3(new_n609), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n708), .A2(new_n715), .A3(new_n607), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n649), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT86), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT86), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n669), .B1(new_n466), .B2(new_n479), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n436), .A2(new_n447), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT24), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n436), .A2(new_n437), .A3(new_n447), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n452), .B1(new_n724), .B2(new_n252), .ZN(new_n725));
  INV_X1    g0525(.A(new_n453), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n486), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT85), .B1(new_n599), .B2(new_n603), .ZN(new_n728));
  INV_X1    g0528(.A(new_n608), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n706), .A2(new_n710), .A3(new_n711), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n607), .B1(new_n720), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n698), .B1(new_n620), .B2(new_n697), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n719), .B(new_n649), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n718), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n648), .B1(new_n617), .B2(new_n621), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n696), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n681), .B1(new_n739), .B2(G1), .ZN(G364));
  NAND3_X1  g0540(.A1(new_n658), .A2(new_n682), .A3(new_n663), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n664), .A2(G330), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT87), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n402), .A2(new_n254), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n743), .B1(new_n678), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n677), .A2(KEYINPUT87), .A3(G1), .A4(new_n745), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n741), .A2(new_n742), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n675), .A2(new_n265), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n751), .A2(G355), .B1(new_n493), .B2(new_n675), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n675), .A2(new_n268), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G45), .B2(new_n215), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n243), .A2(new_n470), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(G20), .B1(KEYINPUT88), .B2(G169), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(KEYINPUT88), .A2(G169), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n214), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n756), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT89), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n213), .B1(new_n768), .B2(G190), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT91), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT91), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT92), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n770), .A2(KEYINPUT92), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n491), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n213), .A2(G190), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n425), .A3(G200), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT90), .Z(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G107), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n207), .A2(new_n290), .A3(new_n484), .A4(G179), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n213), .A2(new_n425), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n268), .B1(new_n784), .B2(new_n220), .C1(new_n787), .C2(new_n202), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n779), .A2(G179), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n788), .B1(G68), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n785), .A2(G190), .A3(new_n484), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G50), .A2(new_n793), .B1(new_n795), .B2(G58), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n779), .A2(new_n768), .ZN(new_n797));
  INV_X1    g0597(.A(G159), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT32), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n782), .A2(new_n791), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n778), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT93), .ZN(new_n804));
  XOR2_X1   g0604(.A(KEYINPUT33), .B(G317), .Z(new_n805));
  INV_X1    g0605(.A(G326), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n265), .B1(new_n789), .B2(new_n805), .C1(new_n806), .C2(new_n792), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G322), .B2(new_n795), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n781), .A2(G283), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n772), .A2(G294), .ZN(new_n810));
  INV_X1    g0610(.A(new_n797), .ZN(new_n811));
  INV_X1    g0611(.A(new_n787), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n811), .A2(G329), .B1(new_n812), .B2(G311), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n783), .B(KEYINPUT94), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G303), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n803), .A2(KEYINPUT93), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n804), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n765), .B(new_n749), .C1(new_n819), .C2(new_n760), .ZN(new_n820));
  INV_X1    g0620(.A(new_n763), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n664), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n750), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  INV_X1    g0624(.A(new_n749), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n406), .A2(new_n649), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n420), .B2(new_n422), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT96), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n428), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n424), .A2(new_n427), .A3(KEYINPUT96), .A4(new_n426), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(KEYINPUT97), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT97), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n827), .A2(new_n829), .A3(new_n834), .A4(new_n830), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n632), .A2(new_n633), .A3(new_n826), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n737), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n683), .A2(new_n695), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G330), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n825), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n842), .B2(new_n840), .ZN(new_n844));
  INV_X1    g0644(.A(new_n760), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n762), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n825), .B1(G77), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n790), .A2(G150), .B1(new_n812), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  INV_X1    g0649(.A(G143), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n848), .B1(new_n849), .B2(new_n792), .C1(new_n850), .C2(new_n794), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n772), .A2(G58), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n811), .A2(G132), .ZN(new_n856));
  INV_X1    g0656(.A(new_n814), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n268), .B(new_n856), .C1(new_n857), .C2(new_n258), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G68), .B2(new_n781), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n857), .A2(new_n444), .B1(new_n493), .B2(new_n787), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n268), .B(new_n861), .C1(G311), .C2(new_n811), .ZN(new_n862));
  AOI22_X1  g0662(.A1(G294), .A2(new_n795), .B1(new_n793), .B2(G303), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n790), .A2(KEYINPUT95), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n790), .A2(KEYINPUT95), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(G283), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n781), .A2(G87), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n862), .A2(new_n863), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n860), .B1(new_n870), .B2(new_n778), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n847), .B1(new_n871), .B2(new_n760), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n839), .B2(new_n762), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n844), .A2(new_n873), .ZN(G384));
  NOR3_X1   g0674(.A1(new_n213), .A2(new_n493), .A3(new_n214), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n590), .A2(new_n594), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT35), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n877), .B2(new_n876), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  OR2_X1    g0680(.A1(new_n215), .A2(new_n202), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n326), .A2(new_n328), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n881), .A2(new_n882), .B1(G50), .B2(new_n218), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(G1), .A3(new_n254), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT98), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n736), .A2(new_n431), .A3(new_n738), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n640), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n646), .B(KEYINPUT99), .Z(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n625), .B2(new_n630), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n372), .A2(new_n648), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n391), .A2(new_n395), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n378), .B1(new_n377), .B2(new_n381), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n383), .A2(KEYINPUT13), .A3(new_n380), .ZN(new_n894));
  OAI21_X1  g0694(.A(G169), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT14), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n388), .A3(new_n387), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n372), .B(new_n648), .C1(new_n897), .C2(new_n394), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n737), .A2(new_n839), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n829), .A2(new_n830), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n648), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n900), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT16), .B1(new_n324), .B2(new_n330), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n316), .B1(new_n332), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n646), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n354), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n338), .A2(new_n889), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n626), .A2(new_n343), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n311), .B2(new_n339), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n907), .B1(new_n351), .B2(new_n908), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n912), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n890), .B1(new_n905), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n897), .A2(new_n372), .A3(new_n649), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n920), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n916), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n625), .A2(new_n630), .A3(new_n636), .ZN(new_n927));
  INV_X1    g0727(.A(new_n911), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n343), .A2(new_n911), .A3(new_n624), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT37), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n912), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n343), .A2(new_n911), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n933), .A2(KEYINPUT81), .A3(KEYINPUT37), .A4(new_n626), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n926), .B1(new_n936), .B2(new_n918), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n924), .B(new_n925), .C1(new_n937), .C2(KEYINPUT39), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n922), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n888), .B(new_n939), .Z(new_n940));
  OAI21_X1  g0740(.A(new_n899), .B1(new_n832), .B2(new_n837), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n683), .B2(new_n695), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n929), .B2(new_n935), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n943), .B2(new_n926), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT40), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT40), .B1(new_n919), .B2(new_n920), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n942), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n430), .B1(new_n683), .B2(new_n695), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n682), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n940), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n206), .B2(new_n744), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n940), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n886), .B1(new_n953), .B2(new_n954), .ZN(G367));
  NAND2_X1  g0755(.A1(new_n705), .A2(new_n648), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n714), .A2(new_n956), .B1(new_n603), .B2(new_n648), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n668), .A2(KEYINPUT102), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT102), .B1(new_n668), .B2(new_n957), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n670), .A2(new_n957), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n714), .A2(new_n616), .A3(new_n956), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n648), .B1(new_n963), .B2(new_n706), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(KEYINPUT42), .B2(new_n961), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT101), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n649), .B1(new_n555), .B2(new_n556), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n607), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n729), .B2(new_n968), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT100), .Z(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT43), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n966), .A2(KEYINPUT101), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n967), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n967), .B2(new_n973), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n960), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n977), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n979), .A2(new_n974), .B1(new_n959), .B2(new_n958), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  INV_X1    g0782(.A(new_n957), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n673), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT44), .B1(new_n672), .B2(new_n957), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n672), .A2(new_n957), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n986), .A2(new_n668), .A3(new_n988), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n990), .A2(new_n991), .B1(new_n984), .B2(new_n985), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n682), .B(new_n666), .C1(new_n658), .C2(new_n663), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n666), .B1(new_n516), .B2(new_n648), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n670), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n742), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n739), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT103), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n676), .B(KEYINPUT41), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n746), .A2(new_n206), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1000), .B1(new_n999), .B2(new_n1001), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n981), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n753), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n236), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n764), .B1(new_n210), .B2(new_n404), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n825), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n867), .A2(G294), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n772), .A2(new_n410), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n783), .A2(G116), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT46), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n268), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(G303), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1015), .B1(new_n491), .B2(new_n780), .C1(new_n1016), .C2(new_n794), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(KEYINPUT104), .B(G311), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1017), .B1(new_n793), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  INV_X1    g0821(.A(G283), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n797), .A2(new_n1021), .B1(new_n787), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1014), .A2(new_n493), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1023), .B1(new_n814), .B2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1011), .A2(new_n1012), .A3(new_n1020), .A4(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n866), .A2(new_n798), .B1(new_n258), .B2(new_n787), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT105), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n265), .B1(new_n783), .B2(G58), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n797), .B2(new_n849), .C1(new_n202), .C2(new_n780), .ZN(new_n1031));
  INV_X1    g0831(.A(G150), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n850), .A2(new_n792), .B1(new_n794), .B2(new_n1032), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n777), .A2(new_n218), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1026), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT47), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1010), .B1(new_n1038), .B2(new_n760), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n821), .B2(new_n971), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1006), .A2(new_n1040), .ZN(G387));
  NAND3_X1  g0841(.A1(new_n742), .A2(new_n670), .A3(new_n996), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n664), .A2(G330), .A3(new_n997), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1003), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n781), .A2(G97), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n265), .B1(new_n783), .B2(G77), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n1032), .C2(new_n797), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT106), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n777), .A2(new_n404), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n790), .A2(new_n401), .B1(new_n812), .B2(G68), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n258), .B2(new_n794), .C1(new_n798), .C2(new_n792), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n268), .B1(new_n811), .B2(G326), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n793), .A2(G322), .B1(new_n812), .B2(G303), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n1021), .B2(new_n794), .C1(new_n866), .C2(new_n1018), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT48), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n772), .A2(G283), .B1(G294), .B2(new_n783), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT49), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1054), .B1(new_n493), .B2(new_n780), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1053), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n845), .B1(new_n1065), .B2(KEYINPUT107), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT107), .B2(new_n1065), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n233), .A2(new_n470), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1068), .A2(new_n753), .B1(new_n679), .B2(new_n751), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n401), .A2(new_n258), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT50), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n470), .B1(new_n218), .B2(new_n202), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1071), .A2(new_n679), .A3(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1069), .A2(new_n1073), .B1(G107), .B2(new_n210), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1074), .A2(new_n764), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n749), .B(new_n1075), .C1(new_n666), .C2(new_n763), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1044), .A2(new_n1045), .B1(new_n1067), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1044), .A2(new_n739), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n676), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1044), .A2(new_n739), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT108), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(KEYINPUT108), .B(new_n1077), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(G393));
  NOR2_X1   g0888(.A1(new_n1078), .A2(new_n995), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(new_n677), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1078), .A2(new_n995), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1007), .A2(new_n240), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n764), .B1(new_n491), .B2(new_n210), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G311), .A2(new_n795), .B1(new_n793), .B2(G317), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  INV_X1    g0896(.A(G294), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n265), .B1(new_n784), .B2(new_n1022), .C1(new_n787), .C2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G322), .B2(new_n811), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n782), .B(new_n1099), .C1(new_n1016), .C2(new_n866), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1096), .B(new_n1100), .C1(G116), .C2(new_n772), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n776), .A2(G77), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n258), .B2(new_n866), .C1(new_n248), .C2(new_n787), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT110), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n265), .B1(new_n783), .B2(G68), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n869), .B(new_n1105), .C1(new_n850), .C2(new_n797), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1032), .A2(new_n792), .B1(new_n794), .B2(new_n798), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1101), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n825), .B1(new_n1093), .B2(new_n1094), .C1(new_n1111), .C2(new_n845), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT111), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1114), .B(new_n1115), .C1(new_n821), .C2(new_n983), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n995), .B2(new_n1003), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT112), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1092), .B1(new_n1119), .B2(new_n1120), .ZN(G390));
  OAI21_X1  g0921(.A(new_n925), .B1(new_n937), .B2(KEYINPUT39), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n903), .B1(new_n737), .B2(new_n839), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n923), .B1(new_n1123), .B2(new_n900), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n734), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n719), .B1(new_n716), .B2(new_n649), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n839), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n900), .B1(new_n1128), .B2(new_n904), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n937), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n923), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n696), .A2(new_n839), .A3(new_n899), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n696), .A2(new_n839), .A3(new_n899), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1125), .B(new_n1135), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT113), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n839), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n900), .B1(new_n842), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1123), .B1(new_n1140), .B2(new_n1135), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n903), .B1(new_n735), .B2(new_n839), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n899), .B1(new_n696), .B2(new_n839), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1133), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1141), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n431), .A2(new_n696), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n887), .A2(new_n640), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1138), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n677), .B1(new_n1137), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1137), .B2(new_n1148), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1122), .A2(new_n761), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n825), .B1(new_n401), .B2(new_n846), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n857), .A2(new_n220), .B1(new_n1097), .B2(new_n797), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n268), .B(new_n1153), .C1(G97), .C2(new_n812), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n781), .A2(G68), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G116), .A2(new_n795), .B1(new_n793), .B2(G283), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n867), .A2(new_n410), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1102), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n777), .A2(new_n798), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n783), .A2(G150), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n265), .B1(new_n1161), .B2(KEYINPUT53), .ZN(new_n1162));
  INV_X1    g0962(.A(G132), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1162), .B1(KEYINPUT53), .B2(new_n1161), .C1(new_n1163), .C2(new_n794), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G128), .B2(new_n793), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n780), .A2(new_n258), .B1(new_n797), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT114), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n812), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1165), .B(new_n1170), .C1(new_n849), .C2(new_n866), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1158), .A2(new_n1159), .B1(new_n1160), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1152), .B1(new_n1172), .B2(new_n760), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT115), .Z(new_n1174));
  AOI22_X1  g0974(.A1(new_n1137), .A2(new_n1045), .B1(new_n1151), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1150), .A2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(KEYINPUT121), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n939), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n262), .A2(new_n646), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n294), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n294), .A2(new_n1182), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n294), .A2(new_n1182), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n294), .A2(new_n1182), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n1179), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n948), .B2(G330), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n944), .A2(KEYINPUT40), .B1(new_n942), .B2(new_n946), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1191), .A2(new_n682), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1178), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n948), .A2(G330), .A3(new_n1189), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1192), .B1(new_n1191), .B2(new_n682), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n939), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1003), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n825), .B1(G50), .B2(new_n846), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n779), .A2(G58), .A3(new_n425), .A4(G200), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT116), .Z(new_n1201));
  OAI22_X1  g1001(.A1(new_n797), .A2(new_n1022), .B1(new_n787), .B2(new_n404), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G41), .B(new_n268), .C1(new_n783), .C2(G77), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n491), .B2(new_n789), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(G107), .C2(new_n795), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1036), .B1(G116), .B2(new_n793), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1206), .A2(KEYINPUT117), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(KEYINPUT117), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1201), .B(new_n1205), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT58), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G33), .A2(G41), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G50), .B(new_n1213), .C1(new_n265), .C2(new_n278), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G125), .A2(new_n793), .B1(new_n795), .B2(G128), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n790), .A2(G132), .B1(new_n783), .B2(new_n1169), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n849), .C2(new_n787), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n776), .B2(G150), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT119), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(G124), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1213), .B1(new_n797), .B2(new_n1222), .C1(new_n798), .C2(new_n780), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1214), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1211), .A2(new_n1212), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1199), .B1(new_n1226), .B2(new_n760), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1192), .A2(new_n761), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1198), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1144), .A2(new_n1142), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1123), .B2(new_n1144), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1134), .A2(new_n1136), .A3(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1147), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT120), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(KEYINPUT120), .A3(new_n1236), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT57), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n677), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1195), .A2(new_n1196), .A3(new_n939), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n939), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1235), .A2(KEYINPUT120), .A3(new_n1236), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT120), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1242), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1177), .B(new_n1232), .C1(new_n1244), .C2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1243), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1247), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n676), .B(new_n1254), .C1(new_n1255), .C2(KEYINPUT57), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT121), .B1(new_n1256), .B2(new_n1231), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1253), .A2(new_n1257), .ZN(G375));
  OAI21_X1  g1058(.A(new_n825), .B1(G68), .B2(new_n846), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n867), .A2(G116), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n797), .A2(new_n1016), .B1(new_n787), .B2(new_n441), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n268), .B(new_n1261), .C1(G97), .C2(new_n814), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G283), .A2(new_n795), .B1(new_n793), .B2(G294), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n781), .A2(G77), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1260), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n777), .A2(new_n258), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n867), .A2(new_n1169), .ZN(new_n1267));
  INV_X1    g1067(.A(G128), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n797), .A2(new_n1268), .B1(new_n787), .B2(new_n1032), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n265), .B(new_n1269), .C1(G159), .C2(new_n814), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G132), .A2(new_n793), .B1(new_n795), .B2(G137), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1267), .A2(new_n1201), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1050), .A2(new_n1265), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1259), .B1(new_n1273), .B2(new_n760), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n762), .B2(new_n899), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1145), .B2(new_n1003), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1001), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1276), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(G381));
  NAND3_X1  g1081(.A1(new_n1083), .A2(new_n823), .A3(new_n1085), .ZN(new_n1282));
  OR4_X1    g1082(.A1(G384), .A2(G390), .A3(new_n1282), .A4(G381), .ZN(new_n1283));
  OR4_X1    g1083(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1283), .ZN(G407));
  NAND2_X1  g1084(.A1(new_n647), .A2(G213), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT122), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G378), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G407), .B(G213), .C1(new_n1287), .C2(new_n1289), .ZN(G409));
  INV_X1    g1090(.A(G390), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G387), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n823), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1006), .A2(G390), .A3(new_n1040), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1292), .A2(new_n1282), .A3(new_n1294), .A4(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1282), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1006), .A2(G390), .A3(new_n1040), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G390), .B1(new_n1006), .B2(new_n1040), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT57), .B1(new_n1241), .B2(new_n1248), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1254), .A2(new_n676), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G378), .B(new_n1231), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT123), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1198), .A2(new_n1305), .A3(new_n1230), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1045), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT123), .B1(new_n1307), .B2(new_n1229), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1001), .B(new_n1248), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1288), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1304), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1145), .A2(new_n1147), .A3(KEYINPUT60), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1314), .A2(new_n676), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT60), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1279), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1276), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  OR2_X1    g1122(.A1(new_n1318), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1313), .A2(new_n1287), .A3(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT125), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1313), .A2(KEYINPUT125), .A3(new_n1287), .A4(new_n1326), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT62), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1286), .A2(G2897), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1325), .A2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1332), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G378), .B1(new_n1310), .B2(new_n1309), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1232), .B1(new_n1244), .B2(new_n1252), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1338), .B2(G378), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1336), .B1(new_n1339), .B2(new_n1286), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT61), .ZN(new_n1341));
  AOI211_X1 g1141(.A(new_n1286), .B(new_n1325), .C1(new_n1304), .C2(new_n1312), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1340), .B(new_n1341), .C1(new_n1342), .C2(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1301), .B1(new_n1331), .B2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT63), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1329), .A2(new_n1346), .A3(new_n1330), .ZN(new_n1347));
  AND2_X1   g1147(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1301), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1342), .A2(KEYINPUT63), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1347), .A2(new_n1348), .A3(new_n1349), .A4(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1345), .A2(new_n1351), .ZN(G405));
  AND2_X1   g1152(.A1(new_n1325), .A2(KEYINPUT126), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1256), .A2(new_n1231), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1177), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1338), .A2(KEYINPUT121), .ZN(new_n1356));
  AOI21_X1  g1156(.A(G378), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1338), .A2(new_n1288), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1353), .B1(new_n1357), .B2(new_n1358), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1325), .A2(KEYINPUT126), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1358), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1360), .B1(new_n1289), .B2(new_n1361), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1359), .B1(new_n1362), .B2(new_n1353), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1301), .B(KEYINPUT127), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT127), .ZN(new_n1366));
  XNOR2_X1  g1166(.A(new_n1301), .B(new_n1366), .ZN(new_n1367));
  OAI211_X1 g1167(.A(new_n1367), .B(new_n1359), .C1(new_n1353), .C2(new_n1362), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1365), .A2(new_n1368), .ZN(G402));
endmodule


