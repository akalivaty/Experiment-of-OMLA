//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n229), .B(new_n232), .Z(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G200), .ZN(new_n241));
  NAND2_X1  g0041(.A1(G33), .A2(G41), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT64), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G33), .A3(G41), .ZN(new_n245));
  INV_X1    g0045(.A(new_n214), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G45), .ZN(new_n249));
  AOI21_X1  g0049(.A(G1), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n247), .A2(G232), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT76), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n214), .B1(KEYINPUT64), .B2(new_n242), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n250), .B1(new_n255), .B2(new_n245), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(KEYINPUT76), .A3(G232), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n260), .A2(new_n262), .A3(G226), .A4(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n260), .A2(new_n262), .A3(G223), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G87), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n255), .B2(new_n245), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n267), .A2(new_n268), .B1(new_n270), .B2(new_n250), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n241), .B1(new_n258), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n260), .A2(new_n262), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT7), .B1(new_n274), .B2(new_n206), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT7), .ZN(new_n276));
  AOI211_X1 g0076(.A(new_n276), .B(G20), .C1(new_n260), .C2(new_n262), .ZN(new_n277));
  OAI21_X1  g0077(.A(G68), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT74), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n206), .A2(new_n259), .ZN(new_n280));
  INV_X1    g0080(.A(G159), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(KEYINPUT74), .A3(G159), .ZN(new_n284));
  XNOR2_X1  g0084(.A(G58), .B(G68), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n282), .A2(new_n284), .B1(new_n285), .B2(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n278), .A2(KEYINPUT16), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n288));
  INV_X1    g0088(.A(G68), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n276), .B1(new_n290), .B2(G20), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n282), .A2(new_n284), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n285), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n288), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n214), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n287), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n205), .B2(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(new_n299), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n302), .A2(new_n305), .B1(new_n301), .B2(new_n304), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n258), .A2(G190), .A3(new_n271), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n273), .A2(new_n300), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT17), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(KEYINPUT78), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n306), .ZN(new_n311));
  INV_X1    g0111(.A(new_n299), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n278), .A2(new_n286), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n288), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n314), .B2(new_n287), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n258), .A2(new_n271), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n272), .B1(new_n317), .B2(G190), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n309), .A2(KEYINPUT78), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n309), .A2(KEYINPUT78), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n315), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n310), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n258), .A2(new_n325), .A3(new_n271), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n315), .A2(new_n327), .A3(KEYINPUT18), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT18), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n258), .A2(new_n325), .A3(new_n271), .ZN(new_n330));
  AOI21_X1  g0130(.A(G169), .B1(new_n258), .B2(new_n271), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n300), .A2(new_n306), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n329), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT77), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT18), .B1(new_n315), .B2(new_n327), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT77), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n333), .A3(new_n329), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n322), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n283), .A2(G50), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT73), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n206), .A2(G33), .ZN(new_n343));
  INV_X1    g0143(.A(G77), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(new_n206), .B2(G68), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n299), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT11), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n347), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n303), .A2(KEYINPUT70), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT70), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n351), .A2(new_n205), .A3(G13), .A4(G20), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n299), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(G68), .C1(G1), .C2(new_n206), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n352), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT12), .B1(new_n355), .B2(G68), .ZN(new_n356));
  INV_X1    g0156(.A(G13), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(G1), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT12), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(G20), .A4(new_n289), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n348), .A2(new_n349), .A3(new_n354), .A4(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(G238), .A2(new_n256), .B1(new_n270), .B2(new_n250), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n260), .A2(new_n262), .A3(G232), .A4(G1698), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n260), .A2(new_n262), .A3(G226), .A4(new_n264), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G97), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT72), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n367), .A2(new_n368), .A3(new_n268), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n367), .B2(new_n268), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n363), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT13), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT13), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n363), .C1(new_n369), .C2(new_n370), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT14), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(G169), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(G179), .A3(new_n374), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n375), .B2(G169), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n362), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n290), .A2(G232), .A3(new_n264), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n290), .A2(G238), .A3(G1698), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT65), .B(G107), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n274), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT66), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n382), .A2(new_n383), .A3(new_n385), .A4(KEYINPUT66), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n268), .A3(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(G244), .A2(new_n256), .B1(new_n270), .B2(new_n250), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(KEYINPUT67), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT67), .B1(new_n390), .B2(new_n391), .ZN(new_n394));
  OAI21_X1  g0194(.A(G190), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n394), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(G200), .A3(new_n392), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G20), .A2(G77), .ZN(new_n398));
  XNOR2_X1  g0198(.A(KEYINPUT15), .B(G87), .ZN(new_n399));
  XOR2_X1   g0199(.A(KEYINPUT8), .B(G58), .Z(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(KEYINPUT68), .B2(new_n283), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n398), .B1(new_n343), .B2(new_n399), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n299), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT69), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT69), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(new_n406), .A3(new_n299), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n355), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n344), .B1(new_n205), .B2(G20), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n409), .A2(new_n344), .B1(new_n353), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n395), .A2(new_n397), .A3(new_n408), .A4(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n325), .B1(new_n393), .B2(new_n394), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n396), .A2(new_n323), .A3(new_n392), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n408), .A2(new_n411), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n340), .B(new_n381), .C1(KEYINPUT71), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(KEYINPUT71), .ZN(new_n419));
  INV_X1    g0219(.A(G150), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n301), .A2(new_n343), .B1(new_n420), .B2(new_n280), .ZN(new_n421));
  INV_X1    g0221(.A(G50), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n206), .B1(new_n201), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n299), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n422), .B1(new_n205), .B2(G20), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n305), .A2(new_n425), .B1(new_n422), .B2(new_n304), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT9), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n424), .A2(KEYINPUT9), .A3(new_n426), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n290), .A2(G222), .A3(new_n264), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n290), .A2(G223), .A3(G1698), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n344), .C2(new_n290), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n268), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n270), .A2(new_n250), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n256), .A2(G226), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n435), .A2(G190), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G200), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n431), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT10), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT10), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n431), .A2(new_n443), .A3(new_n438), .A4(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n439), .A2(new_n323), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n427), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n439), .A2(G179), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n372), .A2(new_n374), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n362), .B1(new_n451), .B2(G190), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n375), .A2(G200), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n419), .A2(new_n445), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n418), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT81), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT81), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT5), .ZN(new_n461));
  AOI21_X1  g0261(.A(G41), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT82), .B1(new_n458), .B2(G41), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT82), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n249), .A2(G1), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n464), .A2(new_n270), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n462), .B2(new_n463), .ZN(new_n469));
  AOI211_X1 g0269(.A(KEYINPUT82), .B(G41), .C1(new_n459), .C2(new_n461), .ZN(new_n470));
  OAI211_X1 g0270(.A(G270), .B(new_n247), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n261), .A2(G33), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n473));
  OAI21_X1  g0273(.A(G303), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n260), .A2(new_n262), .A3(G264), .A4(G1698), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n260), .A2(new_n262), .A3(G257), .A4(new_n264), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT85), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n477), .A2(new_n478), .A3(new_n268), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n477), .B2(new_n268), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n468), .B(new_n471), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n482), .B(new_n206), .C1(G33), .C2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT20), .ZN(new_n485));
  INV_X1    g0285(.A(G116), .ZN(new_n486));
  AOI22_X1  g0286(.A1(KEYINPUT86), .A2(new_n485), .B1(new_n486), .B2(G20), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n487), .A3(new_n299), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(KEYINPUT86), .B2(new_n485), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n485), .A2(KEYINPUT86), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n484), .A2(new_n487), .A3(new_n299), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n486), .B1(new_n205), .B2(G33), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n409), .A2(new_n486), .B1(new_n353), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n323), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n481), .A2(KEYINPUT21), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT87), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n481), .A2(new_n498), .A3(new_n495), .A4(KEYINPUT21), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(G179), .B1(new_n479), .B2(new_n480), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n492), .A2(new_n494), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n471), .A2(new_n468), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT21), .B1(new_n481), .B2(new_n495), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n481), .A2(G200), .ZN(new_n507));
  INV_X1    g0307(.A(G190), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n507), .B(new_n502), .C1(new_n508), .C2(new_n481), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n500), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G264), .B(new_n247), .C1(new_n469), .C2(new_n470), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n260), .A2(new_n262), .A3(G250), .A4(new_n264), .ZN(new_n512));
  INV_X1    g0312(.A(G294), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n259), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n290), .A2(G257), .A3(G1698), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n268), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n325), .A3(new_n468), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n511), .A2(new_n468), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n323), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n290), .A2(new_n206), .A3(G87), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT22), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n290), .A2(new_n523), .A3(new_n206), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n526), .A2(G107), .B1(new_n486), .B2(new_n343), .ZN(new_n527));
  XOR2_X1   g0327(.A(KEYINPUT65), .B(G107), .Z(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G20), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n527), .B1(new_n529), .B2(KEYINPUT23), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n525), .A2(new_n530), .A3(KEYINPUT24), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT24), .B1(new_n525), .B2(new_n530), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n532), .A2(new_n533), .A3(new_n312), .ZN(new_n534));
  OAI211_X1 g0334(.A(KEYINPUT88), .B(KEYINPUT25), .C1(new_n303), .C2(G107), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n205), .A2(G33), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n303), .A2(new_n536), .A3(new_n214), .A4(new_n298), .ZN(new_n537));
  INV_X1    g0337(.A(G107), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n304), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g0339(.A(KEYINPUT88), .B(KEYINPUT25), .ZN(new_n540));
  OAI221_X1 g0340(.A(new_n535), .B1(new_n537), .B2(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n541), .B(KEYINPUT89), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n518), .B(new_n520), .C1(new_n534), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n542), .ZN(new_n544));
  INV_X1    g0344(.A(new_n533), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(new_n299), .A3(new_n531), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n517), .A2(G190), .A3(new_n468), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n519), .A2(G200), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n544), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(G257), .B(new_n247), .C1(new_n469), .C2(new_n470), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n468), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT80), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n260), .A2(new_n262), .A3(G244), .A4(new_n264), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n482), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G250), .A2(G1698), .ZN(new_n558));
  NAND2_X1  g0358(.A1(KEYINPUT4), .A2(G244), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(G1698), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n290), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(new_n561), .A3(KEYINPUT79), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n268), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT79), .B1(new_n556), .B2(new_n561), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n553), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n556), .A2(new_n561), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n568), .A2(KEYINPUT80), .A3(new_n268), .A4(new_n562), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n552), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n325), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n268), .A3(new_n562), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n468), .A3(new_n551), .ZN(new_n573));
  XNOR2_X1  g0373(.A(G97), .B(G107), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT6), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n538), .A2(KEYINPUT6), .A3(G97), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n578), .A2(new_n206), .B1(new_n344), .B2(new_n280), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n384), .B1(new_n275), .B2(new_n277), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n299), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n303), .A2(G97), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n537), .B2(new_n483), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n573), .A2(new_n323), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n571), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(G87), .A2(G97), .ZN(new_n589));
  NAND3_X1  g0389(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n528), .A2(new_n589), .B1(new_n206), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n260), .A2(new_n262), .A3(new_n206), .A4(G68), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n343), .A2(new_n483), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(KEYINPUT19), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n299), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n409), .A2(new_n399), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(new_n596), .C1(new_n399), .C2(new_n537), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n247), .A2(G274), .A3(new_n467), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n270), .A2(KEYINPUT83), .A3(new_n467), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n260), .A2(new_n262), .A3(G244), .A4(G1698), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n260), .A2(new_n262), .A3(G238), .A4(new_n264), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n604), .C1(new_n259), .C2(new_n486), .ZN(new_n605));
  INV_X1    g0405(.A(G250), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n467), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n605), .A2(new_n268), .B1(new_n247), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(new_n608), .A3(new_n325), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n597), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n602), .A2(new_n608), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n323), .ZN(new_n612));
  INV_X1    g0412(.A(G87), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n537), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n595), .A2(new_n596), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n611), .B2(G200), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n602), .A2(new_n608), .A3(G190), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n610), .A2(new_n612), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n552), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(G190), .A3(new_n572), .ZN(new_n620));
  OAI221_X1 g0420(.A(new_n580), .B1(new_n344), .B2(new_n280), .C1(new_n206), .C2(new_n578), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n585), .B1(new_n621), .B2(new_n299), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n620), .B(new_n622), .C1(new_n570), .C2(new_n241), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n588), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT84), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT84), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n588), .A2(new_n618), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR4_X1   g0428(.A1(new_n457), .A2(new_n510), .A3(new_n550), .A4(new_n628), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n336), .A2(new_n338), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n416), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n454), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n381), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n631), .B1(new_n634), .B2(new_n322), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n449), .B1(new_n635), .B2(new_n445), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n612), .A2(new_n609), .A3(new_n597), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT90), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n610), .A2(KEYINPUT90), .A3(new_n612), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n616), .A2(new_n617), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n571), .A2(new_n587), .A3(new_n642), .A4(new_n637), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n618), .A2(new_n645), .A3(new_n571), .A4(new_n587), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n500), .A2(new_n506), .A3(new_n543), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n588), .A2(new_n618), .A3(new_n623), .A4(new_n549), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n644), .B(new_n646), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n636), .B1(new_n457), .B2(new_n651), .ZN(G369));
  NAND2_X1  g0452(.A1(new_n500), .A2(new_n506), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n358), .A2(new_n206), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n502), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n510), .B2(new_n661), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n543), .A2(new_n659), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n659), .B1(new_n534), .B2(new_n542), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n549), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n543), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n663), .A2(G330), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT91), .Z(new_n669));
  AOI211_X1 g0469(.A(new_n505), .B(new_n504), .C1(new_n497), .C2(new_n499), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n659), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n664), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(G399));
  INV_X1    g0473(.A(new_n209), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n528), .A2(new_n486), .A3(new_n589), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n212), .B2(new_n676), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n650), .A2(new_n682), .A3(new_n660), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n650), .B2(new_n660), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n543), .A2(new_n549), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n670), .A2(new_n686), .A3(new_n509), .A4(new_n660), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n628), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n471), .A2(new_n511), .A3(new_n468), .A4(new_n516), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(new_n611), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n477), .A2(new_n268), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT85), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n477), .A2(new_n478), .A3(new_n268), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n325), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n619), .A2(new_n695), .A3(new_n572), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n689), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n565), .A2(new_n569), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n619), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n519), .A2(new_n611), .A3(new_n325), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n481), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n573), .A2(new_n501), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n690), .A2(new_n611), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(KEYINPUT30), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n697), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n659), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(G330), .B1(new_n688), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT92), .B1(new_n685), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n650), .A2(new_n660), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT29), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n650), .A2(new_n682), .A3(new_n660), .ZN(new_n715));
  AND4_X1   g0515(.A1(KEYINPUT92), .A2(new_n711), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n681), .B1(new_n718), .B2(G1), .ZN(G364));
  NAND2_X1  g0519(.A1(new_n663), .A2(G330), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n357), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n205), .B1(new_n722), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n675), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G330), .B2(new_n663), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n209), .A2(new_n290), .ZN(new_n728));
  INV_X1    g0528(.A(G355), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n728), .A2(new_n729), .B1(G116), .B2(new_n209), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n674), .A2(new_n290), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n249), .B2(new_n213), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n236), .A2(new_n249), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n214), .B1(G20), .B2(new_n323), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n725), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n206), .A2(new_n325), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(new_n508), .A3(G200), .ZN(new_n744));
  XOR2_X1   g0544(.A(KEYINPUT33), .B(G317), .Z(new_n745));
  NOR2_X1   g0545(.A1(G190), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G311), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n744), .A2(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n206), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n746), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n290), .B(new_n749), .C1(G329), .C2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n508), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n206), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n743), .A2(G190), .A3(new_n241), .ZN(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n755), .A2(new_n513), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n750), .A2(new_n508), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n758), .B1(G283), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G326), .A2(new_n763), .B1(new_n765), .B2(G303), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n753), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n764), .A2(new_n613), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n274), .B(new_n768), .C1(G107), .C2(new_n760), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT94), .Z(new_n770));
  NOR2_X1   g0570(.A1(new_n751), .A2(new_n281), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT93), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT32), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT32), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n744), .A2(new_n289), .B1(new_n747), .B2(new_n344), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G50), .B2(new_n763), .ZN(new_n776));
  INV_X1    g0576(.A(new_n755), .ZN(new_n777));
  INV_X1    g0577(.A(new_n756), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G97), .A2(new_n777), .B1(new_n778), .B2(G58), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n773), .A2(new_n774), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n767), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT95), .ZN(new_n782));
  INV_X1    g0582(.A(new_n739), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n781), .B2(KEYINPUT95), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n742), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n738), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n663), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n727), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(G396));
  NOR2_X1   g0589(.A1(new_n416), .A2(new_n659), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n415), .A2(new_n659), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n412), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(new_n792), .B2(new_n416), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n713), .B(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n725), .B1(new_n795), .B2(new_n711), .ZN(new_n796));
  INV_X1    g0596(.A(G330), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT31), .B1(new_n705), .B2(new_n659), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n510), .A2(new_n550), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n801), .A2(new_n625), .A3(new_n627), .A4(new_n660), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n797), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n794), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n725), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n806), .A2(new_n762), .B1(new_n744), .B2(new_n420), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT98), .ZN(new_n808));
  INV_X1    g0608(.A(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n809), .B2(new_n756), .C1(new_n281), .C2(new_n747), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT34), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n759), .A2(new_n289), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n274), .B1(new_n752), .B2(G132), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n422), .B2(new_n764), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(G58), .C2(new_n777), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n744), .A2(new_n817), .B1(new_n747), .B2(new_n486), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT96), .Z(new_n819));
  OAI22_X1  g0619(.A1(new_n756), .A2(new_n513), .B1(new_n764), .B2(new_n538), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n274), .B1(new_n755), .B2(new_n483), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(G303), .C2(new_n763), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n759), .A2(new_n613), .B1(new_n751), .B2(new_n748), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT97), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n819), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n783), .B1(new_n816), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n739), .A2(new_n736), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n805), .B(new_n826), .C1(new_n344), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT99), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n793), .A2(new_n737), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n796), .A2(new_n804), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G384));
  NOR2_X1   g0632(.A1(new_n722), .A2(new_n205), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n381), .A2(KEYINPUT100), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT100), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n835), .B(new_n362), .C1(new_n379), .C2(new_n380), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n362), .A2(new_n659), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n452), .B2(new_n453), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n379), .A2(new_n380), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n454), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n837), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n800), .A2(new_n802), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n793), .ZN(new_n845));
  INV_X1    g0645(.A(new_n657), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n333), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT101), .B1(new_n340), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n310), .A2(new_n321), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n337), .B1(new_n336), .B2(new_n338), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT101), .ZN(new_n853));
  INV_X1    g0653(.A(new_n847), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n332), .A2(new_n333), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(new_n847), .A3(new_n308), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n848), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n848), .A2(new_n855), .A3(KEYINPUT38), .A4(new_n858), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n845), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n854), .B1(new_n322), .B2(new_n630), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n857), .A2(KEYINPUT102), .A3(KEYINPUT37), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n864), .B(new_n865), .C1(new_n858), .C2(KEYINPUT102), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n860), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT40), .A4(new_n793), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n863), .A2(KEYINPUT40), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n456), .A2(new_n844), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(G330), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT103), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n861), .A2(KEYINPUT39), .A3(new_n862), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n862), .A2(new_n867), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n659), .B1(new_n834), .B2(new_n836), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n631), .A2(new_n846), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n861), .A2(new_n862), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n839), .A2(new_n842), .ZN(new_n884));
  INV_X1    g0684(.A(new_n790), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n793), .A2(new_n650), .A3(new_n660), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n882), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n456), .B1(new_n683), .B2(new_n684), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n636), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n889), .B(new_n891), .Z(new_n892));
  AOI21_X1  g0692(.A(new_n833), .B1(new_n875), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n875), .B2(new_n892), .ZN(new_n894));
  INV_X1    g0694(.A(new_n578), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(G116), .A3(new_n215), .A4(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  INV_X1    g0699(.A(G58), .ZN(new_n900));
  OAI21_X1  g0700(.A(G77), .B1(new_n900), .B2(new_n289), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n212), .A2(new_n901), .B1(G50), .B2(new_n289), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(G1), .A3(new_n357), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n894), .A2(new_n899), .A3(new_n903), .ZN(G367));
  INV_X1    g0704(.A(new_n615), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(new_n660), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n639), .B2(new_n640), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n618), .B2(new_n907), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n588), .B(new_n623), .C1(new_n622), .C2(new_n660), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n913), .A2(new_n543), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n659), .B1(new_n914), .B2(new_n588), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n667), .A2(new_n671), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n571), .A2(new_n587), .A3(new_n659), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(KEYINPUT105), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT105), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n667), .A2(new_n671), .ZN(new_n922));
  INV_X1    g0722(.A(new_n919), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n920), .A2(new_n924), .A3(KEYINPUT42), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT42), .B1(new_n920), .B2(new_n924), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n916), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n912), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n927), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n915), .B1(new_n931), .B2(new_n925), .ZN(new_n932));
  INV_X1    g0732(.A(new_n912), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT106), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n930), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n929), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n933), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n928), .A2(new_n912), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT106), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n936), .A2(new_n940), .B1(new_n669), .B2(new_n923), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n672), .A2(new_n919), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT45), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(KEYINPUT44), .B(new_n923), .C1(new_n917), .C2(new_n664), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT44), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n672), .B2(new_n919), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n944), .A2(new_n669), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n669), .B1(new_n944), .B2(new_n948), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n667), .B(new_n671), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n721), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n717), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n675), .B(KEYINPUT41), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n723), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n935), .B1(new_n930), .B2(new_n934), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n938), .A2(KEYINPUT106), .A3(new_n939), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n669), .A2(new_n923), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n941), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n731), .A2(new_n232), .ZN(new_n962));
  INV_X1    g0762(.A(new_n399), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n741), .B1(new_n674), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n805), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G303), .A2(new_n778), .B1(new_n763), .B2(G311), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT107), .Z(new_n967));
  OAI22_X1  g0767(.A1(new_n755), .A2(new_n528), .B1(new_n759), .B2(new_n483), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n274), .B1(new_n744), .B2(new_n513), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n747), .A2(new_n817), .B1(new_n751), .B2(new_n970), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n765), .A2(KEYINPUT46), .A3(G116), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT46), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n764), .B2(new_n486), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n290), .B1(new_n755), .B2(new_n289), .ZN(new_n977));
  INV_X1    g0777(.A(new_n744), .ZN(new_n978));
  INV_X1    g0778(.A(new_n747), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n978), .A2(G159), .B1(new_n979), .B2(G50), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT108), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n756), .A2(new_n420), .B1(new_n762), .B2(new_n809), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G77), .B2(new_n760), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(new_n981), .C2(new_n980), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n764), .A2(new_n900), .B1(new_n751), .B2(new_n806), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT109), .Z(new_n987));
  OAI22_X1  g0787(.A1(new_n967), .A2(new_n976), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT110), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT47), .Z(new_n990));
  OAI221_X1 g0790(.A(new_n965), .B1(new_n786), .B2(new_n910), .C1(new_n990), .C2(new_n783), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n961), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT111), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n961), .A2(KEYINPUT111), .A3(new_n991), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(G387));
  OAI21_X1  g0797(.A(new_n953), .B1(new_n712), .B2(new_n716), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n711), .A2(new_n714), .A3(new_n715), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT92), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n685), .A2(KEYINPUT92), .A3(new_n711), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n952), .B(new_n720), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n675), .A3(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n667), .A2(new_n786), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n731), .B1(new_n229), .B2(new_n249), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n678), .B2(new_n728), .ZN(new_n1008));
  AOI21_X1  g0808(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1009));
  OR3_X1    g0809(.A1(new_n301), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT50), .B1(new_n301), .B2(G50), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n678), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1008), .A2(new_n1012), .B1(new_n538), .B2(new_n674), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n725), .B1(new_n1013), .B2(new_n741), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n747), .A2(new_n289), .B1(new_n751), .B2(new_n420), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n274), .B(new_n1015), .C1(new_n400), .C2(new_n978), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n764), .A2(new_n344), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n756), .A2(new_n422), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n963), .C2(new_n777), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G159), .A2(new_n763), .B1(new_n760), .B2(G97), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n290), .B1(new_n752), .B2(G326), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n755), .A2(new_n817), .B1(new_n764), .B2(new_n513), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n978), .A2(G311), .B1(new_n979), .B2(G303), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n970), .B2(new_n756), .C1(new_n757), .C2(new_n762), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT112), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1022), .B1(new_n486), .B2(new_n759), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1021), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1014), .B1(new_n1033), .B2(new_n739), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n953), .A2(new_n724), .B1(new_n1006), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1005), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT113), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1005), .A2(new_n1038), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(G393));
  INV_X1    g0840(.A(new_n998), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n676), .B1(new_n951), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n998), .B1(new_n949), .B2(new_n950), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n951), .A2(new_n724), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n777), .A2(G116), .B1(new_n978), .B2(G303), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1046), .A2(KEYINPUT114), .B1(G294), .B2(new_n979), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT114), .B2(new_n1046), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT115), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n756), .A2(new_n748), .B1(new_n762), .B2(new_n970), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n274), .B1(new_n751), .B2(new_n757), .C1(new_n538), .C2(new_n759), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G283), .B2(new_n765), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1049), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n744), .A2(new_n422), .B1(new_n747), .B2(new_n301), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n274), .B(new_n1055), .C1(G143), .C2(new_n752), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n756), .A2(new_n281), .B1(new_n762), .B2(new_n420), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT51), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n755), .A2(new_n344), .B1(new_n759), .B2(new_n613), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G68), .B2(new_n765), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n783), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n732), .A2(new_n239), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n741), .B(new_n1063), .C1(G97), .C2(new_n674), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1062), .A2(new_n805), .A3(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n919), .B2(new_n786), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1044), .A2(new_n1045), .A3(new_n1066), .ZN(G390));
  NAND2_X1  g0867(.A1(new_n886), .A2(new_n885), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n880), .B1(new_n1068), .B2(new_n843), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n861), .A2(KEYINPUT39), .A3(new_n862), .ZN(new_n1071));
  AOI21_X1  g0871(.A(KEYINPUT39), .B1(new_n862), .B2(new_n867), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n803), .A2(new_n793), .A3(new_n843), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1069), .A2(new_n877), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(G330), .B(new_n793), .C1(new_n688), .C2(new_n710), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n884), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1069), .B1(new_n876), .B2(new_n879), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1069), .A2(new_n877), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1076), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n456), .A2(new_n803), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n890), .A2(new_n636), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1077), .A2(new_n884), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1068), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n1074), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1086), .B2(new_n1074), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1082), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n843), .B1(new_n803), .B2(new_n793), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1068), .B1(new_n1078), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1086), .A2(new_n1087), .A3(new_n1074), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1084), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1076), .A2(new_n1081), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(new_n675), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1076), .A2(new_n1081), .A3(new_n724), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n736), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n805), .B1(new_n301), .B2(new_n827), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G132), .A2(new_n778), .B1(new_n763), .B2(G128), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n422), .B2(new_n759), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n744), .A2(new_n806), .B1(new_n747), .B2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT116), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n765), .A2(G150), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n274), .B1(new_n752), .B2(G125), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n281), .B2(new_n755), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1102), .A2(new_n1105), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n978), .A2(new_n384), .B1(new_n979), .B2(G97), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n817), .B2(new_n762), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT117), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n755), .A2(new_n344), .B1(new_n756), .B2(new_n486), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT118), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n812), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n290), .B(new_n768), .C1(G294), .C2(new_n752), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1110), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1099), .B(new_n1100), .C1(new_n783), .C2(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1098), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1097), .A2(new_n1121), .ZN(G378));
  NAND2_X1  g0922(.A1(new_n445), .A2(new_n450), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n427), .A2(new_n846), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT55), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1123), .B(new_n1125), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1127));
  XOR2_X1   g0927(.A(new_n1126), .B(new_n1127), .Z(new_n1128));
  INV_X1    g0928(.A(new_n845), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT40), .B1(new_n883), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(G330), .B1(new_n868), .B2(new_n869), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1128), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n869), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n797), .B1(new_n1133), .B2(new_n877), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1128), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(KEYINPUT40), .C2(new_n863), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n889), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n889), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1128), .A2(new_n736), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(G33), .A2(G41), .ZN(new_n1143));
  AOI211_X1 g0943(.A(G50), .B(new_n1143), .C1(new_n274), .C2(new_n248), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n762), .A2(new_n486), .B1(new_n759), .B2(new_n900), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G107), .B2(new_n778), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G41), .B(new_n290), .C1(new_n978), .C2(G97), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n963), .A2(new_n979), .B1(new_n752), .B2(G283), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1017), .B1(G68), .B2(new_n777), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT58), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1144), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G150), .A2(new_n777), .B1(new_n763), .B2(G125), .ZN(new_n1153));
  INV_X1    g0953(.A(G128), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n756), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n764), .A2(new_n1103), .ZN(new_n1156));
  INV_X1    g0956(.A(G132), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n744), .A2(new_n1157), .B1(new_n747), .B2(new_n806), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n760), .A2(G159), .ZN(new_n1162));
  OR2_X1    g0962(.A1(KEYINPUT119), .A2(G124), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(KEYINPUT119), .A2(G124), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n752), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1161), .A2(new_n1162), .A3(new_n1165), .A4(new_n1143), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1152), .B1(new_n1151), .B2(new_n1150), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1168), .A2(new_n739), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n805), .B(new_n1169), .C1(new_n422), .C2(new_n827), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1141), .A2(new_n724), .B1(new_n1142), .B2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n889), .A2(new_n1136), .A3(new_n1132), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1132), .A2(new_n1136), .B1(new_n881), .B2(new_n888), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT57), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1096), .A2(new_n1085), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n675), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1096), .A2(new_n1085), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT57), .B1(new_n1141), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1171), .B1(new_n1176), .B2(new_n1178), .ZN(G375));
  OAI21_X1  g0979(.A(new_n724), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n744), .A2(new_n1103), .B1(new_n751), .B2(new_n1154), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n274), .B(new_n1181), .C1(G150), .C2(new_n979), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n755), .A2(new_n422), .B1(new_n756), .B2(new_n806), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G159), .B2(new_n765), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G132), .A2(new_n763), .B1(new_n760), .B2(G58), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n762), .A2(new_n513), .B1(new_n764), .B2(new_n483), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G283), .B2(new_n778), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n290), .B1(new_n978), .B2(G116), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n384), .A2(new_n979), .B1(new_n752), .B2(G303), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n777), .A2(new_n963), .B1(new_n760), .B2(G77), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n783), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n805), .B(new_n1193), .C1(new_n289), .C2(new_n827), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n843), .B2(new_n737), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1180), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n955), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1093), .A2(new_n1084), .A3(new_n1094), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1090), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(G381));
  INV_X1    g1001(.A(KEYINPUT122), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1045), .A2(new_n1066), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(new_n1197), .A3(new_n1200), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(G378), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1037), .A2(new_n788), .A3(new_n1039), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(G384), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT121), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT121), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n996), .A2(new_n1206), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1202), .B1(new_n1211), .B2(G375), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G378), .B(new_n1205), .C1(new_n994), .C2(new_n995), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n724), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1142), .A2(new_n1170), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1141), .A2(new_n1177), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n676), .B1(new_n1221), .B2(new_n1177), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1217), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1213), .A2(new_n1214), .A3(KEYINPUT122), .A4(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1212), .A2(new_n1224), .ZN(G407));
  INV_X1    g1025(.A(G213), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(G343), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(G378), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1223), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(G213), .B1(new_n1230), .B2(KEYINPUT123), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1230), .B2(KEYINPUT123), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G407), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(new_n1235), .A3(new_n1232), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(G409));
  OAI211_X1 g1037(.A(G378), .B(new_n1171), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1141), .A2(new_n1198), .A3(new_n1177), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1097), .B(new_n1121), .C1(new_n1239), .C2(new_n1217), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1093), .A2(new_n1084), .A3(KEYINPUT60), .A4(new_n1094), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1242), .A2(new_n675), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT60), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1199), .B1(new_n1095), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G384), .B1(new_n1246), .B2(new_n1197), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n831), .B(new_n1196), .C1(new_n1243), .C2(new_n1245), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1241), .A2(new_n1228), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT63), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1228), .A4(new_n1249), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1227), .A2(G2897), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT125), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1242), .A2(new_n675), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1090), .A2(KEYINPUT60), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n1199), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n831), .B1(new_n1259), .B2(new_n1196), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1246), .A2(G384), .A3(new_n1197), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1254), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1255), .A2(new_n1256), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1256), .B1(new_n1255), .B2(new_n1263), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1141), .A2(new_n1198), .A3(new_n1177), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G378), .B1(new_n1171), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1223), .B2(G378), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1266), .B1(new_n1269), .B2(new_n1227), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n992), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1039), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1038), .B1(new_n1005), .B2(new_n1035), .ZN(new_n1273));
  OAI21_X1  g1073(.A(G396), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1207), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G390), .B1(new_n1275), .B2(KEYINPUT111), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1204), .B1(new_n1274), .B2(new_n1207), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1271), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(G390), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n993), .B1(new_n1274), .B2(new_n1207), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1280), .B(new_n992), .C1(G390), .C2(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1278), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1252), .A2(new_n1253), .A3(new_n1270), .A4(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1278), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1241), .A2(new_n1228), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1288), .B2(new_n1266), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1289), .A2(KEYINPUT126), .A3(new_n1253), .A4(new_n1252), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1255), .A2(new_n1263), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT61), .B1(new_n1288), .B2(new_n1293), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1294), .B1(new_n1250), .B2(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1250), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1292), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1291), .A2(new_n1298), .ZN(G405));
  XNOR2_X1  g1099(.A(G375), .B(G378), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1249), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1300), .B(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1292), .ZN(G402));
endmodule


