//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n585, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1232, new_n1233,
    new_n1234;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g021(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2106), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n469), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n479), .A2(new_n470), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G124), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT70), .B1(new_n479), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT3), .B(G2104), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G126), .A4(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n470), .C1(new_n477), .C2(new_n478), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n495), .A2(new_n501), .A3(G138), .A4(new_n470), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G88), .ZN(new_n512));
  INV_X1    g087(.A(G75), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT72), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G75), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(G62), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G50), .A3(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n522), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n529), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n529), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(KEYINPUT74), .A2(G89), .ZN(new_n540));
  NAND2_X1  g115(.A1(KEYINPUT74), .A2(G89), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n523), .A2(new_n519), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n523), .A2(G51), .A3(G543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n539), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  AOI22_X1  g121(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n521), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n523), .A2(new_n519), .A3(G90), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n550));
  OAI211_X1 g125(.A(G52), .B(G543), .C1(new_n507), .C2(new_n506), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n548), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(G171));
  NAND3_X1  g130(.A1(new_n523), .A2(G43), .A3(G543), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(new_n510), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n519), .A2(G56), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n521), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT76), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT78), .ZN(new_n568));
  XNOR2_X1  g143(.A(KEYINPUT77), .B(KEYINPUT8), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT79), .Z(G188));
  INV_X1    g147(.A(G78), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n573), .A2(new_n514), .A3(KEYINPUT80), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT80), .B1(new_n573), .B2(new_n514), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n508), .A2(new_n509), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  INV_X1    g154(.A(G91), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(new_n510), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n523), .A2(G53), .A3(G543), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT9), .Z(new_n583));
  OR2_X1    g158(.A1(new_n581), .A2(new_n583), .ZN(G299));
  NAND2_X1  g159(.A1(new_n554), .A2(KEYINPUT81), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n548), .B(new_n586), .C1(new_n552), .C2(new_n553), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G301));
  NAND2_X1  g164(.A1(new_n511), .A2(G87), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n507), .A2(new_n506), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n514), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G49), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(G288));
  NAND3_X1  g170(.A1(new_n523), .A2(G48), .A3(G543), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  OAI221_X1 g173(.A(new_n596), .B1(new_n510), .B2(new_n597), .C1(new_n598), .C2(new_n521), .ZN(G305));
  AND2_X1   g174(.A1(new_n519), .A2(G60), .ZN(new_n600));
  AND2_X1   g175(.A1(G72), .A2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT82), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n604), .B(G651), .C1(new_n600), .C2(new_n601), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n511), .A2(G85), .B1(new_n592), .B2(G47), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(new_n592), .A2(G54), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n519), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n521), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OR3_X1    g186(.A1(new_n510), .A2(KEYINPUT84), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT84), .B1(new_n510), .B2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT83), .B1(new_n619), .B2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n588), .A2(new_n621), .ZN(new_n622));
  MUX2_X1   g197(.A(new_n620), .B(KEYINPUT83), .S(new_n622), .Z(G284));
  MUX2_X1   g198(.A(new_n620), .B(KEYINPUT83), .S(new_n622), .Z(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n581), .A2(new_n583), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n619), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n619), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g208(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n634));
  XNOR2_X1  g209(.A(G323), .B(new_n634), .ZN(G282));
  NAND2_X1  g210(.A1(new_n495), .A2(new_n471), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT13), .Z(new_n638));
  NAND2_X1  g213(.A1(KEYINPUT86), .A2(G2100), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n638), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(KEYINPUT86), .B2(G2100), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n640), .B1(new_n642), .B2(new_n639), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n481), .A2(KEYINPUT87), .A3(G135), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n475), .A2(new_n480), .ZN(new_n646));
  INV_X1    g221(.A(G135), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  INV_X1    g225(.A(G111), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(G2105), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n486), .B2(G123), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n654), .A2(G2096), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(G2096), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n643), .A2(new_n655), .A3(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT14), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2451), .B(G2454), .Z(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT88), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G14), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n667), .A2(new_n670), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(G401));
  XNOR2_X1  g249(.A(KEYINPUT92), .B(G2096), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2084), .B(G2090), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT89), .Z(new_n678));
  NOR2_X1   g253(.A1(G2072), .A2(G2078), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n444), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n680), .B(KEYINPUT17), .Z(new_n683));
  INV_X1    g258(.A(new_n681), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n678), .B(new_n682), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT90), .Z(new_n686));
  INV_X1    g261(.A(new_n678), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n683), .A2(new_n687), .A3(new_n684), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT91), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n687), .A2(new_n681), .A3(new_n680), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT18), .Z(new_n691));
  NAND3_X1  g266(.A1(new_n686), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G2100), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(G2100), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n676), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n675), .A3(new_n693), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(G227));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT95), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1971), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT19), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1956), .B(G2474), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G1961), .B(G1966), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n705), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n708), .A2(KEYINPUT94), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(KEYINPUT20), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n712), .A2(new_n716), .A3(new_n713), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G1981), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n710), .A2(new_n705), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n708), .A2(new_n709), .ZN(new_n721));
  MUX2_X1   g296(.A(new_n705), .B(new_n720), .S(new_n721), .Z(new_n722));
  NAND3_X1  g297(.A1(new_n718), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n719), .B1(new_n718), .B2(new_n722), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n703), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n725), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n727), .A2(G1986), .A3(new_n723), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n702), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(G1991), .B(G1996), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n726), .A2(new_n728), .A3(new_n702), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n731), .ZN(new_n734));
  INV_X1    g309(.A(new_n732), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n729), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n736), .ZN(G229));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G32), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n481), .A2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  NAND3_X1  g317(.A1(new_n495), .A2(G129), .A3(G2105), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n471), .A2(G105), .ZN(new_n744));
  AND3_X1   g319(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n738), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G34), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n751), .B2(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT24), .B2(new_n751), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n473), .B2(new_n738), .ZN(new_n754));
  INV_X1    g329(.A(G2084), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G28), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(KEYINPUT30), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(KEYINPUT30), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G19), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n562), .B2(G16), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1341), .Z(new_n765));
  NAND4_X1  g340(.A1(new_n750), .A2(new_n756), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n738), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n738), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT29), .Z(new_n769));
  INV_X1    g344(.A(G2090), .ZN(new_n770));
  INV_X1    g345(.A(G16), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n619), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G4), .B2(new_n771), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT98), .B(G1348), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n769), .A2(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n766), .B(new_n775), .C1(new_n773), .C2(new_n774), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT101), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n475), .A2(new_n480), .A3(G139), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(KEYINPUT100), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT100), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n475), .A2(new_n480), .A3(new_n780), .A4(G139), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT25), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n777), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n778), .A2(KEYINPUT100), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n786), .A2(KEYINPUT101), .A3(new_n781), .A4(new_n783), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n495), .A2(G127), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n470), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G33), .B(new_n793), .S(G29), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(new_n442), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n654), .A2(new_n738), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT102), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n771), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n626), .B2(new_n771), .ZN(new_n800));
  INV_X1    g375(.A(G1956), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n754), .A2(new_n755), .ZN(new_n803));
  NAND2_X1  g378(.A1(G286), .A2(G16), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n771), .A2(G21), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G1966), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n807), .B2(new_n806), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n797), .A2(new_n802), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n738), .A2(G26), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT28), .Z(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(G116), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n486), .B2(G128), .ZN(new_n816));
  INV_X1    g391(.A(G140), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n646), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT99), .B(G2067), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n738), .A2(G27), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G164), .B2(new_n738), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2078), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n771), .A2(G5), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G171), .B2(new_n771), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1961), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n810), .A2(new_n821), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n769), .A2(new_n770), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT103), .Z(new_n830));
  NAND4_X1  g405(.A1(new_n776), .A2(new_n795), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n738), .A2(G25), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n481), .A2(G131), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n834));
  INV_X1    g409(.A(G107), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(G2105), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n486), .B2(G119), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n832), .B1(new_n839), .B2(new_n738), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G1991), .Z(new_n841));
  XOR2_X1   g416(.A(new_n840), .B(new_n841), .Z(new_n842));
  AND2_X1   g417(.A1(new_n771), .A2(G24), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G290), .B2(G16), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n703), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n703), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n842), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n771), .A2(G22), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G166), .B2(new_n771), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G1971), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT34), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n771), .A2(G6), .ZN(new_n854));
  INV_X1    g429(.A(G305), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n771), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT32), .B(G1981), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n856), .B(new_n857), .Z(new_n858));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n771), .A2(G23), .ZN(new_n862));
  INV_X1    g437(.A(G288), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(new_n771), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT33), .B(G1976), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n860), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n852), .A2(new_n853), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G1971), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n851), .B(new_n869), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n860), .A2(new_n861), .A3(new_n866), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT34), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n847), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT36), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(KEYINPUT36), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n831), .B1(new_n874), .B2(new_n875), .ZN(G311));
  INV_X1    g451(.A(new_n831), .ZN(new_n877));
  INV_X1    g452(.A(new_n875), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n873), .A2(KEYINPUT36), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(G150));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n519), .A2(G67), .ZN(new_n882));
  NAND2_X1  g457(.A1(G80), .A2(G543), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n521), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n523), .A2(new_n519), .A3(G93), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n523), .A2(G55), .A3(G543), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n881), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G67), .ZN(new_n889));
  INV_X1    g464(.A(new_n509), .ZN(new_n890));
  NAND2_X1  g465(.A1(KEYINPUT5), .A2(G543), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n883), .ZN(new_n893));
  OAI21_X1  g468(.A(G651), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n894), .A2(KEYINPUT104), .A3(new_n886), .A4(new_n885), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n888), .A2(new_n562), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n886), .A3(new_n885), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(new_n881), .C1(new_n561), .C2(new_n558), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(KEYINPUT38), .Z(new_n900));
  NAND2_X1  g475(.A1(new_n619), .A2(G559), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n903), .A2(new_n904), .A3(G860), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n897), .A2(G860), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT37), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n905), .A2(new_n907), .ZN(G145));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  INV_X1    g485(.A(new_n818), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n740), .A3(new_n745), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n746), .A2(new_n818), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n788), .A3(new_n792), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n788), .B2(new_n792), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n504), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n793), .A2(new_n913), .A3(new_n912), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(G164), .A3(new_n915), .ZN(new_n920));
  OAI21_X1  g495(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n921));
  INV_X1    g496(.A(G118), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(G2105), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n486), .B2(G130), .ZN(new_n924));
  INV_X1    g499(.A(G142), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n646), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n926), .A2(new_n637), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n637), .ZN(new_n928));
  OR3_X1    g503(.A1(new_n927), .A2(new_n928), .A3(new_n838), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n838), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n918), .A2(new_n920), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n654), .A2(new_n488), .ZN(new_n935));
  NAND3_X1  g510(.A1(G162), .A2(new_n649), .A3(new_n653), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n473), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n473), .B1(new_n935), .B2(new_n936), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n936), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G160), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n937), .A3(new_n933), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n932), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n931), .B1(new_n918), .B2(new_n920), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n910), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n929), .A2(KEYINPUT107), .A3(new_n930), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n918), .A2(new_n920), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n918), .B2(new_n920), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n949), .A2(new_n950), .A3(new_n944), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n909), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n948), .ZN(new_n953));
  INV_X1    g528(.A(new_n920), .ZN(new_n954));
  AOI21_X1  g529(.A(G164), .B1(new_n919), .B2(new_n915), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n918), .A2(new_n920), .A3(new_n948), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n956), .A2(new_n957), .A3(new_n943), .A4(new_n940), .ZN(new_n958));
  INV_X1    g533(.A(new_n931), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n954), .B2(new_n955), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n944), .A3(new_n932), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n958), .A2(new_n961), .A3(KEYINPUT108), .A4(new_n910), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n952), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g539(.A1(G166), .A2(G305), .ZN(new_n965));
  NAND2_X1  g540(.A1(G303), .A2(new_n855), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(G290), .B(new_n863), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(G290), .B(G288), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n970), .A2(new_n965), .A3(new_n966), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT109), .Z(new_n974));
  NOR2_X1   g549(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n975), .B(KEYINPUT110), .Z(new_n976));
  INV_X1    g551(.A(new_n899), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n631), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n618), .A2(G299), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n626), .A2(new_n617), .A3(new_n616), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT41), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT41), .B1(new_n979), .B2(new_n980), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n978), .ZN(new_n988));
  AND4_X1   g563(.A1(new_n974), .A2(new_n976), .A3(new_n983), .A4(new_n988), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n976), .A2(new_n974), .B1(new_n983), .B2(new_n988), .ZN(new_n990));
  OAI21_X1  g565(.A(G868), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n897), .A2(new_n621), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(G295));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n992), .ZN(G331));
  OAI211_X1 g569(.A(G286), .B(new_n548), .C1(new_n552), .C2(new_n553), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT112), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n549), .A2(new_n551), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT75), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(G286), .A4(new_n548), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n585), .A2(G168), .A3(new_n587), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n899), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n982), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n899), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n977), .ZN(new_n1012));
  AOI211_X1 g587(.A(KEYINPUT113), .B(new_n899), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1005), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n985), .A2(new_n986), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1014), .A2(KEYINPUT114), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT114), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n969), .A2(KEYINPUT115), .A3(new_n971), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT115), .B1(new_n969), .B2(new_n971), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT43), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n972), .B(new_n1009), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n910), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1005), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(new_n1007), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1028));
  OAI22_X1  g603(.A1(new_n987), .A2(new_n1027), .B1(new_n1028), .B2(new_n1006), .ZN(new_n1029));
  AOI21_X1  g604(.A(G37), .B1(new_n1029), .B2(new_n1021), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1024), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT43), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1025), .A2(KEYINPUT44), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1011), .A2(new_n977), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT113), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1026), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1034), .B1(new_n1038), .B2(new_n987), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1014), .A2(new_n1015), .A3(KEYINPUT114), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1008), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1021), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1024), .B(new_n910), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT43), .B1(new_n1041), .B2(new_n972), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1043), .A2(KEYINPUT43), .B1(new_n1044), .B2(new_n1030), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1033), .B1(new_n1045), .B2(new_n1046), .ZN(G397));
  NAND3_X1  g622(.A1(new_n468), .A2(new_n472), .A3(G40), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n468), .A2(new_n472), .A3(KEYINPUT116), .A4(G40), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1384), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT45), .B1(new_n504), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(new_n746), .B(G1996), .Z(new_n1057));
  INV_X1    g632(.A(G2067), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n818), .B(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n838), .B(new_n841), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(G290), .B(G1986), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1056), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G1384), .B1(new_n498), .B2(new_n503), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1050), .B(new_n1051), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT122), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1068), .B2(KEYINPUT122), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n801), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n1074));
  XNOR2_X1  g649(.A(G299), .B(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n504), .A2(new_n1053), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT45), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1066), .A2(KEYINPUT45), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1052), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT124), .B(KEYINPUT56), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1081), .B(G2072), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1073), .B(new_n1075), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1348), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1068), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1050), .A2(new_n1066), .A3(new_n1051), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1058), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n618), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1083), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1075), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1072), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1956), .B1(new_n1093), .B2(new_n1069), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT61), .B1(new_n1096), .B2(new_n1083), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1086), .A2(new_n1089), .A3(new_n618), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT60), .B1(new_n1099), .B2(new_n1090), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n618), .A2(KEYINPUT60), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1086), .A2(new_n1089), .A3(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT58), .B(G1341), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1080), .A2(G1996), .B1(new_n1088), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n562), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1104), .B2(new_n562), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1100), .B(new_n1102), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1098), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1096), .A2(new_n1083), .A3(KEYINPUT61), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1097), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1076), .A2(KEYINPUT50), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1052), .A2(new_n1112), .A3(new_n755), .A4(new_n1071), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1077), .B(G1384), .C1(new_n498), .C2(new_n503), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1114), .A2(new_n1054), .A3(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1113), .B(G168), .C1(new_n1116), .C2(G1966), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1080), .A2(new_n807), .ZN(new_n1119));
  AOI21_X1  g694(.A(G168), .B1(new_n1119), .B2(new_n1113), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT51), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1117), .A2(new_n1122), .A3(G8), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1080), .B2(G2078), .ZN(new_n1126));
  INV_X1    g701(.A(G1961), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1068), .B2(new_n1085), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1048), .A2(new_n1125), .A3(G2078), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1078), .A2(new_n1079), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1124), .B1(new_n1131), .B2(G171), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1116), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1126), .A2(new_n1133), .A3(G301), .A4(new_n1128), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1121), .A2(new_n1123), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(G303), .A2(G8), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT55), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1052), .A2(new_n1112), .A3(new_n770), .A4(new_n1071), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1068), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1142), .A2(KEYINPUT117), .A3(new_n770), .A4(new_n1071), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1080), .A2(new_n869), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1138), .A2(new_n1145), .A3(G8), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1087), .A2(G8), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n598), .B2(new_n521), .ZN(new_n1149));
  NAND3_X1  g724(.A1(G305), .A2(G1981), .A3(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n598), .A2(new_n521), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n511), .A2(G86), .B1(new_n592), .B2(G48), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1151), .B(new_n1152), .C1(new_n1148), .C2(new_n719), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT49), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1147), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1150), .A2(new_n1153), .A3(KEYINPUT49), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n590), .A2(new_n593), .A3(G1976), .A4(new_n594), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT118), .ZN(new_n1162));
  INV_X1    g737(.A(G1976), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT52), .B1(G288), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1162), .A2(G8), .A3(new_n1087), .A4(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(G8), .A3(new_n1087), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT52), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1160), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1146), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1093), .A2(new_n770), .A3(new_n1069), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1144), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1138), .B1(new_n1171), .B2(G8), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1126), .A2(new_n1133), .A3(new_n1128), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n588), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1126), .A2(G301), .A3(new_n1130), .A4(new_n1128), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT125), .B1(new_n1177), .B2(new_n1124), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n1179));
  AOI211_X1 g754(.A(new_n1179), .B(KEYINPUT54), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1135), .B(new_n1173), .C1(new_n1178), .C2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1111), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n1183));
  INV_X1    g758(.A(G8), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(new_n1170), .B2(new_n1144), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1146), .B(new_n1168), .C1(new_n1185), .C2(new_n1138), .ZN(new_n1186));
  AOI211_X1 g761(.A(new_n1184), .B(G286), .C1(new_n1119), .C2(new_n1113), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1183), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1146), .A2(new_n1168), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1145), .A2(G8), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1137), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1190), .A2(KEYINPUT63), .A3(new_n1187), .A4(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1189), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(KEYINPUT62), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1175), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1121), .A2(new_n1198), .A3(new_n1123), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1196), .A2(new_n1173), .A3(new_n1197), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n863), .A2(new_n1163), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT121), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1160), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n855), .A2(new_n719), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1147), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1146), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1205), .B1(new_n1206), .B2(new_n1168), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1194), .A2(new_n1200), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1065), .B1(new_n1182), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1055), .B1(new_n747), .B2(new_n1059), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n1210), .B(KEYINPUT127), .Z(new_n1211));
  NOR2_X1   g786(.A1(new_n1055), .A2(G1996), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1212), .B(KEYINPUT46), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  XOR2_X1   g789(.A(new_n1214), .B(KEYINPUT47), .Z(new_n1215));
  NAND3_X1  g790(.A1(new_n1061), .A2(new_n841), .A3(new_n839), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n911), .A2(new_n1058), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1055), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  XOR2_X1   g793(.A(new_n1218), .B(KEYINPUT126), .Z(new_n1219));
  OR3_X1    g794(.A1(new_n1055), .A2(G1986), .A3(G290), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1220), .ZN(new_n1221));
  AOI22_X1  g796(.A1(new_n1063), .A2(new_n1056), .B1(KEYINPUT48), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1222), .B1(KEYINPUT48), .B2(new_n1221), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1215), .A2(new_n1219), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1209), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g800(.A(G319), .B1(new_n672), .B2(new_n673), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n696), .B2(new_n698), .ZN(new_n1228));
  AND3_X1   g802(.A1(new_n1228), .A2(new_n733), .A3(new_n736), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1229), .A2(new_n963), .ZN(new_n1230));
  NOR2_X1   g804(.A1(new_n1230), .A2(new_n1045), .ZN(G308));
  AND2_X1   g805(.A1(new_n1044), .A2(new_n1030), .ZN(new_n1232));
  AOI21_X1  g806(.A(G37), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1233));
  AOI21_X1  g807(.A(new_n1023), .B1(new_n1233), .B2(new_n1024), .ZN(new_n1234));
  OAI211_X1 g808(.A(new_n963), .B(new_n1229), .C1(new_n1232), .C2(new_n1234), .ZN(G225));
endmodule


