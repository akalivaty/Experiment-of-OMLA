//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n556, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  OR4_X1    g026(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g030(.A(G2105), .ZN(new_n456));
  XNOR2_X1  g031(.A(KEYINPUT3), .B(G2104), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G125), .ZN(new_n458));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT66), .B(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n464), .B(new_n466), .C1(new_n467), .C2(new_n465), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n461), .B1(new_n470), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n456), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(new_n456), .B2(G112), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  AND2_X1   g055(.A1(new_n464), .A2(new_n466), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n463), .A2(KEYINPUT66), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n463), .A2(KEYINPUT66), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT3), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(new_n484), .A3(G126), .ZN(new_n485));
  NAND2_X1  g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n456), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(KEYINPUT4), .A2(G138), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n481), .A2(new_n484), .A3(new_n456), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n457), .A2(G138), .A3(new_n456), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n456), .A2(G102), .A3(G2104), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n487), .A2(new_n493), .A3(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n497), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT68), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT69), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n497), .A2(new_n499), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n496), .B1(new_n504), .B2(new_n505), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(G651), .B1(G50), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n517), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n503), .A2(G89), .A3(new_n509), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n523), .B2(new_n526), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n521), .B(new_n522), .C1(new_n527), .C2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n510), .A2(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n515), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G651), .B1(G52), .B2(new_n517), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n515), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(KEYINPUT71), .A3(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n503), .A2(G81), .A3(new_n509), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n517), .A2(G43), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  XOR2_X1   g130(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n556));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G188));
  OAI211_X1 g134(.A(G53), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n506), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n564), .B1(new_n562), .B2(new_n563), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n503), .A2(G91), .A3(new_n509), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n497), .A2(new_n499), .A3(G65), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n569), .B1(new_n572), .B2(G651), .ZN(new_n573));
  INV_X1    g148(.A(G651), .ZN(new_n574));
  AOI211_X1 g149(.A(KEYINPUT75), .B(new_n574), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n568), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT76), .B1(new_n567), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT9), .B1(new_n517), .B2(G53), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n560), .A2(new_n561), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT74), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT75), .B1(new_n584), .B2(new_n574), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n572), .A2(new_n569), .A3(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n582), .A2(new_n583), .A3(new_n568), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n577), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G299));
  NAND2_X1  g165(.A1(new_n510), .A2(G87), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n517), .A2(G49), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT77), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT78), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n591), .A2(new_n593), .A3(new_n595), .ZN(G288));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT79), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n515), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT80), .Z(new_n602));
  NAND2_X1  g177(.A1(new_n517), .A2(G48), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n503), .A2(new_n509), .ZN(new_n604));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n602), .A2(new_n606), .ZN(G305));
  XOR2_X1   g182(.A(KEYINPUT81), .B(G85), .Z(new_n608));
  NAND2_X1  g183(.A1(new_n510), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G60), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n515), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G47), .B2(new_n517), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n503), .A2(G92), .A3(new_n509), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n503), .A2(new_n509), .A3(new_n618), .A4(G92), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G79), .ZN(new_n623));
  OR3_X1    g198(.A1(new_n623), .A2(new_n496), .A3(KEYINPUT83), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT83), .B1(new_n623), .B2(new_n496), .ZN(new_n625));
  INV_X1    g200(.A(G66), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n515), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n627), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n619), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n615), .B1(new_n631), .B2(G868), .ZN(G284));
  OAI21_X1  g207(.A(new_n615), .B1(new_n631), .B2(G868), .ZN(G321));
  NAND2_X1  g208(.A1(G286), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n589), .B2(G868), .ZN(G297));
  OAI21_X1  g210(.A(new_n634), .B1(new_n589), .B2(G868), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n631), .B1(new_n637), .B2(G860), .ZN(G148));
  INV_X1    g213(.A(G868), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n551), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n631), .A2(new_n637), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT84), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n640), .B1(new_n642), .B2(new_n639), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n475), .A2(G135), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(new_n456), .B2(G111), .ZN(new_n648));
  INV_X1    g223(.A(G99), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(new_n456), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n473), .B2(G123), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n475), .A2(KEYINPUT85), .A3(G135), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(G2096), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n457), .A2(new_n467), .A3(new_n456), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT12), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n658), .ZN(G156));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT14), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1341), .B(G1348), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2443), .B(G2446), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G14), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2067), .B(G2678), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2072), .B(G2078), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT88), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n679), .B(KEYINPUT17), .Z(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(new_n677), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n677), .A3(new_n675), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n678), .A2(new_n679), .A3(new_n675), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT18), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G2096), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2100), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G227));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n691), .A2(new_n692), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n694), .A2(new_n696), .A3(new_n698), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n701), .B(new_n702), .C1(new_n700), .C2(new_n699), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT89), .B(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n703), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1991), .B(G1996), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1986), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(G229));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G16), .B2(G23), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n712), .A2(G16), .A3(G23), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n713), .B(new_n714), .C1(G288), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT33), .ZN(new_n717));
  INV_X1    g292(.A(G1976), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n715), .A2(G6), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n602), .A2(new_n606), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n715), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT32), .B(G1981), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G16), .A2(G22), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G166), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT93), .B(G1971), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n719), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n730));
  AOI21_X1  g305(.A(new_n711), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G16), .A2(G24), .ZN(new_n732));
  INV_X1    g307(.A(G290), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1986), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  AOI22_X1  g311(.A1(G119), .A2(new_n473), .B1(new_n475), .B2(G131), .ZN(new_n737));
  OR2_X1    g312(.A1(G95), .A2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n738), .B(G2104), .C1(G107), .C2(new_n456), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT90), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G25), .B(new_n741), .S(G29), .Z(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT35), .B(G1991), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n742), .B(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n730), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n719), .A2(new_n746), .A3(new_n724), .A4(new_n728), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n731), .A2(new_n736), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT95), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n715), .A2(KEYINPUT23), .A3(G20), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT23), .ZN(new_n753));
  INV_X1    g328(.A(G20), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G16), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n755), .C1(new_n589), .C2(new_n715), .ZN(new_n756));
  INV_X1    g331(.A(G1956), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n748), .A2(KEYINPUT95), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n748), .A2(KEYINPUT95), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n759), .A2(KEYINPUT36), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n456), .A2(G103), .A3(G2104), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT25), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n457), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n456), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n763), .B(new_n765), .C1(G139), .C2(new_n475), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT98), .B1(G29), .B2(G33), .ZN(new_n768));
  OR3_X1    g343(.A1(KEYINPUT98), .A2(G29), .A3(G33), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2072), .ZN(new_n771));
  INV_X1    g346(.A(G2084), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT24), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G34), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n471), .B2(G29), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G32), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n469), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(G2105), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n473), .A2(G129), .ZN(new_n782));
  NAND3_X1  g357(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT26), .Z(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT27), .B(G1996), .Z(new_n788));
  OAI221_X1 g363(.A(new_n771), .B1(new_n772), .B2(new_n778), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT99), .ZN(new_n790));
  INV_X1    g365(.A(G1966), .ZN(new_n791));
  NAND2_X1  g366(.A1(G168), .A2(G16), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G16), .B2(G21), .ZN(new_n793));
  INV_X1    g368(.A(G29), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G35), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G162), .B2(new_n794), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT29), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n790), .B1(new_n791), .B2(new_n793), .C1(G2090), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n794), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n794), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G2078), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n653), .A2(new_n794), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n793), .A2(new_n791), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT100), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT31), .B(G11), .Z(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n797), .A2(G2090), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT101), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT30), .B(G28), .Z(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(G29), .ZN(new_n810));
  NOR2_X1   g385(.A1(G5), .A2(G16), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G171), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1961), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n810), .B(new_n813), .C1(new_n772), .C2(new_n778), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n787), .A2(new_n788), .B1(G2078), .B2(new_n800), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n806), .A2(new_n808), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n798), .A2(new_n801), .A3(new_n802), .A4(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n751), .A2(new_n758), .A3(new_n761), .A4(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n794), .A2(G26), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n473), .A2(G128), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n475), .A2(G140), .ZN(new_n821));
  NOR2_X1   g396(.A1(G104), .A2(G2105), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(new_n456), .B2(G116), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n819), .B1(new_n824), .B2(G29), .ZN(new_n825));
  MUX2_X1   g400(.A(new_n819), .B(new_n825), .S(KEYINPUT28), .Z(new_n826));
  XOR2_X1   g401(.A(KEYINPUT96), .B(G2067), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n715), .A2(G4), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n631), .B2(new_n715), .ZN(new_n830));
  INV_X1    g405(.A(G1348), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n715), .A2(G19), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n552), .B2(new_n715), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(G1341), .Z(new_n835));
  NAND3_X1  g410(.A1(new_n828), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT97), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n818), .A2(new_n837), .ZN(G311));
  AND3_X1   g413(.A1(new_n759), .A2(KEYINPUT36), .A3(new_n760), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT36), .B1(new_n759), .B2(new_n760), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n837), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n841), .A2(new_n842), .A3(new_n758), .A4(new_n817), .ZN(G150));
  AND2_X1   g418(.A1(new_n510), .A2(G93), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n517), .A2(G55), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n574), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n630), .A2(new_n637), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT39), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n551), .A2(KEYINPUT102), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(new_n545), .C1(new_n549), .C2(new_n550), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n855), .A2(new_n848), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n848), .B1(new_n855), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n854), .B(new_n860), .Z(new_n861));
  OAI21_X1  g436(.A(new_n851), .B1(new_n861), .B2(G860), .ZN(G145));
  XNOR2_X1  g437(.A(new_n653), .B(new_n471), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  INV_X1    g439(.A(G126), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n486), .B1(new_n468), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n494), .B1(new_n866), .B2(G2105), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n489), .A2(KEYINPUT103), .A3(new_n492), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT103), .B1(new_n489), .B2(new_n492), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n864), .B(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n741), .B(new_n656), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n766), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n473), .A2(G130), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n475), .A2(G142), .ZN(new_n879));
  NOR2_X1   g454(.A1(G106), .A2(G2105), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(new_n456), .B2(G118), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n878), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n785), .B(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(new_n824), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n875), .A2(new_n884), .A3(new_n876), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g465(.A(new_n642), .B(new_n860), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n619), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT10), .B1(new_n617), .B2(new_n619), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n894), .A2(new_n577), .A3(new_n588), .A4(new_n628), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n589), .A2(new_n630), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT104), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n898));
  NAND3_X1  g473(.A1(G299), .A2(new_n631), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n899), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n895), .A2(new_n896), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n901), .B1(new_n905), .B2(new_n891), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  XNOR2_X1  g482(.A(G166), .B(G288), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(new_n721), .ZN(new_n909));
  XNOR2_X1  g484(.A(G288), .B(G303), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(G305), .ZN(new_n911));
  OAI21_X1  g486(.A(G290), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n721), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(G305), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n733), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n907), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n907), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(G868), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g497(.A(new_n921), .B1(G868), .B2(new_n848), .ZN(G331));
  XNOR2_X1  g498(.A(G286), .B(G171), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n858), .B2(new_n859), .ZN(new_n925));
  XNOR2_X1  g500(.A(G286), .B(G301), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n546), .A2(new_n548), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT72), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n856), .B1(new_n930), .B2(new_n545), .ZN(new_n931));
  INV_X1    g506(.A(new_n857), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n849), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n855), .A2(new_n848), .A3(new_n857), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n926), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n925), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n897), .A2(new_n899), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n900), .A2(new_n903), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n895), .A2(new_n896), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT41), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n925), .A2(new_n942), .A3(new_n935), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n938), .B(KEYINPUT105), .C1(new_n940), .C2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n936), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n939), .A4(new_n942), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n917), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n902), .A2(new_n904), .A3(new_n935), .A4(new_n925), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n938), .A2(new_n949), .A3(new_n916), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n950), .A2(new_n887), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT106), .ZN(new_n954));
  INV_X1    g529(.A(new_n951), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n916), .B1(new_n938), .B2(new_n949), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n948), .A2(new_n951), .A3(new_n958), .A4(new_n952), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n948), .A2(new_n951), .A3(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT107), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n962), .A2(new_n969), .A3(new_n966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(G397));
  XNOR2_X1  g546(.A(KEYINPUT108), .B(G1384), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n870), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n870), .A2(KEYINPUT109), .A3(new_n972), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(G40), .B(new_n461), .C1(new_n470), .C2(G2105), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n978), .A2(G1996), .A3(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(KEYINPUT46), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  INV_X1    g557(.A(G2067), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n824), .B(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n982), .B1(new_n785), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n980), .A2(KEYINPUT46), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n982), .A2(new_n735), .A3(new_n733), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT48), .ZN(new_n991));
  INV_X1    g566(.A(G1996), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n786), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n785), .A2(G1996), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n984), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n741), .A2(new_n743), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n737), .A2(new_n744), .A3(new_n740), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n982), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n991), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n997), .B(KEYINPUT126), .ZN(new_n1001));
  OAI22_X1  g576(.A1(new_n995), .A2(new_n1001), .B1(G2067), .B2(new_n824), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n982), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n989), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n1004), .B(KEYINPUT127), .Z(new_n1005));
  NOR3_X1   g580(.A1(new_n602), .A2(new_n606), .A3(G1981), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n606), .A2(KEYINPUT114), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n606), .A2(KEYINPUT114), .ZN(new_n1009));
  INV_X1    g584(.A(new_n601), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1007), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1011), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1006), .B1(new_n1017), .B2(G1981), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT49), .B1(new_n1018), .B2(KEYINPUT115), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT103), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n493), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n489), .A2(new_n492), .A3(KEYINPUT103), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1384), .B1(new_n1023), .B2(new_n867), .ZN(new_n1024));
  INV_X1    g599(.A(new_n979), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1016), .A2(new_n1019), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT112), .B1(G288), .B2(new_n718), .ZN(new_n1031));
  OR3_X1    g606(.A1(G288), .A2(KEYINPUT112), .A3(new_n718), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1030), .A2(G8), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  INV_X1    g611(.A(G288), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n1037), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1029), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n870), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(new_n1025), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n976), .B1(G164), .B2(G1384), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1971), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  INV_X1    g622(.A(G1384), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n870), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n1025), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT111), .B(G2090), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G303), .A2(G8), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT55), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(G8), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1040), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1029), .A2(new_n718), .A3(new_n1037), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1007), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n1028), .B2(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1058), .A2(new_n1029), .A3(new_n1039), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1051), .A2(G2084), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT45), .B1(new_n870), .B2(new_n1048), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n979), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT116), .B(new_n1025), .C1(new_n1024), .C2(KEYINPUT45), .ZN(new_n1068));
  OR3_X1    g643(.A1(G164), .A2(new_n976), .A3(G1384), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1064), .B1(new_n1070), .B2(new_n791), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1071), .A2(new_n1027), .A3(G286), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1054), .A2(G8), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(new_n1056), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1063), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT117), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1063), .A2(new_n1072), .A3(new_n1078), .A4(new_n1075), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OR2_X1    g655(.A1(G164), .A2(G1384), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1025), .B1(new_n1081), .B2(KEYINPUT50), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1024), .A2(new_n1047), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1082), .A2(new_n1052), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1056), .B1(new_n1085), .B2(new_n1027), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(new_n1058), .A3(new_n1029), .A4(new_n1039), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT63), .B1(new_n1088), .B2(new_n1072), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1062), .B1(new_n1080), .B2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT120), .B(KEYINPUT51), .Z(new_n1091));
  NOR2_X1   g666(.A1(new_n1071), .A2(new_n1027), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G286), .A2(G8), .ZN(new_n1093));
  XOR2_X1   g668(.A(new_n1093), .B(KEYINPUT121), .Z(new_n1094));
  OAI21_X1  g669(.A(new_n1091), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1093), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(KEYINPUT51), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1071), .B2(new_n1027), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(KEYINPUT122), .B(new_n1097), .C1(new_n1071), .C2(new_n1027), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1095), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1071), .A2(new_n1093), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1106), .A3(new_n1103), .ZN(new_n1107));
  INV_X1    g682(.A(G2078), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1041), .A2(new_n1043), .A3(new_n1025), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  INV_X1    g685(.A(G1961), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1109), .A2(new_n1110), .B1(new_n1051), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1108), .A2(KEYINPUT53), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1070), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G171), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1105), .A2(new_n1107), .A3(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT124), .B(G2078), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n978), .A2(KEYINPUT53), .A3(new_n1042), .A4(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(new_n1112), .A3(G301), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n562), .A2(new_n563), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n576), .B2(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1127), .A2(KEYINPUT118), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(KEYINPUT118), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n582), .A2(new_n568), .A3(new_n587), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1128), .B(new_n1129), .C1(new_n1125), .C2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n757), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1042), .A2(new_n1043), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n983), .A2(new_n1026), .B1(new_n1051), .B2(new_n831), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n630), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1135), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT58), .B(G1341), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1044), .A2(G1996), .B1(new_n1026), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n552), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(KEYINPUT119), .A3(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1137), .A2(new_n630), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT60), .B1(new_n1145), .B2(new_n1138), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1136), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1132), .A2(KEYINPUT61), .A3(new_n1134), .A4(new_n1131), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1137), .A2(new_n1151), .A3(new_n631), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1144), .A2(new_n1146), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1154));
  NOR2_X1   g729(.A1(new_n1142), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1139), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1120), .A2(new_n1112), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(G171), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1158), .B(KEYINPUT54), .C1(G171), .C2(new_n1114), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1124), .A2(new_n1156), .A3(new_n1104), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1117), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1090), .B1(new_n1161), .B2(new_n1088), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n982), .A2(G1986), .A3(G290), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n990), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT110), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n999), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1005), .B1(new_n1162), .B2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g742(.A1(new_n889), .A2(new_n673), .A3(new_n689), .ZN(new_n1169));
  INV_X1    g743(.A(G229), .ZN(new_n1170));
  NAND4_X1  g744(.A1(new_n1169), .A2(G319), .A3(new_n1170), .A4(new_n960), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


