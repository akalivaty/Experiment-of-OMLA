//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT0), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n188), .B(new_n190), .C1(new_n191), .C2(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n191), .A2(new_n192), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G101), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n198), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(G101), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n200), .A2(new_n203), .A3(new_n210), .A4(new_n204), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n188), .A2(new_n190), .ZN(new_n213));
  OAI211_X1 g027(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n189), .C2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G128), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT67), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n197), .A2(new_n218), .A3(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n199), .A2(G107), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n202), .A2(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n211), .A2(new_n223), .A3(KEYINPUT10), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n208), .A2(new_n212), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n192), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n197), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n218), .B1(G143), .B2(new_n187), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n213), .B(KEYINPUT78), .C1(new_n192), .C2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n231), .A3(new_n219), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n211), .A2(new_n223), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G131), .ZN(new_n237));
  INV_X1    g051(.A(G134), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT11), .B1(new_n238), .B2(G137), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT64), .B1(new_n241), .B2(G134), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n238), .A3(G137), .ZN(new_n246));
  AND4_X1   g060(.A1(new_n237), .A2(new_n243), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n244), .A2(new_n246), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n237), .B1(new_n248), .B2(new_n243), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n226), .A2(new_n236), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G110), .B(G140), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G227), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n252), .B(new_n254), .Z(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n211), .A2(new_n223), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n217), .A2(new_n258), .A3(new_n219), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n257), .B(new_n250), .C1(new_n234), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n234), .A2(new_n259), .ZN(new_n261));
  INV_X1    g075(.A(new_n250), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT12), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n251), .B(new_n256), .C1(new_n260), .C2(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n209), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n198), .A2(new_n207), .ZN(new_n266));
  AND4_X1   g080(.A1(new_n218), .A2(new_n188), .A3(new_n190), .A4(G128), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(G128), .A3(new_n214), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n267), .B1(new_n271), .B2(new_n213), .ZN(new_n272));
  OAI22_X1  g086(.A1(new_n265), .A2(new_n266), .B1(new_n272), .B2(new_n224), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT10), .B1(new_n232), .B2(new_n233), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n273), .A2(new_n262), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n250), .B1(new_n226), .B2(new_n236), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n255), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n264), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G469), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT79), .B1(new_n275), .B2(new_n255), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n262), .B1(new_n273), .B2(new_n274), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT79), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n251), .A2(new_n284), .A3(new_n256), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n251), .B1(new_n260), .B2(new_n263), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n255), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n288), .A3(G469), .ZN(new_n289));
  NAND2_X1  g103(.A1(G469), .A2(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n281), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G210), .B1(G237), .B2(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(KEYINPUT71), .A2(G125), .ZN(new_n294));
  NAND2_X1  g108(.A1(KEYINPUT71), .A2(G125), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n217), .A2(new_n219), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n295), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n193), .B(new_n297), .C1(new_n196), .C2(new_n197), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT82), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n213), .B1(new_n194), .B2(new_n195), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n301), .A2(KEYINPUT82), .A3(new_n193), .A4(new_n297), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n296), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G224), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(G953), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n303), .B(new_n306), .ZN(new_n307));
  OR2_X1    g121(.A1(KEYINPUT2), .A2(G113), .ZN(new_n308));
  AND3_X1   g122(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G116), .ZN(new_n313));
  INV_X1    g127(.A(G116), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G116), .B(G119), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n318), .B(new_n308), .C1(new_n310), .C2(new_n309), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n212), .A2(new_n320), .A3(new_n207), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT5), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n312), .A3(G116), .ZN(new_n323));
  OAI211_X1 g137(.A(G113), .B(new_n323), .C1(new_n316), .C2(new_n322), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n233), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G110), .B(G122), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n326), .A2(new_n328), .B1(new_n329), .B2(KEYINPUT6), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(KEYINPUT6), .ZN(new_n331));
  AOI211_X1 g145(.A(new_n327), .B(new_n331), .C1(new_n321), .C2(new_n325), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n321), .A2(new_n325), .A3(new_n327), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT81), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n321), .A2(new_n336), .A3(new_n325), .A4(new_n327), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(KEYINPUT6), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n307), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(new_n337), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n306), .A2(KEYINPUT7), .ZN(new_n341));
  AND4_X1   g155(.A1(new_n296), .A2(new_n300), .A3(new_n302), .A4(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(new_n327), .B(KEYINPUT8), .Z(new_n343));
  AND3_X1   g157(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT5), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n323), .A2(G113), .ZN(new_n345));
  OAI22_X1  g159(.A1(new_n344), .A2(new_n345), .B1(new_n311), .B2(new_n316), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n258), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n343), .B1(new_n325), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n341), .B1(new_n296), .B2(new_n298), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n342), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n340), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n280), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n293), .B1(new_n339), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n307), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n335), .A2(KEYINPUT6), .A3(new_n337), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n346), .A2(new_n258), .ZN(new_n356));
  INV_X1    g170(.A(new_n209), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n357), .A2(new_n206), .B1(new_n319), .B2(new_n317), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n356), .B1(new_n358), .B2(new_n212), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n331), .B1(new_n359), .B2(new_n327), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n326), .A2(new_n329), .A3(KEYINPUT6), .A4(new_n328), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n354), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(G902), .B1(new_n340), .B2(new_n350), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n292), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n353), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G214), .B1(G237), .B2(G902), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT9), .B(G234), .ZN(new_n368));
  OAI21_X1  g182(.A(G221), .B1(new_n368), .B2(G902), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT77), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n291), .A2(new_n366), .A3(new_n367), .A4(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(G116), .B(G122), .Z(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G107), .ZN(new_n374));
  XNOR2_X1  g188(.A(G116), .B(G122), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n202), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT13), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n189), .A3(G128), .ZN(new_n379));
  XOR2_X1   g193(.A(G128), .B(G143), .Z(new_n380));
  OAI211_X1 g194(.A(G134), .B(new_n379), .C1(new_n380), .C2(new_n378), .ZN(new_n381));
  XNOR2_X1  g195(.A(G128), .B(G143), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n238), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(KEYINPUT86), .A3(new_n238), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n377), .A2(new_n381), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n380), .A2(G134), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n383), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n314), .A2(KEYINPUT14), .A3(G122), .ZN(new_n390));
  OAI211_X1 g204(.A(G107), .B(new_n390), .C1(new_n373), .C2(KEYINPUT14), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n391), .A3(new_n376), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G217), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n368), .A2(new_n394), .A3(G953), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n387), .A2(new_n392), .A3(new_n395), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n280), .ZN(new_n400));
  INV_X1    g214(.A(G478), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(KEYINPUT15), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n400), .B(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n253), .A2(G952), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(G234), .B2(G237), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT21), .B(G898), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(G234), .A2(G237), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(G902), .A3(G953), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n406), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT87), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n403), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n199), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n294), .A2(G140), .A3(new_n295), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT70), .ZN(new_n418));
  INV_X1    g232(.A(G140), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(KEYINPUT70), .A2(G140), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(G125), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n417), .A2(new_n422), .A3(KEYINPUT83), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(G146), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G125), .B(G140), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n187), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(new_n237), .ZN(new_n432));
  NOR2_X1   g246(.A1(G237), .A2(G953), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(G143), .A3(G214), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(G143), .B1(new_n433), .B2(G214), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n253), .A3(G214), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n189), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n440), .B(new_n434), .C1(new_n431), .C2(new_n237), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n430), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT84), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n430), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G131), .B1(new_n435), .B2(new_n436), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(new_n237), .A3(new_n434), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(KEYINPUT17), .B(G131), .C1(new_n435), .C2(new_n436), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n417), .A2(new_n422), .A3(KEYINPUT16), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT16), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n297), .A2(new_n456), .A3(new_n419), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n455), .A2(KEYINPUT72), .A3(G146), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n457), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n187), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(G146), .A3(new_n457), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT72), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n454), .A2(new_n458), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n416), .B1(new_n448), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n446), .B1(new_n430), .B2(new_n443), .ZN(new_n466));
  AOI211_X1 g280(.A(KEYINPUT84), .B(new_n442), .C1(new_n427), .C2(new_n429), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n464), .B(new_n416), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n280), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G475), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT20), .ZN(new_n472));
  INV_X1    g286(.A(new_n416), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n425), .A2(KEYINPUT19), .A3(new_n426), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT19), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n428), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(new_n187), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT73), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n461), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n455), .A2(KEYINPUT73), .A3(G146), .A4(new_n457), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n449), .A2(new_n451), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n474), .A2(KEYINPUT85), .A3(new_n187), .A4(new_n476), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n466), .A2(new_n467), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n473), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n468), .ZN(new_n490));
  NOR2_X1   g304(.A1(G475), .A2(G902), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n472), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n416), .B1(new_n448), .B2(new_n486), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n472), .B(new_n491), .C1(new_n493), .C2(new_n469), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n414), .B(new_n471), .C1(new_n492), .C2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n372), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n198), .B1(new_n247), .B2(new_n249), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n248), .A2(new_n237), .A3(new_n243), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT65), .B1(new_n238), .B2(G137), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n241), .A3(G134), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n238), .A2(G137), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n504), .A2(new_n505), .A3(G131), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n504), .B2(G131), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n499), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n498), .B1(new_n508), .B2(new_n272), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n320), .B1(new_n509), .B2(KEYINPUT69), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n220), .B(new_n499), .C1(new_n506), .C2(new_n507), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT69), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(new_n498), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n433), .A2(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n509), .A2(new_n320), .ZN(new_n521));
  INV_X1    g335(.A(new_n320), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n511), .A2(new_n498), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n515), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n516), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n527));
  INV_X1    g341(.A(new_n520), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n511), .B2(new_n498), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n498), .B(new_n529), .C1(new_n508), .C2(new_n272), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n522), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n523), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n528), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n526), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n280), .B1(new_n526), .B2(new_n527), .ZN(new_n537));
  OAI21_X1  g351(.A(G472), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n532), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n320), .B1(new_n539), .B2(new_n530), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n520), .A3(new_n523), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT31), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n540), .A2(new_n543), .A3(new_n520), .A4(new_n523), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT28), .B1(new_n510), .B2(new_n513), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n528), .B1(new_n545), .B2(new_n524), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n547), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n538), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n192), .A2(G119), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT23), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n556));
  INV_X1    g370(.A(G110), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n312), .A2(G128), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n553), .A2(new_n558), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT24), .B(G110), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n559), .A2(new_n562), .B1(new_n187), .B2(new_n428), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n481), .A2(new_n482), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT74), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT74), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n481), .A2(new_n566), .A3(new_n482), .A4(new_n563), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n463), .A2(new_n458), .A3(new_n460), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n560), .A2(new_n561), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(G110), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(KEYINPUT75), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT22), .B(G137), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n575), .B(new_n576), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n565), .A2(new_n567), .B1(new_n569), .B2(new_n572), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT75), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n573), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n577), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n280), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT25), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n577), .B1(new_n580), .B2(KEYINPUT75), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n584), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n591), .B2(new_n585), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT25), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n394), .B1(G234), .B2(new_n280), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n588), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n585), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n595), .A2(G902), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT76), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT76), .ZN(new_n600));
  INV_X1    g414(.A(new_n598), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n600), .B(new_n601), .C1(new_n591), .C2(new_n585), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n497), .A2(new_n552), .A3(new_n596), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n547), .A2(new_n280), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n606), .A2(G472), .B1(new_n547), .B2(new_n549), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n291), .A2(new_n371), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n596), .A2(new_n607), .A3(new_n603), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n363), .A2(KEYINPUT88), .A3(new_n292), .A4(new_n364), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n367), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n612), .B1(KEYINPUT88), .B2(new_n366), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n491), .B1(new_n493), .B2(new_n469), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT20), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n615), .A2(new_n494), .B1(G475), .B2(new_n470), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  INV_X1    g431(.A(new_n398), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n395), .B1(new_n387), .B2(new_n392), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT89), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n399), .A2(KEYINPUT89), .A3(new_n617), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n619), .A2(new_n617), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT90), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n398), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n387), .A2(new_n392), .A3(KEYINPUT90), .A4(new_n395), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n625), .A2(KEYINPUT91), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT91), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n401), .A2(G902), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n624), .A2(new_n629), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n400), .A2(new_n401), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR4_X1   g450(.A1(new_n613), .A2(new_n616), .A3(new_n413), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n610), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NAND2_X1  g455(.A1(new_n616), .A2(new_n403), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n642), .A2(new_n613), .A3(new_n413), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n610), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n578), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n583), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n598), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n595), .B1(new_n592), .B2(new_n593), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT25), .B(G902), .C1(new_n591), .C2(new_n585), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n497), .A2(new_n607), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  OR2_X1    g469(.A1(new_n410), .A2(G900), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n406), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n642), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n613), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n552), .A2(new_n652), .A3(new_n608), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n192), .ZN(G30));
  XNOR2_X1  g478(.A(new_n657), .B(KEYINPUT39), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n608), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT40), .Z(new_n667));
  INV_X1    g481(.A(new_n652), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n366), .B(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n471), .B1(new_n492), .B2(new_n495), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n403), .ZN(new_n672));
  INV_X1    g486(.A(new_n367), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n667), .A2(new_n668), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n547), .A2(new_n549), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT32), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT94), .Z(new_n681));
  INV_X1    g495(.A(new_n541), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n280), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT95), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n675), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  AOI22_X1  g503(.A1(new_n679), .A2(new_n538), .B1(new_n596), .B2(new_n649), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT96), .ZN(new_n691));
  INV_X1    g505(.A(new_n636), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n671), .A2(new_n692), .A3(new_n657), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n613), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n690), .A2(new_n691), .A3(new_n608), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n615), .A2(new_n494), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n636), .B1(new_n696), .B2(new_n471), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n366), .A2(KEYINPUT88), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n612), .A4(new_n657), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT96), .B1(new_n662), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT97), .B(G146), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G48));
  AOI21_X1  g517(.A(new_n256), .B1(new_n283), .B2(new_n251), .ZN(new_n704));
  INV_X1    g518(.A(new_n263), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n261), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n275), .A2(new_n255), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(G469), .B1(new_n709), .B2(G902), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT98), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n281), .ZN(new_n712));
  OAI211_X1 g526(.A(KEYINPUT98), .B(G469), .C1(new_n709), .C2(G902), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT99), .B1(new_n714), .B2(new_n369), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT99), .ZN(new_n716));
  INV_X1    g530(.A(new_n369), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n716), .B(new_n717), .C1(new_n712), .C2(new_n713), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n545), .A2(new_n524), .A3(new_n528), .ZN(new_n720));
  AOI21_X1  g534(.A(G902), .B1(new_n720), .B2(KEYINPUT29), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n526), .A2(new_n527), .A3(new_n535), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n677), .A2(new_n678), .B1(G472), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n597), .A2(new_n598), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n600), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n597), .A2(KEYINPUT76), .A3(new_n598), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n726), .B(new_n727), .C1(new_n650), .C2(new_n651), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n719), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n637), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n643), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  AND2_X1   g549(.A1(new_n616), .A2(new_n414), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n719), .A2(new_n690), .A3(new_n736), .A4(new_n660), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  INV_X1    g552(.A(new_n607), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT100), .B1(new_n728), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n672), .A2(new_n613), .A3(new_n413), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT100), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n596), .A2(new_n607), .A3(new_n603), .A4(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n740), .A2(new_n719), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  NOR3_X1   g559(.A1(new_n715), .A2(new_n718), .A3(new_n613), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT102), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n697), .B2(new_n657), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n616), .A2(new_n636), .A3(KEYINPUT102), .A4(new_n658), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n652), .A2(new_n607), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT101), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT101), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n652), .A2(new_n753), .A3(new_n607), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n746), .A2(new_n750), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  INV_X1    g570(.A(new_n728), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n291), .A2(new_n369), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n353), .A2(new_n365), .A3(new_n367), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT103), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n353), .A2(new_n365), .A3(new_n367), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT103), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n291), .A4(new_n369), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n757), .A2(new_n764), .A3(new_n552), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT42), .B1(new_n765), .B2(new_n750), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n693), .A2(KEYINPUT102), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n697), .A2(new_n747), .A3(new_n657), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n767), .A3(KEYINPUT42), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n550), .B2(new_n551), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n677), .A2(KEYINPUT104), .A3(new_n678), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n538), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n757), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT105), .B1(new_n766), .B2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n769), .A2(new_n774), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n729), .A2(new_n764), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n767), .A2(new_n768), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT105), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n777), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n776), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n237), .ZN(G33));
  NAND4_X1  g599(.A1(new_n757), .A2(new_n764), .A3(new_n552), .A4(new_n659), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  NAND2_X1  g601(.A1(new_n616), .A2(new_n692), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n739), .A3(new_n652), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT45), .B1(new_n286), .B2(new_n288), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n279), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT45), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n290), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(KEYINPUT106), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(KEYINPUT106), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n290), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n799), .A2(new_n281), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n804), .A2(new_n369), .A3(new_n665), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n791), .A2(new_n792), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n793), .A2(new_n761), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  NAND2_X1  g622(.A1(new_n804), .A2(new_n369), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n804), .B(new_n369), .C1(KEYINPUT107), .C2(new_n813), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n757), .A2(new_n552), .A3(new_n693), .A4(new_n759), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  XOR2_X1   g631(.A(new_n714), .B(KEYINPUT49), .Z(new_n818));
  NAND3_X1  g632(.A1(new_n670), .A2(new_n367), .A3(new_n371), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n818), .A2(new_n788), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n757), .A3(new_n687), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n812), .A2(new_n814), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n714), .A2(new_n370), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n790), .A2(new_n405), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n740), .A3(new_n743), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n759), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n823), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n719), .A2(new_n673), .A3(new_n670), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n827), .A2(new_n832), .A3(new_n740), .A4(new_n743), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n687), .A2(new_n757), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n719), .A2(new_n761), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n406), .B1(new_n837), .B2(KEYINPUT113), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n671), .A2(new_n692), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n836), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n752), .A2(new_n754), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n838), .A2(new_n839), .A3(new_n842), .A4(new_n790), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n831), .A2(new_n835), .A3(new_n844), .ZN(new_n845));
  OR3_X1    g659(.A1(new_n826), .A2(new_n823), .A3(new_n830), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT51), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  INV_X1    g662(.A(new_n826), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n829), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n835), .A2(new_n844), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n774), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n838), .A2(new_n839), .A3(new_n852), .A4(new_n790), .ZN(new_n853));
  XOR2_X1   g667(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n854));
  XOR2_X1   g668(.A(new_n853), .B(new_n854), .Z(new_n855));
  AND4_X1   g669(.A1(new_n697), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n714), .A2(new_n369), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n716), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n714), .A2(KEYINPUT99), .A3(new_n369), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n660), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n828), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n404), .B(KEYINPUT114), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n855), .A2(new_n856), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n851), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n822), .B1(new_n847), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n831), .A2(new_n835), .A3(new_n846), .A4(new_n844), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n848), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(KEYINPUT116), .A3(new_n851), .A4(new_n863), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT108), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n729), .B(new_n719), .C1(new_n637), .C2(new_n643), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n871), .A2(new_n744), .A3(new_n737), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n750), .A2(new_n752), .A3(new_n754), .A4(new_n764), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n671), .A2(new_n759), .A3(new_n403), .A4(new_n658), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n552), .A3(new_n608), .A4(new_n652), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n786), .A2(new_n875), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n413), .B(new_n673), .C1(new_n353), .C2(new_n365), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n696), .A2(new_n471), .A3(new_n403), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n877), .B1(new_n878), .B2(new_n697), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n604), .B(new_n653), .C1(new_n609), .C2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n872), .A2(new_n873), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n870), .B1(new_n784), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n663), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n672), .A2(new_n613), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n758), .A2(new_n658), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n685), .A2(new_n885), .A3(new_n668), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n701), .A2(new_n884), .A3(new_n755), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n786), .A2(new_n875), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n604), .A2(new_n653), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n879), .A2(new_n609), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n891), .A2(new_n894), .A3(new_n873), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n871), .A2(new_n744), .A3(new_n737), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(KEYINPUT108), .A3(new_n776), .A4(new_n783), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n883), .A2(new_n890), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n895), .A2(new_n900), .ZN(new_n903));
  XOR2_X1   g717(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n888), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n860), .A2(new_n780), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n663), .B1(new_n842), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(new_n889), .A3(new_n701), .A4(new_n887), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n903), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n777), .A2(new_n781), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n872), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT111), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n911), .A2(new_n872), .A3(KEYINPUT111), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n901), .A2(new_n902), .A3(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n899), .A2(KEYINPUT110), .A3(new_n900), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT110), .ZN(new_n920));
  AND4_X1   g734(.A1(new_n883), .A2(new_n898), .A3(new_n909), .A4(new_n906), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(KEYINPUT53), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n899), .A2(new_n900), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n918), .B1(new_n924), .B2(new_n902), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n869), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(G952), .A2(G953), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT117), .Z(new_n928));
  OAI21_X1  g742(.A(new_n821), .B1(new_n926), .B2(new_n928), .ZN(G75));
  AOI21_X1  g743(.A(new_n280), .B1(new_n901), .B2(new_n917), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(G210), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n355), .A2(new_n362), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n307), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n363), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n933), .A2(new_n937), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n253), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  INV_X1    g755(.A(KEYINPUT118), .ZN(new_n942));
  INV_X1    g756(.A(new_n940), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n901), .A2(new_n917), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT54), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n918), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n290), .B(KEYINPUT57), .Z(new_n947));
  AOI21_X1  g761(.A(new_n709), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n280), .B(new_n797), .C1(new_n901), .C2(new_n917), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n942), .B(new_n943), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  AOI221_X4 g764(.A(KEYINPUT54), .B1(new_n916), .B2(new_n910), .C1(new_n899), .C2(new_n900), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n902), .B1(new_n901), .B2(new_n917), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n949), .B1(new_n953), .B2(new_n278), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT118), .B1(new_n954), .B2(new_n940), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n950), .A2(new_n955), .ZN(G54));
  NAND3_X1  g770(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n957));
  INV_X1    g771(.A(new_n490), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n940), .ZN(G60));
  INV_X1    g775(.A(new_n946), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n624), .A2(new_n629), .A3(new_n632), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT119), .ZN(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n401), .A2(new_n280), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n965), .B(new_n966), .Z(new_n967));
  OR2_X1    g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n943), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n967), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n925), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n971), .B2(new_n964), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT60), .Z(new_n974));
  AOI21_X1  g788(.A(new_n597), .B1(new_n944), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n975), .A2(new_n940), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT121), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT61), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n944), .A2(new_n648), .A3(new_n974), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n976), .B(new_n979), .C1(new_n977), .C2(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n407), .B2(new_n304), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n896), .A2(new_n880), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n934), .B1(G898), .B2(new_n253), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT122), .Z(new_n988));
  XNOR2_X1  g802(.A(new_n986), .B(new_n988), .ZN(G69));
  NAND3_X1  g803(.A1(new_n701), .A2(new_n884), .A3(new_n755), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n688), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n666), .A2(new_n759), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n729), .B(new_n996), .C1(new_n697), .C2(new_n878), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n807), .A2(new_n816), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n994), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n253), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n531), .A2(new_n532), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n474), .A2(new_n476), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1001), .B(new_n1002), .Z(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT123), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n253), .A2(G900), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n774), .A2(new_n613), .A3(new_n672), .ZN(new_n1008));
  AOI22_X1  g822(.A1(new_n805), .A2(new_n1008), .B1(new_n659), .B2(new_n765), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n807), .A2(new_n816), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n784), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n1010), .A2(new_n1011), .A3(new_n992), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1007), .B1(new_n1012), .B2(G953), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT125), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n1003), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1005), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(G72));
  NAND2_X1  g834(.A1(new_n1012), .A2(new_n985), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT126), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n533), .A2(new_n534), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n528), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1026), .A2(new_n528), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1029), .A2(new_n1023), .A3(new_n1027), .ZN(new_n1030));
  OAI221_X1 g844(.A(new_n943), .B1(new_n1025), .B2(new_n1027), .C1(new_n924), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(new_n985), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1024), .B1(new_n999), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n1028), .ZN(new_n1034));
  OR2_X1    g848(.A1(new_n1034), .A2(KEYINPUT127), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(KEYINPUT127), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1031), .B1(new_n1035), .B2(new_n1036), .ZN(G57));
endmodule


