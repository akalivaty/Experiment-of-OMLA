

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U556 ( .A(G543), .B(KEYINPUT0), .Z(n523) );
  NAND2_X1 U557 ( .A1(G29), .A2(n979), .ZN(n524) );
  AND2_X1 U558 ( .A1(n789), .A2(n788), .ZN(n525) );
  AND2_X1 U559 ( .A1(n790), .A2(n525), .ZN(n526) );
  NOR2_X1 U560 ( .A1(n991), .A2(n714), .ZN(n717) );
  INV_X1 U561 ( .A(KEYINPUT98), .ZN(n715) );
  AND2_X1 U562 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U563 ( .A1(n738), .A2(n737), .ZN(n739) );
  INV_X1 U564 ( .A(KEYINPUT104), .ZN(n772) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n807) );
  NAND2_X1 U566 ( .A1(n588), .A2(n587), .ZN(n991) );
  XNOR2_X1 U567 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n528) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U569 ( .A(n528), .B(n527), .ZN(n611) );
  NAND2_X1 U570 ( .A1(G138), .A2(n611), .ZN(n529) );
  XNOR2_X1 U571 ( .A(n529), .B(KEYINPUT88), .ZN(n533) );
  INV_X1 U572 ( .A(G2105), .ZN(n530) );
  AND2_X1 U573 ( .A1(G2104), .A2(n530), .ZN(n531) );
  XNOR2_X1 U574 ( .A(n531), .B(KEYINPUT64), .ZN(n613) );
  NAND2_X1 U575 ( .A1(G102), .A2(n613), .ZN(n532) );
  NAND2_X1 U576 ( .A1(n533), .A2(n532), .ZN(n540) );
  INV_X1 U577 ( .A(KEYINPUT87), .ZN(n538) );
  NOR2_X1 U578 ( .A1(G2104), .A2(n530), .ZN(n556) );
  NAND2_X1 U579 ( .A1(n556), .A2(G126), .ZN(n534) );
  XNOR2_X1 U580 ( .A(n534), .B(KEYINPUT86), .ZN(n536) );
  AND2_X1 U581 ( .A1(G2104), .A2(G2105), .ZN(n892) );
  NAND2_X1 U582 ( .A1(G114), .A2(n892), .ZN(n535) );
  NAND2_X1 U583 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U584 ( .A(n538), .B(n537), .ZN(n539) );
  NOR2_X1 U585 ( .A1(n540), .A2(n539), .ZN(G164) );
  XNOR2_X1 U586 ( .A(KEYINPUT66), .B(n523), .ZN(n660) );
  NOR2_X2 U587 ( .A1(G651), .A2(n660), .ZN(n658) );
  NAND2_X1 U588 ( .A1(n658), .A2(G51), .ZN(n541) );
  XOR2_X1 U589 ( .A(KEYINPUT71), .B(n541), .Z(n544) );
  INV_X1 U590 ( .A(G651), .ZN(n547) );
  NOR2_X1 U591 ( .A1(G543), .A2(n547), .ZN(n542) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n542), .Z(n664) );
  NAND2_X1 U593 ( .A1(n664), .A2(G63), .ZN(n543) );
  NAND2_X1 U594 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U595 ( .A(KEYINPUT6), .B(n545), .ZN(n553) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U597 ( .A1(n649), .A2(G89), .ZN(n546) );
  XNOR2_X1 U598 ( .A(n546), .B(KEYINPUT4), .ZN(n549) );
  NOR2_X2 U599 ( .A1(n547), .A2(n660), .ZN(n652) );
  NAND2_X1 U600 ( .A1(G76), .A2(n652), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U602 ( .A(KEYINPUT5), .B(n550), .Z(n551) );
  XNOR2_X1 U603 ( .A(KEYINPUT70), .B(n551), .ZN(n552) );
  NOR2_X1 U604 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U605 ( .A(KEYINPUT7), .B(n554), .Z(G168) );
  NAND2_X1 U606 ( .A1(n613), .A2(G101), .ZN(n555) );
  XNOR2_X1 U607 ( .A(KEYINPUT23), .B(n555), .ZN(n562) );
  NAND2_X1 U608 ( .A1(n611), .A2(G137), .ZN(n560) );
  BUF_X1 U609 ( .A(n556), .Z(n890) );
  NAND2_X1 U610 ( .A1(G125), .A2(n890), .ZN(n558) );
  NAND2_X1 U611 ( .A1(G113), .A2(n892), .ZN(n557) );
  AND2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X2 U614 ( .A1(n562), .A2(n561), .ZN(G160) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U616 ( .A(G108), .ZN(G238) );
  INV_X1 U617 ( .A(G120), .ZN(G236) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  NAND2_X1 U621 ( .A1(G65), .A2(n664), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G53), .A2(n658), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U624 ( .A1(G78), .A2(n652), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G91), .A2(n649), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n731) );
  INV_X1 U628 ( .A(n731), .ZN(G299) );
  NAND2_X1 U629 ( .A1(G64), .A2(n664), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G52), .A2(n658), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n575) );
  NAND2_X1 U632 ( .A1(G77), .A2(n652), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G90), .A2(n649), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U636 ( .A1(n575), .A2(n574), .ZN(G171) );
  INV_X1 U637 ( .A(G171), .ZN(G301) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U639 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U640 ( .A(G567), .ZN(n691) );
  NOR2_X1 U641 ( .A1(n691), .A2(G223), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT11), .ZN(G234) );
  XOR2_X1 U643 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n579) );
  NAND2_X1 U644 ( .A1(G56), .A2(n664), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n586) );
  XNOR2_X1 U646 ( .A(KEYINPUT69), .B(KEYINPUT13), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n649), .A2(G81), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT12), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G68), .A2(n652), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U651 ( .A(n584), .B(n583), .ZN(n585) );
  NOR2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n658), .A2(G43), .ZN(n587) );
  INV_X1 U654 ( .A(G860), .ZN(n600) );
  OR2_X1 U655 ( .A1(n991), .A2(n600), .ZN(G153) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U657 ( .A1(G66), .A2(n664), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G92), .A2(n649), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U660 ( .A1(G79), .A2(n652), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G54), .A2(n658), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U664 ( .A(KEYINPUT15), .B(n595), .Z(n988) );
  OR2_X1 U665 ( .A1(n988), .A2(G868), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(G284) );
  XOR2_X1 U667 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n599) );
  INV_X1 U669 ( .A(G868), .ZN(n676) );
  NOR2_X1 U670 ( .A1(G286), .A2(n676), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n601), .A2(n988), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U675 ( .A1(n988), .A2(G868), .ZN(n603) );
  XNOR2_X1 U676 ( .A(KEYINPUT72), .B(n603), .ZN(n604) );
  NOR2_X1 U677 ( .A1(G559), .A2(n604), .ZN(n606) );
  NOR2_X1 U678 ( .A1(G868), .A2(n991), .ZN(n605) );
  NOR2_X1 U679 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G123), .A2(n890), .ZN(n607) );
  XOR2_X1 U681 ( .A(KEYINPUT18), .B(n607), .Z(n608) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT73), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G111), .A2(n892), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n618) );
  INV_X1 U685 ( .A(n611), .ZN(n612) );
  INV_X1 U686 ( .A(n612), .ZN(n896) );
  NAND2_X1 U687 ( .A1(G135), .A2(n896), .ZN(n616) );
  INV_X1 U688 ( .A(n613), .ZN(n614) );
  INV_X1 U689 ( .A(n614), .ZN(n899) );
  NAND2_X1 U690 ( .A1(G99), .A2(n899), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n960) );
  XNOR2_X1 U693 ( .A(n960), .B(G2096), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT74), .ZN(n621) );
  INV_X1 U695 ( .A(G2100), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(G156) );
  XNOR2_X1 U697 ( .A(n991), .B(KEYINPUT75), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n988), .A2(G559), .ZN(n622) );
  XOR2_X1 U699 ( .A(n623), .B(n622), .Z(n673) );
  NOR2_X1 U700 ( .A1(n673), .A2(G860), .ZN(n632) );
  NAND2_X1 U701 ( .A1(G67), .A2(n664), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G55), .A2(n658), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n626), .B(KEYINPUT77), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G93), .A2(n649), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n652), .A2(G80), .ZN(n629) );
  XOR2_X1 U708 ( .A(KEYINPUT76), .B(n629), .Z(n630) );
  NOR2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n675) );
  XNOR2_X1 U710 ( .A(n632), .B(n675), .ZN(G145) );
  NAND2_X1 U711 ( .A1(G73), .A2(n652), .ZN(n633) );
  XNOR2_X1 U712 ( .A(n633), .B(KEYINPUT2), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G61), .A2(n664), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G86), .A2(n649), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G48), .A2(n658), .ZN(n636) );
  XNOR2_X1 U717 ( .A(KEYINPUT79), .B(n636), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U720 ( .A1(G75), .A2(n652), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G88), .A2(n649), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n647) );
  NAND2_X1 U723 ( .A1(G62), .A2(n664), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G50), .A2(n658), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U726 ( .A(KEYINPUT80), .B(n645), .ZN(n646) );
  NOR2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U728 ( .A(n648), .B(KEYINPUT81), .ZN(G303) );
  INV_X1 U729 ( .A(G303), .ZN(G166) );
  NAND2_X1 U730 ( .A1(G85), .A2(n649), .ZN(n651) );
  NAND2_X1 U731 ( .A1(G47), .A2(n658), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U733 ( .A1(G72), .A2(n652), .ZN(n653) );
  XNOR2_X1 U734 ( .A(KEYINPUT67), .B(n653), .ZN(n654) );
  NOR2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U736 ( .A1(n664), .A2(G60), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n657), .A2(n656), .ZN(G290) );
  NAND2_X1 U738 ( .A1(G49), .A2(n658), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n659), .B(KEYINPUT78), .ZN(n666) );
  NAND2_X1 U740 ( .A1(G651), .A2(G74), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G87), .A2(n660), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U743 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n666), .A2(n665), .ZN(G288) );
  XOR2_X1 U745 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n667) );
  XNOR2_X1 U746 ( .A(G305), .B(n667), .ZN(n668) );
  XOR2_X1 U747 ( .A(n668), .B(n675), .Z(n670) );
  XNOR2_X1 U748 ( .A(G166), .B(n731), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n671), .B(G290), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n672), .B(G288), .ZN(n866) );
  XOR2_X1 U752 ( .A(n673), .B(n866), .Z(n674) );
  NAND2_X1 U753 ( .A1(n674), .A2(G868), .ZN(n678) );
  NAND2_X1 U754 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U756 ( .A(KEYINPUT83), .B(n679), .ZN(G295) );
  XOR2_X1 U757 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n681) );
  NAND2_X1 U758 ( .A1(G2084), .A2(G2078), .ZN(n680) );
  XNOR2_X1 U759 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U762 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U766 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U767 ( .A1(G96), .A2(n687), .ZN(n842) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n842), .ZN(n688) );
  XNOR2_X1 U769 ( .A(n688), .B(KEYINPUT85), .ZN(n693) );
  NOR2_X1 U770 ( .A1(G236), .A2(G238), .ZN(n689) );
  NAND2_X1 U771 ( .A1(G69), .A2(n689), .ZN(n690) );
  NOR2_X1 U772 ( .A1(G237), .A2(n690), .ZN(n844) );
  NOR2_X1 U773 ( .A1(n691), .A2(n844), .ZN(n692) );
  NOR2_X1 U774 ( .A1(n693), .A2(n692), .ZN(G319) );
  INV_X1 U775 ( .A(G319), .ZN(n695) );
  NAND2_X1 U776 ( .A1(G483), .A2(G661), .ZN(n694) );
  NOR2_X1 U777 ( .A1(n695), .A2(n694), .ZN(n841) );
  NAND2_X1 U778 ( .A1(n841), .A2(G36), .ZN(G176) );
  XNOR2_X1 U779 ( .A(G1981), .B(G305), .ZN(n997) );
  NAND2_X1 U780 ( .A1(G160), .A2(G40), .ZN(n806) );
  INV_X1 U781 ( .A(n806), .ZN(n696) );
  NAND2_X2 U782 ( .A1(n807), .A2(n696), .ZN(n750) );
  AND2_X1 U783 ( .A1(n750), .A2(G8), .ZN(n697) );
  XNOR2_X1 U784 ( .A(KEYINPUT93), .B(n697), .ZN(n787) );
  NOR2_X1 U785 ( .A1(G1966), .A2(n787), .ZN(n743) );
  OR2_X1 U786 ( .A1(G2084), .A2(n750), .ZN(n698) );
  XNOR2_X1 U787 ( .A(KEYINPUT96), .B(n698), .ZN(n744) );
  NAND2_X1 U788 ( .A1(G8), .A2(n744), .ZN(n699) );
  NOR2_X1 U789 ( .A1(n743), .A2(n699), .ZN(n700) );
  XNOR2_X1 U790 ( .A(n700), .B(KEYINPUT30), .ZN(n702) );
  INV_X1 U791 ( .A(G168), .ZN(n701) );
  XOR2_X1 U792 ( .A(KEYINPUT100), .B(n703), .Z(n708) );
  NAND2_X1 U793 ( .A1(G1961), .A2(n750), .ZN(n706) );
  INV_X1 U794 ( .A(n750), .ZN(n724) );
  XNOR2_X1 U795 ( .A(G2078), .B(KEYINPUT25), .ZN(n704) );
  XNOR2_X1 U796 ( .A(n704), .B(KEYINPUT97), .ZN(n939) );
  NAND2_X1 U797 ( .A1(n724), .A2(n939), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n736) );
  NAND2_X1 U799 ( .A1(G301), .A2(n736), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U801 ( .A(n709), .B(KEYINPUT31), .ZN(n741) );
  INV_X1 U802 ( .A(G1996), .ZN(n934) );
  NOR2_X1 U803 ( .A1(n750), .A2(n934), .ZN(n711) );
  INV_X1 U804 ( .A(KEYINPUT26), .ZN(n710) );
  XNOR2_X1 U805 ( .A(n711), .B(n710), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n750), .A2(G1341), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U808 ( .A1(n717), .A2(n988), .ZN(n716) );
  XNOR2_X1 U809 ( .A(n716), .B(n715), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n717), .A2(n988), .ZN(n721) );
  NOR2_X1 U811 ( .A1(n724), .A2(G1348), .ZN(n719) );
  NOR2_X1 U812 ( .A1(G2067), .A2(n750), .ZN(n718) );
  NOR2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n729) );
  NAND2_X1 U816 ( .A1(n724), .A2(G2072), .ZN(n725) );
  XNOR2_X1 U817 ( .A(n725), .B(KEYINPUT27), .ZN(n727) );
  AND2_X1 U818 ( .A1(G1956), .A2(n750), .ZN(n726) );
  NOR2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n734) );
  NOR2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U823 ( .A(n732), .B(KEYINPUT28), .Z(n733) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U825 ( .A(n735), .B(KEYINPUT29), .ZN(n738) );
  NOR2_X1 U826 ( .A1(G301), .A2(n736), .ZN(n737) );
  XNOR2_X1 U827 ( .A(KEYINPUT99), .B(n739), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n749) );
  XNOR2_X1 U829 ( .A(n749), .B(KEYINPUT101), .ZN(n742) );
  NOR2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n747) );
  INV_X1 U831 ( .A(n744), .ZN(n745) );
  NAND2_X1 U832 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U834 ( .A(n748), .B(KEYINPUT102), .ZN(n782) );
  XOR2_X1 U835 ( .A(KEYINPUT103), .B(KEYINPUT32), .Z(n758) );
  NAND2_X1 U836 ( .A1(G286), .A2(n749), .ZN(n755) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n787), .ZN(n752) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n750), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n753), .A2(G303), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U842 ( .A1(G8), .A2(n756), .ZN(n757) );
  XNOR2_X1 U843 ( .A(n758), .B(n757), .ZN(n781) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n984) );
  INV_X1 U845 ( .A(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n984), .A2(n759), .ZN(n760) );
  INV_X1 U847 ( .A(n787), .ZN(n765) );
  INV_X1 U848 ( .A(n765), .ZN(n779) );
  NOR2_X1 U849 ( .A1(n760), .A2(n779), .ZN(n762) );
  AND2_X1 U850 ( .A1(n781), .A2(n762), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n782), .A2(n761), .ZN(n771) );
  INV_X1 U852 ( .A(n762), .ZN(n764) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NOR2_X1 U854 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U855 ( .A1(n766), .A2(n763), .ZN(n999) );
  OR2_X1 U856 ( .A1(n764), .A2(n999), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U858 ( .A1(n767), .A2(KEYINPUT33), .ZN(n768) );
  AND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n773) );
  XNOR2_X1 U861 ( .A(n773), .B(n772), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n997), .A2(n774), .ZN(n775) );
  XNOR2_X1 U863 ( .A(n775), .B(KEYINPUT105), .ZN(n790) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U865 ( .A(n776), .B(KEYINPUT94), .Z(n777) );
  XNOR2_X1 U866 ( .A(KEYINPUT24), .B(n777), .ZN(n778) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U868 ( .A(n780), .B(KEYINPUT95), .ZN(n789) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n785) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G8), .A2(n783), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G131), .A2(n896), .ZN(n792) );
  NAND2_X1 U875 ( .A1(G95), .A2(n899), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U877 ( .A1(G119), .A2(n890), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G107), .A2(n892), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U880 ( .A1(n796), .A2(n795), .ZN(n907) );
  XNOR2_X1 U881 ( .A(KEYINPUT91), .B(G1991), .ZN(n938) );
  NOR2_X1 U882 ( .A1(n907), .A2(n938), .ZN(n805) );
  NAND2_X1 U883 ( .A1(G129), .A2(n890), .ZN(n798) );
  NAND2_X1 U884 ( .A1(G117), .A2(n892), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U886 ( .A1(n899), .A2(G105), .ZN(n799) );
  XOR2_X1 U887 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n896), .A2(G141), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n911) );
  AND2_X1 U891 ( .A1(G1996), .A2(n911), .ZN(n804) );
  NOR2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n963) );
  NOR2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n833) );
  INV_X1 U894 ( .A(n833), .ZN(n808) );
  NOR2_X1 U895 ( .A1(n963), .A2(n808), .ZN(n826) );
  XOR2_X1 U896 ( .A(KEYINPUT92), .B(n826), .Z(n820) );
  NAND2_X1 U897 ( .A1(G140), .A2(n896), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G104), .A2(n899), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n812) );
  XOR2_X1 U900 ( .A(KEYINPUT89), .B(KEYINPUT34), .Z(n811) );
  XNOR2_X1 U901 ( .A(n812), .B(n811), .ZN(n818) );
  NAND2_X1 U902 ( .A1(n890), .A2(G128), .ZN(n813) );
  XNOR2_X1 U903 ( .A(n813), .B(KEYINPUT90), .ZN(n815) );
  NAND2_X1 U904 ( .A1(G116), .A2(n892), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U906 ( .A(KEYINPUT35), .B(n816), .Z(n817) );
  NOR2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U908 ( .A(KEYINPUT36), .B(n819), .ZN(n914) );
  XNOR2_X1 U909 ( .A(KEYINPUT37), .B(G2067), .ZN(n831) );
  NOR2_X1 U910 ( .A1(n914), .A2(n831), .ZN(n977) );
  NAND2_X1 U911 ( .A1(n833), .A2(n977), .ZN(n829) );
  NAND2_X1 U912 ( .A1(n820), .A2(n829), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n526), .A2(n821), .ZN(n823) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U915 ( .A1(n987), .A2(n833), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n836) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n911), .ZN(n958) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n824) );
  AND2_X1 U919 ( .A1(n938), .A2(n907), .ZN(n961) );
  NOR2_X1 U920 ( .A1(n824), .A2(n961), .ZN(n825) );
  NOR2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U922 ( .A1(n958), .A2(n827), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n828), .B(KEYINPUT39), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n914), .A2(n831), .ZN(n966) );
  NAND2_X1 U926 ( .A1(n832), .A2(n966), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U929 ( .A(n837), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U930 ( .A(G223), .ZN(n838) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U933 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  INV_X1 U938 ( .A(n842), .ZN(n843) );
  NAND2_X1 U939 ( .A1(n844), .A2(n843), .ZN(G261) );
  INV_X1 U940 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U941 ( .A(G1991), .B(G2474), .ZN(n854) );
  XOR2_X1 U942 ( .A(G1981), .B(G1966), .Z(n846) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1956), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U945 ( .A(G1976), .B(G1961), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1971), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U949 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(G229) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2090), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n855), .B(KEYINPUT108), .ZN(n865) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2678), .Z(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT43), .B(G2096), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U957 ( .A(G2100), .B(G2084), .Z(n859) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2072), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U960 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U961 ( .A(KEYINPUT107), .B(KEYINPUT109), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(G227) );
  XNOR2_X1 U964 ( .A(n991), .B(n866), .ZN(n868) );
  XNOR2_X1 U965 ( .A(G171), .B(n988), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U967 ( .A(G286), .B(n869), .Z(n870) );
  NOR2_X1 U968 ( .A1(G37), .A2(n870), .ZN(G397) );
  NAND2_X1 U969 ( .A1(G112), .A2(n892), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G100), .A2(n899), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n878) );
  NAND2_X1 U972 ( .A1(n890), .A2(G124), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G136), .A2(n896), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U976 ( .A(KEYINPUT111), .B(n876), .Z(n877) );
  NOR2_X1 U977 ( .A1(n878), .A2(n877), .ZN(G162) );
  XOR2_X1 U978 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n880) );
  XNOR2_X1 U979 ( .A(G162), .B(KEYINPUT46), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n906) );
  NAND2_X1 U981 ( .A1(G106), .A2(n899), .ZN(n881) );
  XOR2_X1 U982 ( .A(KEYINPUT113), .B(n881), .Z(n883) );
  NAND2_X1 U983 ( .A1(n896), .A2(G142), .ZN(n882) );
  NAND2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n884), .B(KEYINPUT45), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G130), .A2(n890), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G118), .A2(n892), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT112), .B(n887), .Z(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n904) );
  NAND2_X1 U991 ( .A1(n890), .A2(G127), .ZN(n891) );
  XOR2_X1 U992 ( .A(KEYINPUT115), .B(n891), .Z(n894) );
  NAND2_X1 U993 ( .A1(n892), .A2(G115), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n895), .B(KEYINPUT47), .ZN(n898) );
  NAND2_X1 U996 ( .A1(G139), .A2(n896), .ZN(n897) );
  NAND2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n902) );
  NAND2_X1 U998 ( .A1(n899), .A2(G103), .ZN(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT114), .B(n900), .Z(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(KEYINPUT116), .B(n903), .Z(n968) );
  XNOR2_X1 U1002 ( .A(n904), .B(n968), .ZN(n905) );
  XOR2_X1 U1003 ( .A(n906), .B(n905), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G160), .B(n907), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n910), .B(n960), .Z(n913) );
  XOR2_X1 U1007 ( .A(G164), .B(n911), .Z(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(KEYINPUT118), .B(n917), .ZN(G395) );
  XOR2_X1 U1012 ( .A(G2443), .B(G2427), .Z(n919) );
  XNOR2_X1 U1013 ( .A(G2438), .B(G2454), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1015 ( .A(n920), .B(G2435), .Z(n922) );
  XNOR2_X1 U1016 ( .A(G1348), .B(G1341), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(n926) );
  XOR2_X1 U1018 ( .A(G2430), .B(G2446), .Z(n924) );
  XNOR2_X1 U1019 ( .A(KEYINPUT106), .B(G2451), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1021 ( .A(n926), .B(n925), .Z(n927) );
  NAND2_X1 U1022 ( .A1(G14), .A2(n927), .ZN(n933) );
  NAND2_X1 U1023 ( .A1(G319), .A2(n933), .ZN(n930) );
  NOR2_X1 U1024 ( .A1(G229), .A2(G227), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT49), .B(n928), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(G397), .A2(G395), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(G69), .ZN(G235) );
  INV_X1 U1031 ( .A(n933), .ZN(G401) );
  XNOR2_X1 U1032 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n956) );
  XNOR2_X1 U1033 ( .A(G32), .B(n934), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n935), .A2(G28), .ZN(n945) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n943) );
  XOR2_X1 U1038 ( .A(n938), .B(G25), .Z(n941) );
  XNOR2_X1 U1039 ( .A(n939), .B(G27), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(KEYINPUT53), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(n947), .B(KEYINPUT121), .ZN(n950) );
  XOR2_X1 U1045 ( .A(G2084), .B(G34), .Z(n948) );
  XNOR2_X1 U1046 ( .A(KEYINPUT54), .B(n948), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT120), .B(G2090), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(G35), .B(n951), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  OR2_X1 U1051 ( .A1(G29), .A2(n954), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(n956), .B(n955), .ZN(n980) );
  XOR2_X1 U1053 ( .A(G2090), .B(G162), .Z(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1055 ( .A(KEYINPUT51), .B(n959), .Z(n975) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1058 ( .A(G160), .B(G2084), .Z(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n973) );
  XOR2_X1 U1061 ( .A(G164), .B(G2078), .Z(n970) );
  XNOR2_X1 U1062 ( .A(G2072), .B(n968), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1064 ( .A(KEYINPUT50), .B(n971), .Z(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1068 ( .A(n978), .B(KEYINPUT52), .Z(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n524), .ZN(n1034) );
  XOR2_X1 U1070 ( .A(G16), .B(KEYINPUT56), .Z(n981) );
  XNOR2_X1 U1071 ( .A(KEYINPUT122), .B(n981), .ZN(n1004) );
  XNOR2_X1 U1072 ( .A(G301), .B(G1961), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(G299), .B(G1956), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n995) );
  XNOR2_X1 U1077 ( .A(n988), .B(G1348), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(G1971), .A2(G303), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G1341), .B(n991), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n1002) );
  XOR2_X1 U1083 ( .A(G1966), .B(G168), .Z(n996) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1085 ( .A(KEYINPUT57), .B(n998), .Z(n1000) );
  NAND2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1087 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1088 ( .A1(n1004), .A2(n1003), .ZN(n1031) );
  XNOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(n1005), .B(G4), .ZN(n1009) );
  XNOR2_X1 U1091 ( .A(G1956), .B(G20), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G1981), .B(G6), .ZN(n1006) );
  NOR2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1095 ( .A(KEYINPUT123), .B(G1341), .Z(n1010) );
  XNOR2_X1 U1096 ( .A(G19), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1013), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1014), .B(KEYINPUT124), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(G1961), .B(G5), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1026) );
  XNOR2_X1 U1104 ( .A(G1986), .B(G24), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(G22), .B(G1971), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(G1976), .B(KEYINPUT125), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1021), .B(G23), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT58), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1027), .Z(n1028) );
  NOR2_X1 U1113 ( .A1(G16), .A2(n1028), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(n1029), .B(KEYINPUT126), .ZN(n1030) );
  NOR2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1116 ( .A(n1032), .B(KEYINPUT127), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1035), .A2(G11), .ZN(n1036) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1036), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

