

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  XNOR2_X1 U324 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U325 ( .A(n359), .B(n358), .Z(n292) );
  XOR2_X1 U326 ( .A(G183GAT), .B(KEYINPUT17), .Z(n293) );
  XOR2_X1 U327 ( .A(n433), .B(n372), .Z(n294) );
  INV_X1 U328 ( .A(KEYINPUT93), .ZN(n398) );
  XNOR2_X1 U329 ( .A(n548), .B(n398), .ZN(n401) );
  INV_X1 U330 ( .A(KEYINPUT119), .ZN(n467) );
  XNOR2_X1 U331 ( .A(n467), .B(KEYINPUT54), .ZN(n468) );
  XNOR2_X1 U332 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U333 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U334 ( .A(n360), .B(n292), .ZN(n361) );
  NOR2_X1 U335 ( .A1(n472), .A2(n520), .ZN(n395) );
  XNOR2_X1 U336 ( .A(n362), .B(n361), .ZN(n364) );
  NOR2_X1 U337 ( .A1(n399), .A2(n475), .ZN(n568) );
  XNOR2_X1 U338 ( .A(KEYINPUT99), .B(n452), .ZN(n498) );
  XNOR2_X1 U339 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n476) );
  XNOR2_X1 U340 ( .A(G36GAT), .B(KEYINPUT100), .ZN(n453) );
  XNOR2_X1 U341 ( .A(n477), .B(n476), .ZN(G1350GAT) );
  XNOR2_X1 U342 ( .A(n454), .B(n453), .ZN(G1329GAT) );
  XOR2_X1 U343 ( .A(G78GAT), .B(G64GAT), .Z(n296) );
  XNOR2_X1 U344 ( .A(G183GAT), .B(G71GAT), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U346 ( .A(n297), .B(G211GAT), .Z(n299) );
  XOR2_X1 U347 ( .A(KEYINPUT13), .B(G57GAT), .Z(n432) );
  XNOR2_X1 U348 ( .A(G8GAT), .B(n432), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n305) );
  XOR2_X1 U350 ( .A(G1GAT), .B(G15GAT), .Z(n301) );
  XNOR2_X1 U351 ( .A(KEYINPUT68), .B(G22GAT), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n441) );
  XOR2_X1 U353 ( .A(G127GAT), .B(n441), .Z(n303) );
  NAND2_X1 U354 ( .A1(G231GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U356 ( .A(n305), .B(n304), .Z(n313) );
  XOR2_X1 U357 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n307) );
  XNOR2_X1 U358 ( .A(KEYINPUT77), .B(KEYINPUT76), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U360 ( .A(G155GAT), .B(KEYINPUT12), .Z(n309) );
  XNOR2_X1 U361 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U364 ( .A(n313), .B(n312), .Z(n584) );
  INV_X1 U365 ( .A(n584), .ZN(n538) );
  XOR2_X1 U366 ( .A(G50GAT), .B(G162GAT), .Z(n377) );
  XNOR2_X1 U367 ( .A(G36GAT), .B(G190GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n314), .B(G218GAT), .ZN(n369) );
  XOR2_X1 U369 ( .A(G92GAT), .B(n369), .Z(n316) );
  NAND2_X1 U370 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n377), .B(n317), .ZN(n321) );
  XOR2_X1 U373 ( .A(G29GAT), .B(G43GAT), .Z(n319) );
  XNOR2_X1 U374 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n442) );
  XOR2_X1 U376 ( .A(G99GAT), .B(G85GAT), .Z(n416) );
  XOR2_X1 U377 ( .A(n442), .B(n416), .Z(n320) );
  XNOR2_X1 U378 ( .A(n321), .B(n320), .ZN(n329) );
  XOR2_X1 U379 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n323) );
  XNOR2_X1 U380 ( .A(KEYINPUT10), .B(KEYINPUT65), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U382 ( .A(KEYINPUT9), .B(KEYINPUT73), .Z(n325) );
  XNOR2_X1 U383 ( .A(G134GAT), .B(G106GAT), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U385 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n567) );
  XOR2_X1 U387 ( .A(KEYINPUT36), .B(n567), .Z(n589) );
  XOR2_X1 U388 ( .A(KEYINPUT0), .B(G127GAT), .Z(n331) );
  XNOR2_X1 U389 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n333) );
  XOR2_X1 U391 ( .A(G113GAT), .B(G134GAT), .Z(n332) );
  XOR2_X1 U392 ( .A(n333), .B(n332), .Z(n363) );
  XOR2_X1 U393 ( .A(KEYINPUT4), .B(G148GAT), .Z(n335) );
  XNOR2_X1 U394 ( .A(G1GAT), .B(G120GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U396 ( .A(KEYINPUT6), .B(KEYINPUT87), .Z(n337) );
  XNOR2_X1 U397 ( .A(KEYINPUT88), .B(KEYINPUT5), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U399 ( .A(n339), .B(n338), .Z(n351) );
  XNOR2_X1 U400 ( .A(KEYINPUT2), .B(KEYINPUT85), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n340), .B(KEYINPUT3), .ZN(n341) );
  XOR2_X1 U402 ( .A(n341), .B(KEYINPUT86), .Z(n343) );
  XNOR2_X1 U403 ( .A(G141GAT), .B(G155GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n389) );
  XOR2_X1 U405 ( .A(G162GAT), .B(G85GAT), .Z(n345) );
  XNOR2_X1 U406 ( .A(G29GAT), .B(G57GAT), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U408 ( .A(KEYINPUT1), .B(n346), .Z(n348) );
  NAND2_X1 U409 ( .A1(G225GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n389), .B(n349), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n363), .B(n352), .ZN(n545) );
  XOR2_X1 U414 ( .A(G120GAT), .B(G71GAT), .Z(n433) );
  XNOR2_X1 U415 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n293), .B(n353), .ZN(n372) );
  XNOR2_X1 U417 ( .A(G190GAT), .B(G99GAT), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n294), .B(n354), .ZN(n362) );
  XOR2_X1 U419 ( .A(G176GAT), .B(G15GAT), .Z(n356) );
  XNOR2_X1 U420 ( .A(G169GAT), .B(G43GAT), .ZN(n355) );
  XNOR2_X1 U421 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n357), .B(KEYINPUT82), .ZN(n360) );
  XOR2_X1 U423 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n359) );
  NAND2_X1 U424 ( .A1(G227GAT), .A2(G233GAT), .ZN(n358) );
  XOR2_X1 U425 ( .A(n364), .B(n363), .Z(n399) );
  INV_X1 U426 ( .A(n399), .ZN(n520) );
  XOR2_X1 U427 ( .A(G169GAT), .B(G8GAT), .Z(n445) );
  XOR2_X1 U428 ( .A(KEYINPUT89), .B(n445), .Z(n366) );
  NAND2_X1 U429 ( .A1(G226GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n376) );
  XOR2_X1 U431 ( .A(KEYINPUT21), .B(KEYINPUT84), .Z(n368) );
  XNOR2_X1 U432 ( .A(G197GAT), .B(G211GAT), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n381) );
  XOR2_X1 U434 ( .A(n381), .B(n369), .Z(n374) );
  XOR2_X1 U435 ( .A(G64GAT), .B(G204GAT), .Z(n371) );
  XNOR2_X1 U436 ( .A(G176GAT), .B(G92GAT), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n425) );
  XNOR2_X1 U438 ( .A(n372), .B(n425), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U440 ( .A(n376), .B(n375), .Z(n517) );
  NAND2_X1 U441 ( .A1(n520), .A2(n517), .ZN(n392) );
  XOR2_X1 U442 ( .A(n377), .B(G218GAT), .Z(n380) );
  XNOR2_X1 U443 ( .A(G106GAT), .B(G78GAT), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n378), .B(G148GAT), .ZN(n417) );
  XNOR2_X1 U445 ( .A(G204GAT), .B(n417), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n385) );
  XOR2_X1 U447 ( .A(n381), .B(KEYINPUT22), .Z(n383) );
  NAND2_X1 U448 ( .A1(G228GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U450 ( .A(n385), .B(n384), .Z(n391) );
  XOR2_X1 U451 ( .A(KEYINPUT23), .B(KEYINPUT83), .Z(n387) );
  XNOR2_X1 U452 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n472) );
  NAND2_X1 U456 ( .A1(n392), .A2(n472), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n393), .B(KEYINPUT25), .ZN(n403) );
  XNOR2_X1 U458 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n574) );
  XNOR2_X1 U460 ( .A(n517), .B(KEYINPUT90), .ZN(n396) );
  XOR2_X1 U461 ( .A(n396), .B(KEYINPUT27), .Z(n405) );
  INV_X1 U462 ( .A(n405), .ZN(n397) );
  NAND2_X1 U463 ( .A1(n574), .A2(n397), .ZN(n548) );
  NAND2_X1 U464 ( .A1(n399), .A2(KEYINPUT91), .ZN(n400) );
  NAND2_X1 U465 ( .A1(n401), .A2(n400), .ZN(n402) );
  NOR2_X1 U466 ( .A1(n403), .A2(n402), .ZN(n404) );
  NOR2_X1 U467 ( .A1(n545), .A2(n404), .ZN(n412) );
  INV_X1 U468 ( .A(KEYINPUT91), .ZN(n406) );
  XOR2_X1 U469 ( .A(n472), .B(KEYINPUT28), .Z(n523) );
  NOR2_X1 U470 ( .A1(n523), .A2(n405), .ZN(n407) );
  NAND2_X1 U471 ( .A1(n407), .A2(n545), .ZN(n528) );
  NAND2_X1 U472 ( .A1(n406), .A2(n528), .ZN(n409) );
  NAND2_X1 U473 ( .A1(n407), .A2(KEYINPUT91), .ZN(n408) );
  NAND2_X1 U474 ( .A1(n409), .A2(n408), .ZN(n410) );
  NOR2_X1 U475 ( .A1(n410), .A2(n520), .ZN(n411) );
  NOR2_X1 U476 ( .A1(n412), .A2(n411), .ZN(n481) );
  NOR2_X1 U477 ( .A1(n589), .A2(n481), .ZN(n413) );
  NAND2_X1 U478 ( .A1(n538), .A2(n413), .ZN(n414) );
  XNOR2_X1 U479 ( .A(KEYINPUT98), .B(n414), .ZN(n415) );
  XNOR2_X1 U480 ( .A(n415), .B(KEYINPUT37), .ZN(n514) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n421) );
  INV_X1 U482 ( .A(n421), .ZN(n419) );
  AND2_X1 U483 ( .A1(G230GAT), .A2(G233GAT), .ZN(n420) );
  INV_X1 U484 ( .A(n420), .ZN(n418) );
  NAND2_X1 U485 ( .A1(n419), .A2(n418), .ZN(n423) );
  NAND2_X1 U486 ( .A1(n421), .A2(n420), .ZN(n422) );
  NAND2_X1 U487 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n424), .B(KEYINPUT32), .ZN(n431) );
  XOR2_X1 U489 ( .A(n425), .B(KEYINPUT31), .Z(n429) );
  XOR2_X1 U490 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n427) );
  XNOR2_X1 U491 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U493 ( .A(n433), .B(n432), .Z(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n580) );
  XOR2_X1 U495 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n437) );
  XNOR2_X1 U496 ( .A(G197GAT), .B(KEYINPUT67), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n450) );
  XOR2_X1 U498 ( .A(G141GAT), .B(G113GAT), .Z(n439) );
  NAND2_X1 U499 ( .A1(G229GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U501 ( .A(n440), .B(KEYINPUT29), .Z(n444) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n446) );
  XOR2_X1 U504 ( .A(n446), .B(n445), .Z(n448) );
  XNOR2_X1 U505 ( .A(G50GAT), .B(G36GAT), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n575) );
  NOR2_X1 U508 ( .A1(n580), .A2(n575), .ZN(n482) );
  NAND2_X1 U509 ( .A1(n514), .A2(n482), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n451), .B(KEYINPUT38), .ZN(n452) );
  NAND2_X1 U511 ( .A1(n498), .A2(n517), .ZN(n454) );
  XNOR2_X1 U512 ( .A(KEYINPUT118), .B(n517), .ZN(n466) );
  INV_X1 U513 ( .A(n575), .ZN(n560) );
  INV_X1 U514 ( .A(KEYINPUT41), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n580), .B(n455), .ZN(n563) );
  NAND2_X1 U516 ( .A1(n560), .A2(n563), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n456), .B(KEYINPUT46), .ZN(n458) );
  INV_X1 U518 ( .A(n567), .ZN(n542) );
  AND2_X1 U519 ( .A1(n538), .A2(n542), .ZN(n457) );
  AND2_X1 U520 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U521 ( .A(n459), .B(KEYINPUT47), .ZN(n464) );
  NOR2_X1 U522 ( .A1(n538), .A2(n589), .ZN(n460) );
  XOR2_X1 U523 ( .A(KEYINPUT45), .B(n460), .Z(n461) );
  NOR2_X1 U524 ( .A1(n580), .A2(n461), .ZN(n462) );
  NAND2_X1 U525 ( .A1(n462), .A2(n575), .ZN(n463) );
  NAND2_X1 U526 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U527 ( .A(KEYINPUT48), .B(n465), .ZN(n546) );
  NAND2_X1 U528 ( .A1(n466), .A2(n546), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n545), .A2(n470), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT64), .ZN(n573) );
  NAND2_X1 U531 ( .A1(n573), .A2(n472), .ZN(n474) );
  XOR2_X1 U532 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n584), .A2(n568), .ZN(n477) );
  NAND2_X1 U535 ( .A1(n584), .A2(n542), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT16), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n479), .B(KEYINPUT78), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n481), .A2(n480), .ZN(n501) );
  NAND2_X1 U539 ( .A1(n501), .A2(n482), .ZN(n483) );
  XOR2_X1 U540 ( .A(KEYINPUT94), .B(n483), .Z(n490) );
  NAND2_X1 U541 ( .A1(n490), .A2(n545), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(KEYINPUT34), .ZN(n485) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U544 ( .A1(n490), .A2(n517), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT35), .B(KEYINPUT95), .Z(n488) );
  NAND2_X1 U547 ( .A1(n490), .A2(n520), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U549 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n492) );
  NAND2_X1 U551 ( .A1(n523), .A2(n490), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G22GAT), .B(n493), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U555 ( .A1(n498), .A2(n545), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n498), .A2(n520), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n523), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U562 ( .A(n563), .ZN(n533) );
  NOR2_X1 U563 ( .A1(n533), .A2(n560), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(KEYINPUT102), .ZN(n513) );
  NAND2_X1 U565 ( .A1(n513), .A2(n501), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(KEYINPUT103), .ZN(n510) );
  NAND2_X1 U567 ( .A1(n545), .A2(n510), .ZN(n505) );
  XOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT101), .Z(n503) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n510), .A2(n517), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(KEYINPUT104), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  XOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT105), .Z(n509) );
  NAND2_X1 U575 ( .A1(n510), .A2(n520), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U578 ( .A1(n510), .A2(n523), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  AND2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n524) );
  NAND2_X1 U581 ( .A1(n524), .A2(n545), .ZN(n515) );
  XNOR2_X1 U582 ( .A(KEYINPUT106), .B(n515), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  XOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT107), .Z(n519) );
  NAND2_X1 U585 ( .A1(n524), .A2(n517), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n520), .A2(n524), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(KEYINPUT108), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n526) );
  NAND2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n399), .A2(n528), .ZN(n529) );
  NAND2_X1 U595 ( .A1(n546), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(KEYINPUT110), .B(n530), .ZN(n541) );
  NOR2_X1 U597 ( .A1(n541), .A2(n575), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(KEYINPUT111), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  NOR2_X1 U600 ( .A1(n533), .A2(n541), .ZN(n537) );
  XOR2_X1 U601 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n535) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT113), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n541), .ZN(n539) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(n539), .Z(n540) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n544) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n557), .A2(n560), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(KEYINPUT114), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n552) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U619 ( .A(KEYINPUT115), .B(n553), .Z(n555) );
  NAND2_X1 U620 ( .A1(n557), .A2(n563), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n584), .A2(n557), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U624 ( .A(G162GAT), .B(KEYINPUT117), .Z(n559) );
  NAND2_X1 U625 ( .A1(n557), .A2(n567), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1347GAT) );
  XOR2_X1 U627 ( .A(G169GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U628 ( .A1(n568), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n568), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1351GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n588) );
  NOR2_X1 U640 ( .A1(n588), .A2(n575), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U646 ( .A(n588), .ZN(n585) );
  NAND2_X1 U647 ( .A1(n585), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

