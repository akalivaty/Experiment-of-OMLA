//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n634, new_n636, new_n637, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1247, new_n1248;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .A3(G101), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n463), .A2(G137), .A3(new_n462), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n466), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n463), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n462), .B1(new_n478), .B2(new_n480), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(new_n462), .A2(G138), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n463), .A2(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n463), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n494), .A2(new_n500), .A3(new_n501), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(G50), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(KEYINPUT72), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT6), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n514), .A2(new_n524), .ZN(G166));
  OR2_X1    g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n532), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n528), .A2(new_n529), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n523), .A2(new_n528), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT74), .B(G51), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n521), .A2(KEYINPUT6), .A3(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(KEYINPUT6), .B1(new_n521), .B2(G651), .ZN(new_n540));
  OAI21_X1  g115(.A(KEYINPUT73), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n520), .A2(new_n542), .A3(new_n522), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n541), .A2(G543), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n537), .B1(new_n538), .B2(new_n544), .ZN(G168));
  NAND4_X1  g120(.A1(new_n541), .A2(G52), .A3(G543), .A4(new_n543), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n520), .A2(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n526), .B2(new_n527), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT75), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n556), .B(new_n553), .C1(new_n511), .C2(new_n551), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(G651), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n550), .A2(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  INV_X1    g135(.A(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n523), .B2(KEYINPUT73), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n562), .A2(G43), .A3(new_n543), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G56), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n511), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n547), .B2(G81), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  NAND4_X1  g149(.A1(new_n541), .A2(G53), .A3(G543), .A4(new_n543), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n562), .A2(KEYINPUT9), .A3(G53), .A4(new_n543), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n511), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n547), .B2(G91), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND3_X1  g160(.A1(new_n562), .A2(G49), .A3(new_n543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n547), .A2(KEYINPUT76), .A3(G87), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT76), .B1(new_n547), .B2(G87), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(G288));
  OAI21_X1  g165(.A(G61), .B1(new_n509), .B2(new_n510), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n519), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(KEYINPUT77), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  AOI211_X1 g170(.A(new_n595), .B(new_n519), .C1(new_n591), .C2(new_n592), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G48), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n511), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(new_n523), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(new_n544), .A2(G47), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n547), .A2(G85), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  INV_X1    g182(.A(G72), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n511), .A2(new_n607), .B1(new_n608), .B2(new_n561), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n605), .B(new_n606), .C1(new_n611), .C2(new_n613), .ZN(G290));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NOR2_X1   g190(.A1(G301), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n562), .A2(G54), .A3(new_n543), .ZN(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT79), .B(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n511), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G651), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n547), .A2(KEYINPUT10), .A3(G92), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT10), .B1(new_n547), .B2(G92), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n617), .B(new_n621), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(KEYINPUT80), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(KEYINPUT80), .ZN(new_n627));
  AND2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n616), .B1(new_n628), .B2(new_n615), .ZN(G284));
  AOI21_X1  g204(.A(new_n616), .B1(new_n628), .B2(new_n615), .ZN(G321));
  NAND2_X1  g205(.A1(G299), .A2(new_n615), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n615), .B2(G168), .ZN(G297));
  OAI21_X1  g207(.A(new_n631), .B1(new_n615), .B2(G168), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n628), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n568), .A2(new_n615), .ZN(new_n636));
  AND3_X1   g211(.A1(new_n626), .A2(new_n634), .A3(new_n627), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(new_n615), .ZN(G323));
  XOR2_X1   g213(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n639));
  XNOR2_X1  g214(.A(G323), .B(new_n639), .ZN(G282));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(KEYINPUT83), .ZN(new_n642));
  INV_X1    g217(.A(G111), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n641), .A2(KEYINPUT83), .B1(new_n643), .B2(G2105), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n481), .A2(G135), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n483), .A2(new_n646), .A3(G123), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n646), .B1(new_n483), .B2(G123), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2096), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT13), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(G156));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT84), .ZN(new_n670));
  OAI21_X1  g245(.A(G14), .B1(new_n667), .B2(new_n668), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(G401));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT85), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  XOR2_X1   g254(.A(new_n676), .B(KEYINPUT86), .Z(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n680), .B2(new_n674), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n674), .B(KEYINPUT17), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(new_n680), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n680), .A3(new_n677), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT19), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n691), .A2(new_n692), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(new_n698), .B(new_n697), .S(new_n690), .Z(new_n699));
  NOR2_X1   g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT87), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(G229));
  INV_X1    g282(.A(KEYINPUT101), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G6), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n603), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT32), .B(G1981), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n712), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n714), .B(new_n710), .C1(new_n603), .C2(new_n709), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n709), .A2(G22), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n717), .B(new_n718), .C1(G166), .C2(new_n709), .ZN(new_n719));
  INV_X1    g294(.A(G1971), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n709), .B1(new_n514), .B2(new_n524), .ZN(new_n721));
  INV_X1    g296(.A(new_n718), .ZN(new_n722));
  OAI21_X1  g297(.A(KEYINPUT91), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n719), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n720), .B1(new_n719), .B2(new_n723), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n716), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G23), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT89), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G288), .B2(new_n709), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT33), .B(G1976), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n727), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT34), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n727), .A2(new_n740), .A3(new_n736), .A4(new_n737), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  OR2_X1    g317(.A1(G95), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT88), .Z(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G119), .B2(new_n483), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n481), .A2(G131), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n742), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT35), .B(G1991), .Z(new_n749));
  AND2_X1   g324(.A1(new_n742), .A2(G25), .ZN(new_n750));
  OR3_X1    g325(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n709), .A2(G24), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G290), .B2(G16), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G1986), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G1986), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n751), .A2(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n741), .A2(KEYINPUT92), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(KEYINPUT92), .B1(new_n741), .B2(new_n757), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n739), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(KEYINPUT93), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n739), .B1(KEYINPUT93), .B2(new_n762), .C1(new_n759), .C2(new_n760), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n709), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n481), .A2(G140), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n483), .A2(G128), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n462), .A2(G116), .ZN(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n771), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AND3_X1   g350(.A1(new_n775), .A2(KEYINPUT94), .A3(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(KEYINPUT94), .B1(new_n775), .B2(G29), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n742), .A2(G26), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT28), .ZN(new_n780));
  AOI21_X1  g355(.A(G2067), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(G2067), .B(new_n780), .C1(new_n776), .C2(new_n777), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n770), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n709), .A2(G4), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n628), .B2(new_n709), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1348), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n742), .A2(G35), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n487), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT29), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  OAI21_X1  g369(.A(G2090), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n794), .ZN(new_n796));
  INV_X1    g371(.A(G2090), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n796), .A2(new_n797), .A3(new_n792), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n709), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n569), .B2(new_n709), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G1341), .Z(new_n801));
  NAND3_X1  g376(.A1(new_n795), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n784), .A2(new_n787), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n709), .A2(G21), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G168), .B2(new_n709), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G1966), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT97), .ZN(new_n808));
  OR2_X1    g383(.A1(G29), .A2(G33), .ZN(new_n809));
  NAND2_X1  g384(.A1(G115), .A2(G2104), .ZN(new_n810));
  INV_X1    g385(.A(G127), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n477), .B2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n462), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT25), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n481), .B2(G139), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n809), .B1(new_n819), .B2(new_n742), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT96), .B(G2072), .Z(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n742), .A2(G27), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n506), .B2(G29), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT99), .B(G2078), .Z(new_n825));
  AOI22_X1  g400(.A1(new_n820), .A2(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n808), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G34), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT24), .ZN(new_n829));
  AOI21_X1  g404(.A(G29), .B1(new_n828), .B2(KEYINPUT24), .ZN(new_n830));
  AOI22_X1  g405(.A1(G160), .A2(G29), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n831), .A2(G2084), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(G2084), .ZN(new_n833));
  INV_X1    g408(.A(G28), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT30), .ZN(new_n835));
  AOI21_X1  g410(.A(G29), .B1(new_n834), .B2(KEYINPUT30), .ZN(new_n836));
  OR2_X1    g411(.A1(KEYINPUT31), .A2(G11), .ZN(new_n837));
  NAND2_X1  g412(.A1(KEYINPUT31), .A2(G11), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n832), .A2(new_n833), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g415(.A(G29), .B(new_n645), .C1(new_n647), .C2(new_n648), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n824), .A2(new_n825), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n806), .A2(G1966), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n709), .A2(G5), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G301), .B2(G16), .ZN(new_n846));
  INV_X1    g421(.A(G1961), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n742), .A2(G32), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n481), .A2(G141), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n483), .A2(G129), .ZN(new_n851));
  NAND3_X1  g426(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT26), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n854), .A2(new_n855), .B1(G105), .B2(new_n468), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n849), .B1(new_n857), .B2(G29), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT27), .B(G1996), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n858), .A2(new_n860), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n848), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n827), .A2(new_n844), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n846), .A2(new_n847), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT98), .Z(new_n866));
  AOI21_X1  g441(.A(new_n804), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n844), .A2(new_n863), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n808), .A2(new_n822), .A3(new_n826), .ZN(new_n869));
  AND4_X1   g444(.A1(new_n804), .A2(new_n868), .A3(new_n869), .A4(new_n866), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n803), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n708), .B1(new_n766), .B2(new_n872), .ZN(new_n873));
  AOI211_X1 g448(.A(KEYINPUT101), .B(new_n871), .C1(new_n764), .C2(new_n765), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(G311));
  NAND2_X1  g450(.A1(new_n766), .A2(new_n872), .ZN(G150));
  NAND3_X1  g451(.A1(new_n562), .A2(G55), .A3(new_n543), .ZN(new_n877));
  NAND2_X1  g452(.A1(G80), .A2(G543), .ZN(new_n878));
  INV_X1    g453(.A(G67), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n511), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n880), .A2(G651), .B1(new_n547), .B2(G93), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n628), .A2(G559), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT102), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n568), .A2(new_n882), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n563), .A2(new_n567), .A3(new_n877), .A4(new_n881), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n887), .B(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n891), .A2(KEYINPUT39), .ZN(new_n892));
  INV_X1    g467(.A(G860), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n891), .B2(KEYINPUT39), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n884), .B1(new_n892), .B2(new_n894), .ZN(G145));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n746), .A2(new_n747), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n653), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n819), .B(new_n857), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n775), .B(new_n502), .Z(new_n903));
  NAND2_X1  g478(.A1(new_n481), .A2(G142), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n483), .A2(G130), .ZN(new_n905));
  OAI21_X1  g480(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n907));
  INV_X1    g482(.A(G118), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n906), .A2(new_n907), .B1(new_n908), .B2(G2105), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n907), .B2(new_n906), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n904), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n903), .A2(new_n911), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n902), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n900), .A2(new_n912), .A3(new_n913), .A4(new_n901), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n487), .B(G160), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n918), .B(new_n649), .Z(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n896), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT104), .A4(new_n919), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n917), .B2(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g501(.A1(new_n882), .A2(new_n615), .ZN(new_n927));
  INV_X1    g502(.A(G288), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(new_n603), .ZN(new_n929));
  XNOR2_X1  g504(.A(G290), .B(G303), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(G290), .B(G166), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n603), .B(G288), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n936));
  OR2_X1    g511(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n931), .A2(new_n934), .A3(KEYINPUT107), .A4(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n637), .B(new_n890), .ZN(new_n943));
  AND2_X1   g518(.A1(G299), .A2(new_n625), .ZN(new_n944));
  NOR2_X1   g519(.A1(G299), .A2(new_n625), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(KEYINPUT105), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n578), .A2(new_n582), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT10), .ZN(new_n951));
  INV_X1    g526(.A(G92), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n535), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n953), .A2(new_n622), .B1(G651), .B2(new_n620), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n950), .A2(new_n577), .A3(new_n617), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G299), .A2(new_n625), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n948), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n949), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n956), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT106), .B1(new_n961), .B2(KEYINPUT41), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n963));
  AOI211_X1 g538(.A(new_n963), .B(new_n948), .C1(new_n955), .C2(new_n956), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n943), .A2(new_n960), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n947), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(new_n941), .A3(new_n940), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n940), .A2(new_n941), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(new_n947), .A3(new_n966), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n942), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n927), .B1(new_n971), .B2(new_n615), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n974), .B(new_n927), .C1(new_n971), .C2(new_n615), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(G295));
  NAND2_X1  g551(.A1(new_n972), .A2(KEYINPUT110), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n927), .C1(new_n971), .C2(new_n615), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(G331));
  INV_X1    g555(.A(new_n935), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n550), .A2(KEYINPUT111), .A3(new_n558), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G168), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n555), .A2(G651), .A3(new_n557), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(new_n549), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n986), .A2(new_n888), .A3(new_n889), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n888), .B2(new_n889), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n890), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n982), .A2(G168), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n986), .A2(new_n888), .A3(new_n889), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(new_n946), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT112), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n989), .A2(new_n994), .A3(new_n997), .A4(new_n946), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n965), .A2(new_n960), .B1(new_n994), .B2(new_n989), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n981), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G37), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n989), .A2(new_n994), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n957), .B(KEYINPUT105), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT41), .B1(new_n944), .B2(new_n945), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n963), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n961), .A2(KEYINPUT106), .A3(KEYINPUT41), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1003), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(new_n935), .A3(new_n996), .A4(new_n998), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1001), .A2(new_n1002), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1003), .B1(KEYINPUT113), .B2(new_n1005), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1005), .A2(KEYINPUT113), .A3(new_n957), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n995), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n981), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1017), .A2(KEYINPUT43), .A3(new_n1002), .A4(new_n1010), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT44), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1010), .A2(new_n1002), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1012), .B1(new_n1022), .B2(new_n1001), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1017), .A2(new_n1012), .A3(new_n1002), .A4(new_n1010), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1020), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1021), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT44), .B1(new_n1030), .B2(new_n1024), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT114), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1028), .A2(new_n1032), .ZN(G397));
  INV_X1    g608(.A(G40), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n466), .A2(new_n475), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n502), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n775), .B(G2067), .Z(new_n1041));
  INV_X1    g616(.A(G1996), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n857), .B(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n746), .A2(new_n749), .A3(new_n747), .ZN(new_n1044));
  INV_X1    g619(.A(new_n749), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n897), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(G290), .B(G1986), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1040), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1035), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n502), .A2(KEYINPUT115), .A3(new_n1037), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT115), .B1(new_n502), .B2(new_n1037), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n506), .A2(new_n1037), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1036), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n1037), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1035), .ZN(new_n1062));
  INV_X1    g637(.A(G1966), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1059), .A2(new_n1064), .A3(KEYINPUT124), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT124), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1065), .A2(new_n1066), .A3(G286), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n1068));
  INV_X1    g643(.A(G8), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1069), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1072));
  NOR2_X1   g647(.A1(G168), .A2(new_n1069), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1068), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1067), .A2(new_n1071), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1059), .A2(new_n1064), .A3(KEYINPUT124), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1074), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1076), .A2(new_n1077), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1080), .A2(G168), .A3(new_n1081), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1086), .B2(new_n1070), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT62), .B1(new_n1087), .B2(new_n1082), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1038), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n502), .A2(KEYINPUT115), .A3(new_n1037), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1054), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1058), .A2(new_n1035), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n1037), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1035), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G2078), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1384), .B1(new_n503), .B2(new_n505), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1095), .B(new_n1096), .C1(KEYINPUT45), .C2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1093), .A2(new_n847), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1060), .A2(new_n1061), .A3(new_n1096), .A4(new_n1035), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1101), .A2(KEYINPUT125), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT53), .B1(new_n1101), .B2(KEYINPUT125), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1104), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT126), .B1(new_n1104), .B2(G171), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT118), .B(G1981), .Z(new_n1111));
  OAI211_X1 g686(.A(new_n601), .B(new_n1111), .C1(new_n594), .C2(new_n596), .ZN(new_n1112));
  OAI21_X1  g687(.A(G1981), .B1(new_n602), .B2(new_n593), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT49), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1110), .A2(new_n1069), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1113), .A3(KEYINPUT49), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1090), .A2(new_n1035), .A3(new_n1091), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n588), .A2(new_n589), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(G1976), .A3(new_n586), .A4(new_n587), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1119), .A3(G8), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1115), .A2(new_n1116), .B1(KEYINPUT52), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1069), .B1(new_n1053), .B2(new_n1035), .ZN(new_n1122));
  INV_X1    g697(.A(G1976), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT52), .B1(G288), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1122), .A2(KEYINPUT117), .A3(new_n1119), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1124), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1095), .B1(KEYINPUT45), .B2(new_n1097), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n720), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1050), .B1(new_n1097), .B2(new_n1054), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT50), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n797), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1069), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(G303), .A2(G8), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1136), .B(KEYINPUT55), .Z(new_n1137));
  OAI211_X1 g712(.A(new_n1121), .B(new_n1129), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1131), .B(new_n1139), .C1(new_n1093), .C2(G2090), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(G8), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1055), .A2(new_n797), .A3(new_n1058), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1139), .B1(new_n1142), .B2(new_n1131), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1138), .B1(new_n1144), .B2(new_n1137), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1084), .A2(new_n1088), .A3(new_n1109), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n1147));
  AND4_X1   g722(.A1(G168), .A2(new_n1072), .A3(new_n1129), .A4(new_n1121), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1137), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1147), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1121), .A2(new_n1129), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1142), .A2(new_n1131), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT116), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1154), .A2(G8), .A3(new_n1137), .A4(new_n1140), .ZN(new_n1155));
  NOR2_X1   g730(.A1(G286), .A2(KEYINPUT63), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1072), .B(new_n1156), .C1(new_n1137), .C2(new_n1135), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1152), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(new_n1123), .A3(new_n928), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1069), .B(new_n1110), .C1(new_n1160), .C2(new_n1112), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1151), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1146), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1164));
  AOI211_X1 g739(.A(new_n1099), .B(G2078), .C1(new_n1038), .C2(new_n1036), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1095), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1100), .A2(G301), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT54), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1100), .B(G301), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1092), .A2(new_n1035), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1097), .A2(new_n1054), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n847), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1166), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(G171), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1177));
  OAI211_X1 g752(.A(KEYINPUT54), .B(new_n1169), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1178), .B(new_n1145), .C1(new_n1087), .C2(new_n1082), .ZN(new_n1179));
  XNOR2_X1  g754(.A(G299), .B(KEYINPUT57), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT120), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT57), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G299), .B(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(G1956), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1186));
  XNOR2_X1  g761(.A(KEYINPUT56), .B(G2072), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1095), .B(new_n1187), .C1(KEYINPUT45), .C2(new_n1097), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1188), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1181), .B(new_n1185), .C1(new_n1186), .C2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1191));
  INV_X1    g766(.A(G1956), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1193), .A2(new_n1188), .A3(new_n1183), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n625), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT119), .ZN(new_n1197));
  OR3_X1    g772(.A1(new_n1117), .A2(new_n1197), .A3(G2067), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1197), .B1(new_n1117), .B2(G2067), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(G1348), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1196), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1190), .B1(new_n1195), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1190), .A2(new_n1194), .A3(KEYINPUT61), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1201), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1196), .A2(KEYINPUT60), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1196), .A2(KEYINPUT60), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OAI211_X1 g784(.A(new_n1095), .B(new_n1042), .C1(KEYINPUT45), .C2(new_n1097), .ZN(new_n1210));
  XOR2_X1   g785(.A(KEYINPUT58), .B(G1341), .Z(new_n1211));
  NAND2_X1  g786(.A1(new_n1117), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n568), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT59), .ZN(new_n1214));
  OAI21_X1  g789(.A(KEYINPUT122), .B1(new_n1214), .B2(KEYINPUT121), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(KEYINPUT122), .B2(new_n1214), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1215), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1217), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g794(.A(KEYINPUT60), .B(new_n1196), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1220));
  AND4_X1   g795(.A1(new_n1204), .A2(new_n1209), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1193), .A2(new_n1188), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1222), .A2(new_n1180), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1223), .A2(new_n1224), .A3(new_n1194), .ZN(new_n1225));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1222), .A2(KEYINPUT123), .A3(new_n1180), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1203), .B1(new_n1221), .B2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g804(.A1(new_n1168), .A2(new_n1179), .A3(new_n1229), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1049), .B1(new_n1163), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g806(.A1(new_n1039), .A2(G1996), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1232), .B(KEYINPUT46), .ZN(new_n1233));
  INV_X1    g808(.A(new_n857), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1041), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1233), .B1(new_n1235), .B2(new_n1040), .ZN(new_n1236));
  XOR2_X1   g811(.A(new_n1236), .B(KEYINPUT47), .Z(new_n1237));
  NAND2_X1  g812(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1238));
  OAI22_X1  g813(.A1(new_n1238), .A2(new_n1044), .B1(G2067), .B2(new_n775), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1047), .A2(new_n1040), .ZN(new_n1240));
  NOR3_X1   g815(.A1(G290), .A2(new_n1039), .A3(G1986), .ZN(new_n1241));
  XOR2_X1   g816(.A(new_n1241), .B(KEYINPUT48), .Z(new_n1242));
  AOI22_X1  g817(.A1(new_n1040), .A2(new_n1239), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  AND2_X1   g818(.A1(new_n1237), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1231), .A2(new_n1244), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g820(.A1(G227), .A2(new_n460), .ZN(new_n1247));
  NOR3_X1   g821(.A1(G401), .A2(G229), .A3(new_n1247), .ZN(new_n1248));
  OAI211_X1 g822(.A(new_n925), .B(new_n1248), .C1(new_n1023), .C2(new_n1025), .ZN(G225));
  INV_X1    g823(.A(G225), .ZN(G308));
endmodule


