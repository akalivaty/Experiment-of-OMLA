//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1312, new_n1313, new_n1314, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1388, new_n1389,
    new_n1390;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n209), .B(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G179), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT66), .B(G1), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(KEYINPUT67), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G1), .ZN(new_n256));
  AND4_X1   g0056(.A1(KEYINPUT67), .A2(new_n251), .A3(new_n254), .A4(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(G238), .B(new_n247), .C1(new_n252), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n219), .A2(G1698), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n259), .B1(G226), .B2(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G97), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n213), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT65), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n253), .B(G274), .C1(G41), .C2(G45), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT74), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n247), .A2(KEYINPUT65), .A3(new_n251), .A4(new_n273), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n270), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n271), .B1(new_n270), .B2(new_n274), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n258), .B(new_n267), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n270), .A2(new_n274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n270), .A2(new_n271), .A3(new_n274), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n278), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n283), .A2(new_n258), .A3(new_n267), .A4(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n245), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT13), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n247), .B1(new_n262), .B2(new_n263), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n281), .B2(new_n282), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(new_n289), .B2(new_n258), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n277), .A2(KEYINPUT13), .ZN(new_n291));
  OAI21_X1  g0091(.A(G169), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n286), .B1(new_n292), .B2(KEYINPUT14), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n277), .B(KEYINPUT13), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT14), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n294), .A2(KEYINPUT76), .A3(new_n295), .A4(G169), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n295), .B(G169), .C1(new_n290), .C2(new_n291), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT76), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n293), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n254), .A2(new_n256), .A3(G13), .A4(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G68), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT12), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n213), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n214), .A2(G33), .ZN(new_n308));
  INV_X1    g0108(.A(G77), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n308), .A2(new_n309), .B1(new_n214), .B2(G68), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n202), .A2(G20), .A3(G33), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT11), .ZN(new_n313));
  INV_X1    g0113(.A(new_n307), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n254), .A2(new_n256), .A3(G20), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n305), .B(new_n313), .C1(new_n303), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n300), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(KEYINPUT8), .A2(G58), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT68), .B(G58), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n321), .B2(KEYINPUT8), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT79), .B1(new_n322), .B2(new_n315), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT68), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(G58), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n218), .A2(KEYINPUT68), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT8), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n319), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n327), .A2(KEYINPUT79), .A3(new_n315), .A4(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n301), .A2(new_n314), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n323), .A2(new_n331), .B1(new_n301), .B2(new_n322), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n260), .A2(new_n261), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(new_n214), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT3), .ZN(new_n336));
  INV_X1    g0136(.A(G33), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n214), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT7), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n335), .A2(new_n341), .A3(G68), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n210), .B1(new_n320), .B2(new_n303), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G20), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT78), .ZN(new_n345));
  NOR2_X1   g0145(.A1(G20), .A2(G33), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G159), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(KEYINPUT78), .A3(G159), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT16), .A4(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n352), .A2(new_n307), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n340), .A2(new_n334), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n333), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G68), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n343), .A2(G20), .B1(new_n349), .B2(new_n350), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n332), .B1(new_n353), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(G232), .B(new_n247), .C1(new_n252), .C2(new_n257), .ZN(new_n363));
  OR2_X1    g0163(.A1(G223), .A2(G1698), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G1698), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n364), .B(new_n366), .C1(new_n260), .C2(new_n261), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G87), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n266), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n363), .A2(new_n280), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(G223), .A2(G1698), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n365), .B2(G1698), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n338), .A2(new_n339), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(G33), .B2(G87), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT80), .B1(new_n375), .B2(new_n247), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT80), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n369), .A2(new_n377), .A3(new_n266), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT70), .B(G179), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n363), .A2(new_n280), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n371), .A2(G169), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT18), .B1(new_n362), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT17), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n322), .A2(new_n301), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n329), .A2(new_n330), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT79), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n327), .A2(new_n328), .ZN(new_n388));
  INV_X1    g0188(.A(new_n315), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n385), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n352), .A2(new_n307), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT16), .B1(new_n357), .B2(new_n358), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n377), .B1(new_n369), .B2(new_n266), .ZN(new_n395));
  AOI211_X1 g0195(.A(KEYINPUT80), .B(new_n247), .C1(new_n367), .C2(new_n368), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT81), .B(G190), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n363), .A2(new_n280), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n363), .A2(new_n280), .A3(new_n370), .ZN(new_n400));
  INV_X1    g0200(.A(G200), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n398), .A2(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n384), .B1(new_n394), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n379), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n395), .A2(new_n396), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G169), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n405), .A2(new_n399), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n394), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n397), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n376), .A2(new_n378), .A3(new_n410), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n371), .A2(G200), .B1(new_n411), .B2(new_n381), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n361), .A2(new_n307), .A3(new_n352), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT17), .A4(new_n391), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n383), .A2(new_n403), .A3(new_n409), .A4(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT67), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n254), .A2(new_n256), .ZN(new_n417));
  INV_X1    g0217(.A(new_n251), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n248), .A2(KEYINPUT67), .A3(new_n251), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n266), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G244), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(G232), .A2(G1698), .ZN(new_n424));
  INV_X1    g0224(.A(G1698), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G238), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n374), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n266), .C1(G107), .C2(new_n374), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n280), .ZN(new_n429));
  OAI21_X1  g0229(.A(G200), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT8), .B(G58), .Z(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n346), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G20), .A2(G77), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT71), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n432), .B(new_n433), .C1(new_n435), .C2(new_n308), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n307), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n301), .A2(G77), .ZN(new_n438));
  INV_X1    g0238(.A(new_n316), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(G77), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n422), .A2(G190), .A3(new_n280), .A4(new_n428), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n430), .A2(new_n437), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n406), .B1(new_n423), .B2(new_n429), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n437), .A2(new_n440), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n422), .A2(new_n280), .A3(new_n379), .A4(new_n428), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(KEYINPUT72), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT72), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n442), .B2(new_n446), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n415), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G190), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n279), .B2(new_n285), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n317), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n294), .A2(G200), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n425), .B1(new_n338), .B2(new_n339), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(G223), .B1(new_n333), .B2(G77), .ZN(new_n459));
  AOI21_X1  g0259(.A(G1698), .B1(new_n338), .B2(new_n339), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G222), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n462), .A2(new_n266), .B1(new_n270), .B2(new_n274), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n421), .A2(G226), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n465), .A2(G169), .ZN(new_n466));
  INV_X1    g0266(.A(new_n308), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n322), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n346), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n314), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n301), .A2(new_n202), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n439), .B2(new_n202), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT69), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(KEYINPUT69), .B(new_n471), .C1(new_n439), .C2(new_n202), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n465), .A2(new_n379), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n466), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n401), .B1(new_n463), .B2(new_n464), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(G190), .B2(new_n465), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT9), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  AOI211_X1 g0284(.A(KEYINPUT9), .B(new_n470), .C1(new_n474), .C2(new_n475), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT10), .B1(new_n481), .B2(KEYINPUT73), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n482), .B(new_n487), .C1(new_n484), .C2(new_n485), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n480), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND4_X1   g0291(.A1(new_n318), .A2(new_n451), .A3(new_n457), .A4(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n214), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT22), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT22), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n374), .A2(new_n495), .A3(new_n214), .A4(G87), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT23), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n214), .B2(G107), .ZN(new_n500));
  INV_X1    g0300(.A(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(KEYINPUT23), .A3(G20), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n467), .A2(G116), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n497), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n498), .B1(new_n497), .B2(new_n503), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n307), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n501), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT25), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n301), .B2(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n254), .A2(new_n256), .A3(G33), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n301), .A2(new_n314), .A3(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n507), .A2(new_n509), .B1(new_n511), .B2(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n254), .A2(new_n256), .A3(G45), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G41), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G264), .B(new_n247), .C1(new_n513), .C2(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(G1), .A2(G13), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n272), .B1(new_n519), .B2(new_n246), .ZN(new_n520));
  XNOR2_X1  g0320(.A(KEYINPUT5), .B(G41), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n248), .A3(new_n521), .A4(G45), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G250), .A2(G1698), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n221), .B2(G1698), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n374), .B1(G33), .B2(G294), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n518), .B(new_n522), .C1(new_n525), .C2(new_n247), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n401), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n221), .A2(G1698), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(G250), .B2(G1698), .ZN(new_n529));
  INV_X1    g0329(.A(G294), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n529), .A2(new_n333), .B1(new_n337), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n266), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(new_n452), .A3(new_n518), .A4(new_n522), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n506), .A2(new_n512), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n512), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n497), .A2(new_n503), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT24), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n497), .A2(new_n498), .A3(new_n503), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n536), .B1(new_n540), .B2(new_n307), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n526), .A2(new_n406), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n532), .A2(new_n245), .A3(new_n518), .A4(new_n522), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n535), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G270), .B(new_n247), .C1(new_n513), .C2(new_n517), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n546), .A2(new_n522), .ZN(new_n547));
  OAI211_X1 g0347(.A(G257), .B(new_n425), .C1(new_n260), .C2(new_n261), .ZN(new_n548));
  OAI211_X1 g0348(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n549));
  XNOR2_X1  g0349(.A(KEYINPUT91), .B(G303), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n548), .B(new_n549), .C1(new_n374), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n266), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G116), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n302), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n301), .A2(new_n314), .A3(new_n510), .A4(G116), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n306), .A2(new_n213), .B1(G20), .B2(new_n554), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n558), .B(new_n214), .C1(G33), .C2(new_n220), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n557), .A2(KEYINPUT20), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT20), .B1(new_n557), .B2(new_n559), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n555), .B(new_n556), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n553), .A2(G169), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT92), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n551), .A2(new_n266), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n546), .A2(new_n522), .ZN(new_n568));
  OAI21_X1  g0368(.A(G200), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n562), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n547), .A2(new_n397), .A3(new_n552), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n562), .A2(G179), .A3(new_n552), .A4(new_n547), .ZN(new_n573));
  INV_X1    g0373(.A(new_n565), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n553), .A2(G169), .A3(new_n562), .A4(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n566), .A2(new_n572), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n545), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n214), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT88), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT88), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n581), .A3(new_n214), .ZN(new_n582));
  NOR3_X1   g0382(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n214), .B(G68), .C1(new_n260), .C2(new_n261), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n308), .B2(new_n220), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(new_n307), .B1(new_n302), .B2(new_n435), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT89), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT71), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n434), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n511), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n578), .A2(new_n581), .A3(new_n214), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n581), .B1(new_n578), .B2(new_n214), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n596), .A2(new_n597), .A3(new_n583), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n586), .A2(new_n588), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n307), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n435), .A2(new_n302), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n594), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT89), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G116), .ZN(new_n605));
  INV_X1    g0405(.A(G244), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G1698), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(G238), .B2(G1698), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n605), .B1(new_n608), .B2(new_n333), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n247), .A2(G250), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n609), .A2(new_n266), .B1(new_n513), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(G274), .B1(new_n265), .B2(new_n213), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT87), .B1(new_n513), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT87), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n520), .A2(new_n614), .A3(new_n248), .A4(G45), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(G169), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n611), .A2(new_n616), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n379), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n611), .A2(G190), .A3(new_n616), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT90), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n611), .A2(KEYINPUT90), .A3(G190), .A4(new_n616), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n511), .A2(G87), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n600), .A2(new_n601), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n401), .B1(new_n611), .B2(new_n616), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n604), .A2(new_n619), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(G244), .B(new_n425), .C1(new_n260), .C2(new_n261), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT4), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n606), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n374), .A2(new_n425), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n558), .A3(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(G250), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT84), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n374), .A2(new_n638), .A3(G250), .A4(G1698), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n266), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(G257), .B(new_n247), .C1(new_n513), .C2(new_n517), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n522), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT6), .ZN(new_n646));
  AND2_X1   g0446(.A1(G97), .A2(G107), .ZN(new_n647));
  NOR2_X1   g0447(.A1(G97), .A2(G107), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n501), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(G97), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT82), .ZN(new_n651));
  NAND2_X1  g0451(.A1(KEYINPUT6), .A2(G97), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(G107), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n346), .A2(G77), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n501), .B1(new_n354), .B2(new_n355), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n307), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n302), .A2(KEYINPUT83), .A3(new_n220), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT83), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n301), .B2(G97), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n660), .A2(new_n662), .B1(new_n511), .B2(G97), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n645), .A2(new_n406), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n558), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n460), .B2(new_n633), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n632), .A3(new_n637), .A4(new_n639), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n643), .B1(new_n667), .B2(new_n266), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT86), .B1(new_n668), .B2(new_n379), .ZN(new_n669));
  AND4_X1   g0469(.A1(KEYINPUT86), .A2(new_n641), .A3(new_n379), .A4(new_n644), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n645), .A2(KEYINPUT85), .A3(G200), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT85), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n668), .B2(new_n401), .ZN(new_n674));
  INV_X1    g0474(.A(new_n658), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n654), .A2(G20), .B1(G77), .B2(new_n346), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n314), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n660), .A2(new_n662), .ZN(new_n678));
  INV_X1    g0478(.A(new_n511), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n220), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n668), .A2(G190), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n672), .A2(new_n674), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n671), .A2(new_n683), .ZN(new_n684));
  AND4_X1   g0484(.A1(new_n492), .A2(new_n577), .A3(new_n629), .A4(new_n684), .ZN(G372));
  AND3_X1   g0485(.A1(new_n394), .A2(new_n407), .A3(new_n408), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n408), .B1(new_n394), .B2(new_n407), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n446), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n300), .B2(new_n317), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n403), .A2(new_n414), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n457), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n688), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT96), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n489), .A2(new_n490), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT96), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n696), .B(new_n688), .C1(new_n690), .C2(new_n692), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(new_n479), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n611), .A2(new_n616), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n406), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n701), .A2(KEYINPUT93), .B1(new_n618), .B2(new_n379), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n617), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n604), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n617), .A2(new_n703), .B1(new_n700), .B2(new_n404), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n617), .A2(new_n703), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(new_n604), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n671), .A2(new_n535), .A3(new_n683), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n566), .A2(new_n573), .A3(new_n575), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n544), .B1(new_n506), .B2(new_n512), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n600), .A2(new_n601), .A3(new_n625), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n718), .B(KEYINPUT94), .C1(new_n401), .C2(new_n618), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT94), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n626), .B2(new_n627), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n624), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n705), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n712), .B1(new_n717), .B2(new_n724), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n677), .A2(new_n680), .B1(new_n668), .B2(G169), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT86), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n645), .B2(new_n404), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n668), .A2(KEYINPUT86), .A3(new_n379), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n705), .A3(new_n722), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT26), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n629), .A2(new_n730), .A3(KEYINPUT26), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n725), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n492), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n699), .A2(new_n737), .ZN(G369));
  INV_X1    g0538(.A(KEYINPUT98), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n214), .A2(G13), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n248), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n741), .A2(KEYINPUT27), .ZN(new_n742));
  OAI21_X1  g0542(.A(G213), .B1(new_n741), .B2(KEYINPUT27), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(KEYINPUT97), .B(G343), .Z(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n541), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n545), .B1(new_n739), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n739), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n714), .A2(new_n748), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n715), .A2(new_n748), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n506), .A2(new_n512), .ZN(new_n758));
  INV_X1    g0558(.A(new_n544), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n751), .B1(new_n760), .B2(new_n748), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n748), .A2(new_n570), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n714), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n576), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G330), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n757), .A2(new_n767), .ZN(G399));
  NOR2_X1   g0568(.A1(new_n584), .A2(G116), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n207), .A2(new_n249), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(new_n770), .A3(G1), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n211), .B2(new_n770), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT28), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n684), .A2(new_n577), .A3(new_n629), .A4(new_n748), .ZN(new_n774));
  AND3_X1   g0574(.A1(new_n700), .A2(new_n379), .A3(new_n526), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT100), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n775), .A2(new_n776), .A3(new_n553), .A4(new_n645), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n553), .A2(new_n700), .A3(new_n379), .A4(new_n526), .ZN(new_n778));
  OAI21_X1  g0578(.A(KEYINPUT100), .B1(new_n778), .B2(new_n668), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n611), .A2(new_n518), .A3(new_n532), .A4(new_n616), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n567), .A2(new_n245), .A3(new_n568), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n782), .A2(new_n783), .A3(KEYINPUT30), .A4(new_n668), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n547), .A2(G179), .A3(new_n552), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n645), .A2(new_n785), .A3(new_n781), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT99), .B(KEYINPUT30), .Z(new_n787));
  OAI21_X1  g0587(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n747), .B1(new_n780), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT31), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n778), .A2(new_n668), .ZN(new_n792));
  OAI211_X1 g0592(.A(KEYINPUT31), .B(new_n747), .C1(new_n788), .C2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n774), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G330), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT101), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n794), .A2(KEYINPUT101), .A3(G330), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n747), .B1(new_n725), .B2(new_n735), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT29), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n710), .B1(new_n709), .B2(new_n604), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n575), .A2(new_n573), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n760), .A2(new_n805), .A3(new_n566), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n806), .A2(new_n535), .A3(new_n671), .A4(new_n683), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n804), .B1(new_n807), .B2(new_n723), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n591), .B1(new_n590), .B2(new_n594), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n602), .A2(KEYINPUT89), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n619), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n624), .A2(new_n628), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n732), .B1(new_n813), .B2(new_n671), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n730), .A2(new_n705), .A3(new_n722), .A4(KEYINPUT26), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(KEYINPUT29), .B(new_n748), .C1(new_n808), .C2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n799), .B1(new_n801), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n773), .B1(new_n818), .B2(G1), .ZN(G364));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n213), .B1(G20), .B2(new_n406), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT103), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n333), .A2(new_n207), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n240), .A2(new_n250), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT102), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n827), .B(new_n829), .C1(new_n250), .C2(new_n212), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n374), .A2(new_n207), .ZN(new_n831));
  INV_X1    g0631(.A(G355), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n831), .A2(new_n832), .B1(G116), .B2(new_n207), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n826), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n253), .B1(new_n740), .B2(G45), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n770), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n379), .A2(new_n214), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n401), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(G190), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n840), .A2(G200), .A3(new_n397), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n842), .A2(G77), .B1(new_n844), .B2(G50), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n840), .A2(new_n452), .A3(G200), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n841), .A2(new_n410), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n845), .B1(new_n303), .B2(new_n846), .C1(new_n320), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(G179), .A2(G200), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n214), .B1(new_n850), .B2(G190), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n220), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n850), .A2(G20), .A3(new_n452), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(new_n348), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n852), .B1(new_n855), .B2(KEYINPUT32), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n214), .A2(G179), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(G190), .A3(G200), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT32), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G87), .A2(new_n859), .B1(new_n854), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n857), .A2(new_n452), .A3(G200), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n501), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(new_n333), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n856), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(G283), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n853), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n374), .B(new_n867), .C1(G329), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n851), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n859), .A2(G303), .B1(new_n870), .B2(G294), .ZN(new_n871));
  XNOR2_X1  g0671(.A(KEYINPUT104), .B(G326), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n869), .B(new_n871), .C1(new_n843), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n847), .A2(G322), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n842), .A2(G311), .ZN(new_n875));
  XOR2_X1   g0675(.A(KEYINPUT33), .B(G317), .Z(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n875), .C1(new_n846), .C2(new_n876), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n849), .A2(new_n865), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n839), .B1(new_n823), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n822), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n879), .B1(new_n764), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n766), .A2(new_n838), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(G330), .B2(new_n764), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(G396));
  INV_X1    g0685(.A(new_n838), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n823), .A2(new_n820), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n309), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n444), .A2(new_n747), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n442), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n446), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n689), .A2(new_n748), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(G132), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n374), .B1(new_n853), .B2(new_n895), .C1(new_n862), .C2(new_n303), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n858), .A2(new_n202), .B1(new_n851), .B2(new_n320), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n847), .A2(G143), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n844), .A2(G137), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(G150), .ZN(new_n901));
  INV_X1    g0701(.A(new_n842), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n900), .B1(new_n901), .B2(new_n846), .C1(new_n348), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(KEYINPUT106), .B(KEYINPUT34), .Z(new_n905));
  AOI211_X1 g0705(.A(new_n896), .B(new_n897), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n902), .A2(new_n554), .B1(new_n866), .B2(new_n846), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n908), .A2(KEYINPUT105), .ZN(new_n909));
  INV_X1    g0709(.A(new_n862), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(G87), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(G107), .B2(new_n859), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n374), .B(new_n852), .C1(G311), .C2(new_n868), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(G303), .B2(new_n844), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n530), .B2(new_n848), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(KEYINPUT105), .B2(new_n908), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n906), .A2(new_n907), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n823), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n888), .B1(new_n821), .B2(new_n894), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n442), .A2(new_n446), .A3(new_n748), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n813), .A2(new_n732), .A3(new_n671), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n732), .B2(new_n731), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n922), .B1(new_n924), .B2(new_n808), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n800), .B2(new_n894), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n886), .B1(new_n927), .B2(new_n799), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n797), .B2(new_n798), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n920), .B1(new_n928), .B2(new_n929), .ZN(G384));
  OR2_X1    g0730(.A1(new_n654), .A2(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n654), .A2(KEYINPUT35), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(G116), .A3(new_n215), .A4(new_n932), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT36), .Z(new_n934));
  OAI211_X1 g0734(.A(new_n212), .B(G77), .C1(new_n303), .C2(new_n320), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n202), .A2(G68), .ZN(new_n936));
  AOI211_X1 g0736(.A(G13), .B(new_n248), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n492), .B(new_n817), .C1(new_n800), .C2(KEYINPUT29), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n699), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n925), .A2(new_n892), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT38), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT16), .B1(new_n358), .B2(new_n342), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n391), .B1(new_n392), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n744), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n691), .B2(new_n688), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n412), .A2(new_n413), .A3(new_n391), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n394), .A2(new_n407), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT37), .B1(new_n394), .B2(new_n744), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n944), .A2(new_n407), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n951), .A3(new_n945), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n949), .A2(new_n950), .B1(new_n952), .B2(KEYINPUT37), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n942), .B1(new_n946), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(KEYINPUT37), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(new_n947), .A3(new_n948), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n945), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n415), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT38), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n317), .A2(new_n747), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n318), .A2(new_n457), .A3(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n317), .B(new_n747), .C1(new_n300), .C2(new_n456), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n941), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT39), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n956), .A2(KEYINPUT107), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n394), .A2(new_n744), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n947), .A2(new_n948), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(KEYINPUT37), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT107), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n950), .A2(new_n947), .A3(new_n972), .A4(new_n948), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n968), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n415), .A2(new_n394), .A3(new_n744), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT38), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT38), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n967), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n300), .A2(new_n317), .A3(new_n748), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n954), .A2(KEYINPUT39), .A3(new_n960), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n745), .B1(new_n686), .B2(new_n687), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n966), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n940), .B(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n782), .A2(new_n783), .A3(new_n668), .ZN(new_n986));
  INV_X1    g0786(.A(new_n787), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n988), .A2(new_n777), .A3(new_n779), .A4(new_n784), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(KEYINPUT31), .A3(new_n747), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT31), .B1(new_n989), .B2(new_n747), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n893), .B1(new_n993), .B2(new_n774), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(new_n961), .A3(new_n965), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT40), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n965), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT40), .B1(new_n976), .B2(new_n977), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n774), .A2(new_n791), .A3(new_n990), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n492), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1003), .A2(G330), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n985), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n248), .B2(new_n740), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n985), .A2(new_n1005), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n938), .B1(new_n1007), .B2(new_n1008), .ZN(G367));
  OAI21_X1  g0809(.A(new_n684), .B1(new_n681), .B2(new_n748), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n730), .A2(new_n747), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n754), .A2(new_n755), .A3(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT45), .Z(new_n1014));
  INV_X1    g0814(.A(new_n1012), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT44), .B1(new_n756), .B2(new_n1015), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n756), .A2(KEYINPUT44), .A3(new_n1015), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n767), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n752), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n754), .B1(new_n761), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(new_n766), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n818), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n818), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n770), .B(KEYINPUT41), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n836), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT108), .B1(new_n754), .B2(new_n1015), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT108), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n753), .A2(new_n1030), .A3(new_n1012), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT42), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1010), .A2(new_n760), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n747), .B1(new_n1034), .B2(new_n671), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n1032), .B2(KEYINPUT42), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n748), .A2(new_n718), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n723), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n712), .B2(new_n1038), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT43), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1037), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1033), .A2(new_n1036), .A3(new_n1041), .A4(new_n1040), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n767), .A2(new_n1015), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1040), .A2(new_n822), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n236), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n826), .B1(new_n207), .B2(new_n435), .C1(new_n1051), .C2(new_n827), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n851), .A2(new_n303), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n910), .A2(G77), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n374), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(new_n847), .C2(G150), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT111), .ZN(new_n1057));
  INV_X1    g0857(.A(G137), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n858), .A2(new_n320), .B1(new_n1058), .B2(new_n853), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n842), .A2(G50), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n846), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1062), .A2(G159), .B1(new_n844), .B2(G143), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1059), .A2(KEYINPUT111), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1056), .A2(new_n1061), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n842), .A2(G283), .B1(G107), .B2(new_n870), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT109), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT109), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1062), .A2(G294), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n374), .B1(new_n868), .B2(G317), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n220), .B2(new_n862), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n859), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT46), .B1(new_n859), .B2(G116), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n550), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1076), .A2(new_n847), .B1(new_n844), .B2(G311), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT110), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1065), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT47), .Z(new_n1080));
  OAI211_X1 g0880(.A(new_n838), .B(new_n1052), .C1(new_n1080), .C2(new_n919), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1028), .A2(new_n1049), .B1(new_n1050), .B2(new_n1081), .ZN(G387));
  OR2_X1    g0882(.A1(new_n761), .A2(new_n880), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n769), .A2(new_n831), .B1(G107), .B2(new_n207), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n233), .A2(G45), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n769), .ZN(new_n1086));
  AOI211_X1 g0886(.A(G45), .B(new_n1086), .C1(G68), .C2(G77), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n431), .A2(new_n202), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT50), .Z(new_n1089));
  AOI21_X1  g0889(.A(new_n827), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1084), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n838), .B1(new_n1091), .B2(new_n825), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT112), .Z(new_n1093));
  NOR2_X1   g0893(.A1(new_n858), .A2(new_n309), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n374), .B1(new_n853), .B2(new_n901), .C1(new_n862), .C2(new_n220), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n593), .C2(new_n870), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n842), .A2(G68), .B1(new_n847), .B2(G50), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1062), .A2(new_n322), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n844), .A2(G159), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G317), .A2(new_n847), .B1(new_n1062), .B2(G311), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT114), .B(G322), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1101), .B1(new_n550), .B2(new_n902), .C1(new_n843), .C2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT48), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n858), .A2(new_n530), .B1(new_n851), .B2(new_n866), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT113), .Z(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(KEYINPUT49), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n333), .B1(new_n872), .B2(new_n853), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G116), .B2(new_n910), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT49), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1100), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1093), .B1(new_n1114), .B2(new_n823), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1023), .A2(new_n836), .B1(new_n1083), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1024), .A2(new_n837), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1023), .A2(new_n818), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(G393));
  XNOR2_X1  g0919(.A(new_n1018), .B(new_n767), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(new_n818), .A3(new_n1023), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n837), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1015), .A2(new_n822), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n826), .B1(new_n220), .B2(new_n207), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n243), .A2(new_n827), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n838), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n858), .A2(new_n866), .B1(new_n851), .B2(new_n554), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n333), .B1(new_n1102), .B2(new_n853), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1128), .A2(new_n863), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n902), .B2(new_n530), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G311), .A2(new_n847), .B1(new_n844), .B2(G317), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT52), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(new_n1076), .C2(new_n1062), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(KEYINPUT116), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(KEYINPUT116), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n333), .B(new_n911), .C1(G143), .C2(new_n868), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n303), .B2(new_n858), .C1(new_n309), .C2(new_n851), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n431), .B2(new_n842), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G159), .A2(new_n847), .B1(new_n844), .B2(G150), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1139), .B(new_n1142), .C1(new_n202), .C2(new_n846), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1135), .A2(new_n1136), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1127), .B1(new_n1144), .B2(new_n823), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1120), .A2(new_n836), .B1(new_n1124), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1123), .A2(new_n1146), .ZN(G390));
  AND3_X1   g0947(.A1(new_n794), .A2(KEYINPUT101), .A3(G330), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT101), .B1(new_n794), .B2(G330), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n894), .B(new_n965), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n748), .B(new_n891), .C1(new_n808), .C2(new_n816), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n892), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n963), .A2(new_n964), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1001), .A2(G330), .A3(new_n894), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1150), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n894), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n1154), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n941), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n492), .A2(G330), .A3(new_n1001), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n698), .A2(new_n939), .A3(new_n479), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n921), .B1(new_n725), .B2(new_n735), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n892), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n965), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1169), .A2(new_n979), .B1(new_n978), .B2(new_n981), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n979), .B1(new_n976), .B2(new_n977), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n1152), .B2(new_n965), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1158), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n925), .A2(new_n892), .B1(new_n963), .B2(new_n964), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n974), .A2(new_n975), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n942), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT39), .B1(new_n1176), .B2(new_n960), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n954), .A2(KEYINPUT39), .A3(new_n960), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1174), .A2(new_n980), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1152), .A2(new_n965), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1171), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1179), .A2(new_n1182), .A3(new_n1150), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1173), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1166), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1162), .A2(new_n1183), .A3(new_n1173), .A4(new_n1165), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n837), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n820), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n887), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n838), .B1(new_n322), .B2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1062), .A2(G137), .B1(new_n844), .B2(G128), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1191), .B1(new_n895), .B2(new_n848), .C1(new_n902), .C2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n858), .A2(new_n901), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1195));
  XNOR2_X1  g0995(.A(new_n1194), .B(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(G125), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n374), .B1(new_n853), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G50), .B2(new_n910), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1196), .B(new_n1199), .C1(new_n348), .C2(new_n851), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1062), .A2(G107), .B1(new_n844), .B2(G283), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n220), .B2(new_n902), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n862), .A2(new_n303), .B1(new_n530), .B2(new_n853), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT118), .Z(new_n1204));
  NOR2_X1   g1004(.A1(new_n851), .A2(new_n309), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n374), .B(new_n1205), .C1(G87), .C2(new_n859), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n554), .C2(new_n848), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n1193), .A2(new_n1200), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1190), .B1(new_n1208), .B2(new_n823), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1188), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1184), .B2(new_n835), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1187), .A2(new_n1212), .ZN(G378));
  NAND2_X1  g1013(.A1(new_n695), .A2(new_n479), .ZN(new_n1214));
  XOR2_X1   g1014(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1215), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n491), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n477), .A2(new_n744), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT121), .Z(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1216), .A2(new_n1221), .A3(new_n1218), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1001), .A2(new_n894), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n963), .B2(new_n964), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT40), .B1(new_n1227), .B2(new_n961), .ZN(new_n1228));
  OAI21_X1  g1028(.A(G330), .B1(new_n998), .B2(new_n999), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1225), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(G330), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n996), .B1(new_n1176), .B2(new_n960), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n997), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1230), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n984), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n984), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1230), .A2(new_n1238), .A3(new_n1235), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1225), .A2(new_n820), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n838), .B1(G50), .B2(new_n1189), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n858), .A2(new_n1192), .B1(new_n851), .B2(new_n901), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n842), .A2(G137), .B1(new_n847), .B2(G128), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1197), .B2(new_n843), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(G132), .C2(new_n1062), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT59), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1249));
  OR2_X1    g1049(.A1(KEYINPUT120), .A2(G124), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(KEYINPUT120), .A2(G124), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n868), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(new_n337), .A3(new_n249), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G159), .B2(new_n910), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1248), .A2(new_n1249), .A3(new_n1254), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n848), .A2(new_n501), .B1(new_n220), .B2(new_n846), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n333), .B(new_n249), .C1(new_n853), .C2(new_n866), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n862), .A2(new_n320), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1094), .A2(new_n1257), .A3(new_n1258), .A4(new_n1053), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n435), .B2(new_n902), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1256), .B(new_n1260), .C1(G116), .C2(new_n844), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1261), .A2(KEYINPUT58), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(KEYINPUT58), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G50), .B1(new_n337), .B2(new_n249), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n374), .B2(G41), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT119), .Z(new_n1266));
  NAND4_X1  g1066(.A1(new_n1255), .A2(new_n1262), .A3(new_n1263), .A4(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1242), .B1(new_n1267), .B2(new_n823), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1240), .A2(new_n836), .B1(new_n1241), .B2(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1230), .A2(new_n1238), .A3(new_n1235), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1238), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT57), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1173), .A2(new_n1183), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1164), .B1(new_n1273), .B2(new_n1162), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n837), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n994), .A2(new_n965), .A3(G330), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n893), .B1(new_n797), .B2(new_n798), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1276), .B1(new_n1277), .B2(new_n965), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1278), .A2(new_n941), .B1(new_n1279), .B2(new_n1150), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1165), .B1(new_n1184), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1269), .B1(new_n1275), .B2(new_n1282), .ZN(G375));
  OAI211_X1 g1083(.A(new_n1164), .B(new_n1157), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1166), .A2(new_n1027), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1154), .A2(new_n820), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n838), .B1(G68), .B2(new_n1189), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1062), .A2(G116), .B1(new_n844), .B2(G294), .ZN(new_n1288));
  OAI221_X1 g1088(.A(new_n1288), .B1(new_n501), .B2(new_n902), .C1(new_n866), .C2(new_n848), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n374), .B1(new_n868), .B2(G303), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1054), .A2(new_n1290), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1291), .B1(new_n220), .B2(new_n858), .C1(new_n435), .C2(new_n851), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n842), .A2(G150), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1258), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n333), .B1(new_n868), .B2(G128), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n859), .A2(G159), .B1(new_n870), .B2(G50), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n844), .A2(G132), .ZN(new_n1298));
  OAI221_X1 g1098(.A(new_n1298), .B1(new_n846), .B2(new_n1192), .C1(new_n848), .C2(new_n1058), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n1289), .A2(new_n1292), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1287), .B1(new_n1300), .B2(new_n823), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1162), .A2(new_n836), .B1(new_n1286), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1285), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(KEYINPUT122), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(G381));
  NOR4_X1   g1105(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1306));
  INV_X1    g1106(.A(G387), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n770), .B1(new_n1166), .B2(new_n1184), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1211), .B1(new_n1308), .B2(new_n1186), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1306), .A2(new_n1307), .A3(new_n1309), .A4(new_n1304), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1310), .A2(G375), .ZN(G407));
  NAND2_X1  g1111(.A1(new_n746), .A2(G213), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G407), .B(G213), .C1(G375), .C2(new_n1314), .ZN(G409));
  OAI211_X1 g1115(.A(G378), .B(new_n1269), .C1(new_n1275), .C2(new_n1282), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1240), .A2(new_n1027), .A3(new_n1281), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n836), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1241), .A2(new_n1268), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1309), .B1(new_n1317), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1316), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n770), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT60), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1284), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1278), .A2(new_n941), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1326), .A2(KEYINPUT60), .A3(new_n1164), .A4(new_n1157), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1323), .A2(new_n1325), .A3(new_n1327), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1328), .A2(G384), .A3(new_n1302), .ZN(new_n1329));
  AOI21_X1  g1129(.A(G384), .B1(new_n1328), .B2(new_n1302), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1322), .A2(new_n1312), .A3(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT123), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1313), .B1(new_n1316), .B2(new_n1321), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(KEYINPUT123), .A3(new_n1331), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT62), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1322), .A2(new_n1312), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT124), .ZN(new_n1339));
  INV_X1    g1139(.A(G2897), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1312), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1329), .A2(new_n1330), .A3(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1328), .A2(new_n1302), .ZN(new_n1344));
  INV_X1    g1144(.A(G384), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1328), .A2(G384), .A3(new_n1302), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1341), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1339), .B1(new_n1343), .B2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1342), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1346), .A2(new_n1347), .A3(new_n1341), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1350), .A2(new_n1351), .A3(KEYINPUT124), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1338), .A2(new_n1349), .A3(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1332), .A2(KEYINPUT62), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT61), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1353), .A2(new_n1354), .A3(new_n1355), .ZN(new_n1356));
  OAI21_X1  g1156(.A(KEYINPUT127), .B1(new_n1337), .B2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT62), .ZN(new_n1358));
  AND4_X1   g1158(.A1(KEYINPUT123), .A2(new_n1322), .A3(new_n1312), .A4(new_n1331), .ZN(new_n1359));
  AOI21_X1  g1159(.A(KEYINPUT123), .B1(new_n1335), .B2(new_n1331), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1358), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT127), .ZN(new_n1362));
  AOI21_X1  g1162(.A(KEYINPUT124), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1363), .A2(new_n1335), .ZN(new_n1364));
  AOI21_X1  g1164(.A(KEYINPUT61), .B1(new_n1364), .B2(new_n1352), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1361), .A2(new_n1362), .A3(new_n1365), .A4(new_n1354), .ZN(new_n1366));
  XNOR2_X1  g1166(.A(G393), .B(new_n884), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(G387), .A2(KEYINPUT126), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1367), .B1(new_n1368), .B2(G390), .ZN(new_n1369));
  INV_X1    g1169(.A(G390), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(G387), .A2(KEYINPUT126), .A3(new_n1370), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT125), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1370), .A2(new_n1372), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1372), .B1(new_n1123), .B2(new_n1146), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1374), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1307), .A2(new_n1373), .A3(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1367), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1377), .B1(G387), .B2(new_n1374), .ZN(new_n1378));
  AOI22_X1  g1178(.A1(new_n1369), .A2(new_n1371), .B1(new_n1376), .B2(new_n1378), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1357), .A2(new_n1366), .A3(new_n1379), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1369), .A2(new_n1371), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1376), .A2(new_n1378), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1381), .A2(new_n1382), .ZN(new_n1383));
  OR3_X1    g1183(.A1(new_n1359), .A2(new_n1360), .A3(KEYINPUT63), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1335), .A2(KEYINPUT63), .A3(new_n1331), .ZN(new_n1385));
  NAND4_X1  g1185(.A1(new_n1383), .A2(new_n1384), .A3(new_n1365), .A4(new_n1385), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1380), .A2(new_n1386), .ZN(G405));
  NAND2_X1  g1187(.A1(G375), .A2(new_n1309), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1388), .A2(new_n1316), .ZN(new_n1389));
  XNOR2_X1  g1189(.A(new_n1389), .B(new_n1331), .ZN(new_n1390));
  XNOR2_X1  g1190(.A(new_n1379), .B(new_n1390), .ZN(G402));
endmodule


