//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1069, new_n1070, new_n1071, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(new_n190), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT11), .B1(new_n194), .B2(G137), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(G137), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n200), .B1(new_n199), .B2(new_n201), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT79), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  AOI21_X1  g022(.A(G104), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G107), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n210), .A2(KEYINPUT3), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n206), .A3(new_n208), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n216));
  AOI21_X1  g030(.A(G101), .B1(new_n210), .B2(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n212), .A2(new_n213), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n213), .B1(new_n212), .B2(new_n218), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(G128), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT66), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G143), .B(G146), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(G128), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n228), .B1(new_n233), .B2(new_n234), .ZN(new_n240));
  OR2_X1    g054(.A1(KEYINPUT67), .A2(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT67), .A2(G128), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n231), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT69), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n232), .A2(new_n238), .B1(new_n244), .B2(new_n231), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n221), .A2(KEYINPUT10), .A3(new_n247), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT10), .ZN(new_n252));
  OAI22_X1  g066(.A1(new_n236), .A2(G128), .B1(new_n223), .B2(new_n230), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n232), .B2(new_n238), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n212), .A2(new_n218), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n231), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n236), .A2(KEYINPUT0), .A3(G128), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n210), .A2(G107), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n215), .A2(new_n216), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G101), .ZN(new_n265));
  INV_X1    g079(.A(G101), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT3), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(G104), .B2(new_n205), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT79), .B(G107), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(new_n214), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n266), .B1(new_n270), .B2(new_n262), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n218), .A2(KEYINPUT4), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n261), .B(new_n265), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n256), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n204), .B1(new_n251), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n256), .A2(new_n273), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n239), .A2(new_n249), .A3(new_n245), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n249), .B1(new_n239), .B2(new_n245), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n219), .A2(new_n220), .A3(new_n252), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT81), .B1(new_n282), .B2(new_n204), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n251), .A2(new_n274), .A3(KEYINPUT81), .A4(new_n204), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n276), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(G110), .B(G140), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n288), .A2(G227), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n287), .B(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n251), .A2(new_n274), .A3(new_n204), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT81), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n290), .B1(new_n294), .B2(new_n284), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n248), .A2(new_n255), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT82), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n254), .A2(new_n255), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT82), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n248), .A2(new_n299), .A3(new_n255), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n199), .A2(new_n201), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G131), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT83), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT12), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n301), .B(new_n305), .C1(new_n307), .C2(KEYINPUT12), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n295), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(G902), .B1(new_n291), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n193), .B1(new_n313), .B2(new_n192), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n294), .A2(new_n284), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n311), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n290), .ZN(new_n317));
  INV_X1    g131(.A(new_n290), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT84), .B(new_n318), .C1(new_n283), .C2(new_n285), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n276), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n295), .A2(KEYINPUT84), .ZN(new_n321));
  OAI211_X1 g135(.A(G469), .B(new_n317), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n191), .B1(new_n314), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G475), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT18), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(new_n200), .ZN(new_n326));
  NOR2_X1   g140(.A1(G237), .A2(G953), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(G143), .A3(G214), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(G143), .B1(new_n327), .B2(G214), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G125), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G146), .ZN(new_n337));
  XNOR2_X1  g151(.A(G125), .B(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n227), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G237), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n288), .A3(G214), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n229), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n343), .B(new_n328), .C1(new_n325), .C2(new_n200), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n331), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT88), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n331), .A2(new_n340), .A3(new_n344), .A4(KEYINPUT88), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G113), .B(G122), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(new_n210), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n343), .A2(new_n328), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G131), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT17), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n343), .A2(new_n200), .A3(new_n328), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n338), .A2(KEYINPUT16), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n333), .A2(KEYINPUT16), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n227), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n352), .A2(KEYINPUT17), .A3(G131), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(G146), .A3(new_n358), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n356), .A2(new_n360), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n349), .A2(new_n351), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n351), .B1(new_n349), .B2(new_n363), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n324), .B1(new_n366), .B2(new_n190), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n338), .B(KEYINPUT19), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n227), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n353), .A2(new_n355), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n362), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n351), .B1(new_n349), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT89), .B1(new_n364), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(G475), .A2(G902), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n349), .A2(new_n351), .A3(new_n363), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT89), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n369), .A2(new_n362), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n377), .A2(new_n370), .B1(new_n347), .B2(new_n348), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n375), .B(new_n376), .C1(new_n378), .C2(new_n351), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT20), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(new_n374), .C1(new_n364), .C2(new_n372), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n367), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n385));
  INV_X1    g199(.A(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G116), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT14), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT92), .ZN(new_n390));
  INV_X1    g204(.A(G116), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G122), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n389), .A2(new_n392), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT92), .B1(new_n392), .B2(KEYINPUT14), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n393), .B(G107), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n241), .A2(G143), .A3(new_n242), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n229), .A2(G128), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n194), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n269), .A2(new_n387), .A3(new_n392), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(G134), .A3(new_n398), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n396), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT13), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G134), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n399), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n397), .A2(KEYINPUT13), .A3(G134), .A4(new_n398), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n206), .A2(new_n208), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n387), .A2(new_n392), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n401), .A2(new_n413), .A3(KEYINPUT90), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n411), .A2(new_n412), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n206), .A2(new_n208), .B1(new_n387), .B2(new_n392), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n410), .A2(KEYINPUT91), .A3(new_n414), .A4(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n406), .A2(G134), .B1(new_n398), .B2(new_n397), .ZN(new_n421));
  INV_X1    g235(.A(new_n409), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n418), .A2(new_n414), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n404), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n189), .A2(G217), .A3(new_n288), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n385), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n419), .A2(new_n425), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n403), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT94), .A3(new_n427), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n426), .A2(KEYINPUT93), .A3(new_n428), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT93), .B1(new_n426), .B2(new_n428), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n429), .B(new_n432), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  NOR2_X1   g250(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n440), .B(KEYINPUT96), .Z(new_n441));
  AND3_X1   g255(.A1(new_n435), .A2(new_n190), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n440), .A2(KEYINPUT96), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n435), .B2(new_n190), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n384), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G952), .ZN(new_n448));
  AOI211_X1 g262(.A(G953), .B(new_n448), .C1(G234), .C2(G237), .ZN(new_n449));
  INV_X1    g263(.A(G234), .ZN(new_n450));
  OAI211_X1 g264(.A(G902), .B(G953), .C1(new_n450), .C2(new_n341), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT97), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(G898), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G214), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n255), .A2(KEYINPUT80), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n212), .A2(new_n213), .A3(new_n218), .ZN(new_n460));
  INV_X1    g274(.A(G113), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT2), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT2), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G113), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G116), .B(G119), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT68), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(KEYINPUT5), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n391), .A2(KEYINPUT5), .A3(G119), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(new_n461), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n468), .A2(new_n470), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n459), .A2(new_n460), .A3(new_n474), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n465), .A2(new_n466), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n469), .B1(new_n465), .B2(new_n466), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n479), .B(new_n265), .C1(new_n271), .C2(new_n272), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT85), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n483), .A3(new_n480), .ZN(new_n484));
  XNOR2_X1  g298(.A(G110), .B(G122), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n480), .A3(new_n485), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT6), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n485), .B1(new_n481), .B2(KEYINPUT85), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT6), .A3(new_n484), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n259), .A2(new_n260), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G125), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n246), .B2(G125), .ZN(new_n495));
  INV_X1    g309(.A(G224), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G953), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n497), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n490), .A2(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n488), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n485), .B(KEYINPUT8), .Z(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n474), .B2(new_n255), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n473), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n468), .A2(new_n470), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n504), .B1(new_n509), .B2(new_n255), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n495), .A2(new_n501), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n499), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n190), .B1(new_n502), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT87), .B(new_n458), .C1(new_n500), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n498), .A2(new_n499), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n491), .A2(KEYINPUT6), .A3(new_n484), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n491), .A2(new_n484), .B1(KEYINPUT6), .B2(new_n488), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n513), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n458), .A2(KEYINPUT87), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n454), .B(new_n456), .C1(new_n514), .C2(new_n521), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n323), .A2(new_n447), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT22), .B(G137), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n187), .A2(new_n450), .A3(G953), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n524), .B(new_n525), .Z(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n360), .A2(new_n362), .ZN(new_n528));
  AND2_X1   g342(.A1(KEYINPUT67), .A2(G128), .ZN(new_n529));
  NOR2_X1   g343(.A1(KEYINPUT67), .A2(G128), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT23), .A3(G119), .ZN(new_n532));
  INV_X1    g346(.A(G128), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT23), .B1(new_n533), .B2(G119), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(G119), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G110), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(G119), .ZN(new_n539));
  INV_X1    g353(.A(new_n535), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT24), .B(G110), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n528), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT78), .ZN(new_n545));
  INV_X1    g359(.A(G119), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n243), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n541), .B1(new_n547), .B2(new_n535), .ZN(new_n548));
  INV_X1    g362(.A(G110), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n532), .A2(new_n549), .A3(new_n536), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n550), .A3(KEYINPUT77), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n362), .A2(new_n339), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT77), .B1(new_n548), .B2(new_n550), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n544), .B(new_n545), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT77), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n532), .A2(new_n536), .A3(new_n549), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n542), .B1(new_n539), .B2(new_n540), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n551), .A3(new_n552), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n545), .B1(new_n561), .B2(new_n544), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n527), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n544), .B1(new_n553), .B2(new_n554), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n526), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G217), .B1(new_n450), .B2(G902), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n190), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n565), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n564), .A2(KEYINPUT78), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n555), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(new_n573), .B2(new_n527), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT25), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n574), .A2(new_n575), .A3(G902), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT25), .B1(new_n566), .B2(new_n190), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n567), .B(KEYINPUT76), .Z(new_n579));
  OAI21_X1  g393(.A(new_n570), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT32), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT64), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n201), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n197), .A2(G134), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n194), .A2(KEYINPUT64), .A3(G137), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G131), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(new_n304), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n247), .A2(new_n588), .A3(new_n250), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n204), .A2(new_n493), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT30), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n479), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n587), .A2(new_n304), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n204), .A2(new_n493), .B1(new_n248), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n596), .B2(new_n591), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n327), .A2(G210), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT27), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT26), .B(G101), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n305), .A2(new_n261), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n479), .A2(KEYINPUT70), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT70), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n508), .A2(new_n606), .A3(new_n476), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n603), .B1(new_n608), .B2(new_n589), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n598), .A2(KEYINPUT71), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT71), .B1(new_n598), .B2(new_n609), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT31), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n598), .A2(new_n609), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT31), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n278), .A2(new_n279), .A3(new_n595), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT73), .B1(new_n616), .B2(new_n590), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT73), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n589), .A2(new_n618), .A3(new_n604), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n605), .A2(new_n607), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT28), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n608), .A2(new_n589), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT72), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n596), .A2(new_n626), .A3(new_n479), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n246), .A2(new_n588), .B1(new_n305), .B2(new_n261), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT72), .B1(new_n628), .B2(new_n594), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n625), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT28), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n612), .A2(new_n615), .B1(new_n632), .B2(new_n603), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT74), .B1(G472), .B2(G902), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(KEYINPUT74), .A2(G472), .A3(G902), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n581), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n631), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n589), .A2(new_n604), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n620), .B1(new_n640), .B2(KEYINPUT73), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT28), .B1(new_n641), .B2(new_n619), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n603), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT71), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n613), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n598), .A2(KEYINPUT71), .A3(new_n609), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n614), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n615), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n637), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(KEYINPUT32), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n638), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n603), .B1(new_n630), .B2(KEYINPUT28), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT75), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n624), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n624), .B2(new_n653), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT29), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n593), .A2(new_n597), .B1(new_n589), .B2(new_n608), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n657), .B1(new_n658), .B2(new_n602), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n625), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n621), .B1(new_n589), .B2(new_n604), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT28), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n603), .A2(new_n657), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n624), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n190), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n660), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n580), .B1(new_n652), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n523), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT98), .B(G101), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G3));
  OAI21_X1  g485(.A(new_n318), .B1(new_n283), .B2(new_n285), .ZN(new_n672));
  INV_X1    g486(.A(new_n311), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n275), .B1(new_n294), .B2(new_n284), .ZN(new_n674));
  OAI22_X1  g488(.A1(new_n672), .A2(new_n673), .B1(new_n674), .B2(new_n318), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n192), .A3(new_n190), .ZN(new_n676));
  INV_X1    g490(.A(new_n193), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n322), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n191), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(G472), .B1(new_n633), .B2(G902), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n649), .A2(new_n650), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n575), .B1(new_n574), .B2(G902), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n566), .A2(KEYINPUT25), .A3(new_n190), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n579), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n685), .A2(new_n686), .B1(new_n566), .B2(new_n569), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n681), .A2(new_n682), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT99), .B1(new_n680), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(G472), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n649), .B2(new_n190), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n612), .A2(new_n615), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n637), .B1(new_n692), .B2(new_n643), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n323), .A2(new_n694), .A3(new_n695), .A4(new_n687), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n457), .B1(new_n500), .B2(new_n513), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n518), .A2(new_n519), .A3(new_n458), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n455), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n381), .A2(new_n383), .ZN(new_n701));
  INV_X1    g515(.A(new_n367), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n454), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n190), .A2(G478), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT93), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n431), .B2(new_n427), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n426), .A2(KEYINPUT93), .A3(new_n428), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT33), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n429), .A4(new_n432), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT100), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n426), .B2(new_n428), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n426), .A2(new_n428), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n426), .A2(new_n712), .A3(new_n428), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT33), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n705), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT101), .B(G478), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n435), .B2(new_n190), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n703), .B(new_n704), .C1(new_n718), .C2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n697), .A2(new_n700), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT102), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT34), .B(G104), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G6));
  NAND2_X1  g539(.A1(new_n435), .A2(new_n190), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n443), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n435), .A2(new_n190), .A3(new_n441), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n373), .A2(new_n382), .A3(new_n379), .A4(new_n374), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n367), .B1(new_n381), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n727), .A2(new_n728), .A3(new_n704), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n700), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n689), .A2(new_n696), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT35), .B(G107), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G9));
  NAND2_X1  g549(.A1(new_n681), .A2(new_n682), .ZN(new_n736));
  OR3_X1    g550(.A1(new_n573), .A2(KEYINPUT36), .A3(new_n527), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n573), .B1(KEYINPUT36), .B2(new_n527), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n568), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n685), .B2(new_n686), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n523), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT37), .B(G110), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G12));
  NAND2_X1  g558(.A1(new_n624), .A2(new_n653), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n659), .B1(new_n745), .B2(KEYINPUT75), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n624), .A2(new_n653), .A3(new_n654), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n666), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n638), .B(new_n651), .C1(new_n690), .C2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(G900), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n449), .B1(new_n452), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT103), .Z(new_n752));
  NAND4_X1  g566(.A1(new_n727), .A2(new_n728), .A3(new_n730), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n740), .A2(new_n700), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n749), .A2(new_n323), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G128), .ZN(G30));
  NOR2_X1   g571(.A1(new_n610), .A2(new_n611), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n603), .B1(new_n661), .B2(new_n662), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(G902), .B1(new_n760), .B2(KEYINPUT104), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(KEYINPUT104), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(G472), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n652), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n514), .A2(KEYINPUT38), .A3(new_n521), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT38), .B1(new_n514), .B2(new_n521), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n740), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n703), .A2(new_n727), .A3(new_n728), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n769), .A2(new_n770), .A3(new_n456), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n764), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n752), .B(KEYINPUT39), .Z(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n191), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n678), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(KEYINPUT40), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n775), .A2(KEYINPUT40), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n772), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n229), .ZN(G45));
  OAI211_X1 g593(.A(new_n703), .B(new_n752), .C1(new_n718), .C2(new_n720), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n749), .A2(new_n323), .A3(new_n755), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G146), .ZN(G48));
  AOI22_X1  g597(.A1(new_n286), .A2(new_n290), .B1(new_n295), .B2(new_n311), .ZN(new_n784));
  OAI21_X1  g598(.A(G469), .B1(new_n784), .B2(G902), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n679), .A3(new_n676), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n700), .ZN(new_n787));
  INV_X1    g601(.A(new_n721), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n749), .A3(new_n687), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT41), .B(G113), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G15));
  AND3_X1   g605(.A1(new_n785), .A2(new_n679), .A3(new_n676), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n749), .A2(new_n687), .A3(new_n732), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G116), .ZN(G18));
  NOR3_X1   g608(.A1(new_n446), .A2(new_n740), .A3(new_n454), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n787), .A2(new_n749), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G119), .ZN(G21));
  INV_X1    g611(.A(KEYINPUT107), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n770), .A2(new_n700), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n792), .A2(new_n799), .A3(new_n704), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n640), .A2(new_n620), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n623), .B1(new_n801), .B2(new_n625), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT106), .B1(new_n642), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT106), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n624), .A2(new_n804), .A3(new_n663), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n805), .A3(new_n603), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n692), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n637), .B(KEYINPUT105), .Z(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n681), .B(new_n687), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n798), .B1(new_n800), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n442), .A2(new_n445), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n518), .A2(new_n519), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n456), .B1(new_n813), .B2(new_n457), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n812), .A2(new_n814), .A3(new_n703), .A4(new_n699), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n785), .A2(new_n679), .A3(new_n676), .A4(new_n704), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n809), .B1(new_n806), .B2(new_n692), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n691), .A2(new_n580), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(KEYINPUT107), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n811), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G122), .ZN(G24));
  NOR3_X1   g636(.A1(new_n691), .A2(new_n818), .A3(new_n740), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n787), .A2(new_n823), .A3(new_n781), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G125), .ZN(G27));
  INV_X1    g639(.A(KEYINPUT109), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n693), .B2(KEYINPUT32), .ZN(new_n827));
  OAI211_X1 g641(.A(KEYINPUT109), .B(new_n581), .C1(new_n633), .C2(new_n637), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n667), .A3(new_n651), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n191), .A2(new_n456), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n514), .A2(new_n521), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT108), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n320), .A2(new_n321), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n275), .B1(new_n295), .B2(KEYINPUT84), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT84), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n672), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT108), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(G469), .B(new_n317), .C1(new_n833), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n831), .B1(new_n838), .B2(new_n314), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n829), .A2(new_n839), .A3(new_n687), .A4(new_n781), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT42), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n780), .A2(KEYINPUT42), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n668), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(G131), .ZN(G33));
  INV_X1    g659(.A(KEYINPUT110), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n753), .B(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n668), .A2(new_n839), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G134), .ZN(G36));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n677), .A2(KEYINPUT46), .ZN(new_n851));
  OAI211_X1 g665(.A(KEYINPUT45), .B(new_n317), .C1(new_n833), .C2(new_n837), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT45), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n192), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n851), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n676), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n850), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n318), .B1(new_n315), .B2(new_n311), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n834), .B2(new_n836), .ZN(new_n860));
  OAI21_X1  g674(.A(G469), .B1(new_n860), .B2(KEYINPUT45), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n832), .B1(new_n320), .B2(new_n321), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT108), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n861), .B1(KEYINPUT45), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(KEYINPUT111), .B(new_n676), .C1(new_n865), .C2(new_n851), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT46), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n865), .B2(new_n193), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n858), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n774), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT112), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n514), .A2(new_n521), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n456), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n384), .B1(new_n718), .B2(new_n720), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n874), .A2(KEYINPUT43), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(KEYINPUT43), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n736), .A3(new_n769), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT44), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n881), .A2(new_n882), .B1(new_n878), .B2(new_n877), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n871), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(G137), .ZN(G39));
  INV_X1    g699(.A(KEYINPUT47), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n869), .A2(new_n886), .A3(new_n679), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n886), .B1(new_n869), .B2(new_n679), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n873), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n749), .A2(new_n890), .A3(new_n687), .A4(new_n780), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(G140), .ZN(G42));
  AOI21_X1  g707(.A(KEYINPUT114), .B1(new_n687), .B2(new_n830), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n764), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n768), .A2(new_n874), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n785), .A2(new_n676), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT49), .Z(new_n898));
  NAND3_X1  g712(.A1(new_n687), .A2(KEYINPUT114), .A3(new_n830), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n895), .A2(new_n896), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n652), .A2(new_n687), .A3(new_n763), .ZN(new_n901));
  INV_X1    g715(.A(new_n449), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n897), .A2(new_n831), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n720), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n711), .A2(new_n717), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n705), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n703), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(G952), .A3(new_n288), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n903), .A2(new_n875), .A3(new_n876), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n829), .A2(new_n687), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT48), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n449), .A2(new_n819), .A3(new_n875), .A4(new_n876), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n910), .B(new_n914), .C1(new_n787), .C2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n823), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n908), .A2(new_n703), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n905), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n456), .B1(new_n766), .B2(new_n767), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT119), .B1(new_n921), .B2(new_n786), .ZN(new_n922));
  INV_X1    g736(.A(new_n767), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n455), .B1(new_n923), .B2(new_n765), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n925), .A3(new_n792), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n927), .A2(KEYINPUT50), .A3(new_n915), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT50), .B1(new_n927), .B2(new_n915), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n920), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI22_X1  g744(.A1(new_n887), .A2(new_n888), .B1(new_n679), .B2(new_n897), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n915), .A2(new_n873), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT51), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI211_X1 g749(.A(KEYINPUT51), .B(new_n930), .C1(new_n931), .C2(new_n932), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n916), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n789), .A2(new_n793), .A3(new_n796), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n703), .B(new_n906), .C1(new_n907), .C2(new_n705), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n522), .A2(new_n446), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n689), .A2(new_n696), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n523), .B1(new_n668), .B2(new_n741), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(new_n821), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n680), .B1(new_n652), .B2(new_n667), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n730), .B(new_n752), .C1(new_n442), .C2(new_n445), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n946), .A2(new_n740), .A3(new_n872), .A4(new_n456), .ZN(new_n947));
  NOR4_X1   g761(.A1(new_n780), .A2(new_n691), .A3(new_n818), .A4(new_n740), .ZN(new_n948));
  AOI22_X1  g762(.A1(new_n945), .A2(new_n947), .B1(new_n948), .B2(new_n839), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n841), .A2(new_n949), .A3(new_n843), .A4(new_n848), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT52), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT115), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n676), .A2(new_n677), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n864), .B2(G469), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n740), .A2(new_n679), .A3(new_n752), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n815), .B1(new_n652), .B2(new_n763), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n838), .A2(new_n314), .ZN(new_n959));
  INV_X1    g773(.A(new_n956), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(KEYINPUT115), .A3(new_n960), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n756), .A2(new_n782), .A3(new_n824), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n952), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n756), .A2(new_n782), .A3(new_n824), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(KEYINPUT52), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n951), .A2(KEYINPUT53), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT117), .ZN(new_n970));
  INV_X1    g784(.A(new_n944), .ZN(new_n971));
  INV_X1    g785(.A(new_n950), .ZN(new_n972));
  NAND2_X1  g786(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n962), .B2(new_n963), .ZN(new_n975));
  NOR2_X1   g789(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n965), .A2(new_n966), .A3(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n971), .A2(new_n972), .A3(new_n975), .A4(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT53), .ZN(new_n980));
  AOI22_X1  g794(.A1(new_n969), .A2(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n951), .A2(KEYINPUT117), .A3(new_n968), .A4(KEYINPUT53), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n938), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR4_X1   g797(.A1(new_n810), .A2(new_n815), .A3(new_n816), .A4(new_n798), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT107), .B1(new_n817), .B2(new_n819), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n789), .A2(new_n793), .A3(new_n796), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT118), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT118), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n939), .A2(new_n989), .A3(new_n821), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n943), .A2(new_n942), .A3(KEYINPUT53), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n975), .A2(new_n978), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n992), .A2(new_n993), .A3(new_n950), .ZN(new_n994));
  AOI21_X1  g808(.A(KEYINPUT53), .B1(new_n951), .B2(new_n968), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT54), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n937), .A2(new_n983), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(G952), .A2(G953), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n900), .B1(new_n997), .B2(new_n998), .ZN(G75));
  AND2_X1   g813(.A1(new_n964), .A2(new_n967), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n986), .A2(new_n987), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n943), .A2(new_n942), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n945), .A2(new_n947), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n948), .A2(new_n839), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n848), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n844), .A2(new_n1001), .A3(new_n1002), .A4(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n980), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n975), .A2(new_n978), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n943), .A2(new_n942), .A3(KEYINPUT53), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n939), .A2(new_n821), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(KEYINPUT118), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1008), .A2(new_n972), .A3(new_n990), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1013), .A2(G210), .A3(G902), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n490), .A2(new_n492), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(new_n515), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT55), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g832(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1019));
  AND3_X1   g833(.A1(new_n1014), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT56), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1018), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n288), .A2(G952), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(G51));
  XNOR2_X1  g838(.A(new_n193), .B(KEYINPUT57), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n938), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n996), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n675), .ZN(new_n1028));
  OAI211_X1 g842(.A(G902), .B(new_n865), .C1(new_n994), .C2(new_n995), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT121), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1023), .B1(new_n1028), .B2(new_n1031), .ZN(G54));
  NAND2_X1  g846(.A1(new_n373), .A2(new_n379), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1013), .A2(G902), .ZN(new_n1034));
  NAND2_X1  g848(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1023), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g852(.A1(new_n1034), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1038), .A2(new_n1039), .ZN(G60));
  XNOR2_X1  g854(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n436), .A2(new_n190), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1041), .B(new_n1042), .Z(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n907), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1045), .B1(new_n996), .B2(new_n1026), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n1037), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1043), .B1(new_n983), .B2(new_n996), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1047), .B1(new_n907), .B2(new_n1048), .ZN(G63));
  XOR2_X1   g863(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n1050));
  NAND2_X1  g864(.A1(G217), .A2(G902), .ZN(new_n1051));
  XNOR2_X1  g865(.A(new_n1051), .B(KEYINPUT60), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1052), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n1053), .A2(new_n566), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n737), .A2(new_n738), .ZN(new_n1055));
  INV_X1    g869(.A(new_n1052), .ZN(new_n1056));
  OAI211_X1 g870(.A(new_n1055), .B(new_n1056), .C1(new_n994), .C2(new_n995), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1057), .A2(new_n1037), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1050), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g873(.A(KEYINPUT61), .B1(new_n1053), .B2(new_n566), .ZN(new_n1060));
  INV_X1    g874(.A(KEYINPUT124), .ZN(new_n1061));
  NOR3_X1   g875(.A1(new_n1060), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1023), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1063));
  INV_X1    g877(.A(KEYINPUT61), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1056), .B1(new_n994), .B2(new_n995), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n1064), .B1(new_n1065), .B2(new_n574), .ZN(new_n1066));
  AOI21_X1  g880(.A(KEYINPUT124), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n1059), .B1(new_n1062), .B2(new_n1067), .ZN(G66));
  OAI21_X1  g882(.A(G953), .B1(new_n453), .B2(new_n496), .ZN(new_n1069));
  OAI21_X1  g883(.A(new_n1069), .B1(new_n971), .B2(G953), .ZN(new_n1070));
  OAI211_X1 g884(.A(new_n490), .B(new_n492), .C1(G898), .C2(new_n288), .ZN(new_n1071));
  XNOR2_X1  g885(.A(new_n1070), .B(new_n1071), .ZN(G69));
  AOI21_X1  g886(.A(new_n288), .B1(G227), .B2(G900), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n593), .B1(KEYINPUT30), .B2(new_n628), .ZN(new_n1074));
  XOR2_X1   g888(.A(new_n1074), .B(KEYINPUT125), .Z(new_n1075));
  XNOR2_X1  g889(.A(new_n1075), .B(new_n368), .ZN(new_n1076));
  AOI21_X1  g890(.A(new_n1076), .B1(G900), .B2(G953), .ZN(new_n1077));
  INV_X1    g891(.A(new_n1077), .ZN(new_n1078));
  NOR2_X1   g892(.A1(new_n912), .A2(new_n815), .ZN(new_n1079));
  NAND2_X1  g893(.A1(new_n871), .A2(new_n1079), .ZN(new_n1080));
  AND3_X1   g894(.A1(new_n844), .A2(new_n848), .A3(new_n965), .ZN(new_n1081));
  AND4_X1   g895(.A1(new_n884), .A2(new_n1080), .A3(new_n892), .A4(new_n1081), .ZN(new_n1082));
  AOI21_X1  g896(.A(new_n1078), .B1(new_n1082), .B2(new_n288), .ZN(new_n1083));
  INV_X1    g897(.A(new_n1076), .ZN(new_n1084));
  INV_X1    g898(.A(KEYINPUT62), .ZN(new_n1085));
  OR3_X1    g899(.A1(new_n778), .A2(new_n1085), .A3(new_n963), .ZN(new_n1086));
  OAI21_X1  g900(.A(new_n1085), .B1(new_n778), .B2(new_n963), .ZN(new_n1087));
  NAND3_X1  g901(.A1(new_n873), .A2(new_n940), .A3(new_n446), .ZN(new_n1088));
  NOR2_X1   g902(.A1(new_n1088), .A2(new_n775), .ZN(new_n1089));
  AOI22_X1  g903(.A1(new_n1086), .A2(new_n1087), .B1(new_n668), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g904(.A1(new_n884), .A2(new_n892), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g905(.A(new_n1084), .B1(new_n1091), .B2(new_n288), .ZN(new_n1092));
  OAI21_X1  g906(.A(new_n1073), .B1(new_n1083), .B2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g907(.A1(new_n884), .A2(new_n1080), .A3(new_n892), .A4(new_n1081), .ZN(new_n1094));
  OAI21_X1  g908(.A(new_n1077), .B1(new_n1094), .B2(G953), .ZN(new_n1095));
  INV_X1    g909(.A(new_n1073), .ZN(new_n1096));
  AND2_X1   g910(.A1(new_n1091), .A2(new_n288), .ZN(new_n1097));
  OAI211_X1 g911(.A(new_n1095), .B(new_n1096), .C1(new_n1097), .C2(new_n1084), .ZN(new_n1098));
  NAND2_X1  g912(.A1(new_n1093), .A2(new_n1098), .ZN(G72));
  XNOR2_X1  g913(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1100));
  NOR2_X1   g914(.A1(new_n690), .A2(new_n190), .ZN(new_n1101));
  XOR2_X1   g915(.A(new_n1100), .B(new_n1101), .Z(new_n1102));
  OAI21_X1  g916(.A(new_n1102), .B1(new_n1094), .B2(new_n944), .ZN(new_n1103));
  NAND2_X1  g917(.A1(new_n658), .A2(new_n603), .ZN(new_n1104));
  XNOR2_X1  g918(.A(new_n1104), .B(KEYINPUT127), .ZN(new_n1105));
  NAND2_X1  g919(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g920(.A(new_n1102), .B1(new_n1091), .B2(new_n944), .ZN(new_n1107));
  INV_X1    g921(.A(new_n658), .ZN(new_n1108));
  NAND3_X1  g922(.A1(new_n1107), .A2(new_n602), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g923(.A1(new_n981), .A2(new_n982), .ZN(new_n1110));
  INV_X1    g924(.A(new_n1102), .ZN(new_n1111));
  NAND2_X1  g925(.A1(new_n1108), .A2(new_n603), .ZN(new_n1112));
  AOI21_X1  g926(.A(new_n1111), .B1(new_n758), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g927(.A(new_n1023), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  AND3_X1   g928(.A1(new_n1106), .A2(new_n1109), .A3(new_n1114), .ZN(G57));
endmodule


