//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g024(.A(G2106), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT69), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n453), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  OR2_X1    g034(.A1(new_n456), .A2(new_n450), .ZN(new_n460));
  INV_X1    g035(.A(new_n457), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G125), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n468), .B1(new_n472), .B2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n473), .A2(new_n474), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n471), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n471), .B2(G112), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G138), .B(new_n471), .C1(new_n473), .C2(new_n474), .ZN(new_n489));
  OR2_X1    g064(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n465), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(new_n471), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n495));
  OAI21_X1  g070(.A(G138), .B1(KEYINPUT71), .B2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n465), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G102), .A2(G2104), .ZN(new_n499));
  AOI21_X1  g074(.A(G2105), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n494), .A2(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(G543), .B1(new_n502), .B2(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OR3_X1    g083(.A1(new_n507), .A2(KEYINPUT73), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT73), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(G50), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n507), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n512), .A2(G651), .B1(new_n513), .B2(new_n516), .ZN(G166));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n507), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(G89), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n527));
  INV_X1    g102(.A(G63), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n507), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n522), .A2(KEYINPUT74), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n513), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n532), .A2(new_n534), .A3(G543), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT75), .B(G51), .Z(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n531), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND3_X1  g114(.A1(new_n532), .A2(new_n534), .A3(G543), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n503), .A2(new_n506), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(new_n513), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n540), .A2(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n542), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n518), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n507), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n518), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n553), .B1(new_n552), .B2(new_n551), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n535), .A2(G43), .B1(G81), .B2(new_n523), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n540), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n505), .B1(new_n522), .B2(KEYINPUT74), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .A3(G53), .A4(new_n534), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT77), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n565), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n507), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(new_n523), .B2(G91), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n569), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n577));
  INV_X1    g152(.A(new_n575), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n568), .B2(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(new_n571), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND2_X1  g160(.A1(new_n523), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n542), .B2(G74), .ZN(new_n587));
  INV_X1    g162(.A(G49), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n586), .B(new_n587), .C1(new_n540), .C2(new_n588), .ZN(G288));
  NAND4_X1  g164(.A1(new_n513), .A2(G86), .A3(new_n503), .A4(new_n506), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n513), .A2(G48), .A3(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n503), .A2(new_n506), .A3(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n518), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n592), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n535), .A2(G47), .B1(G85), .B2(new_n523), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n542), .A2(G60), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n518), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n540), .A2(new_n604), .B1(new_n543), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT79), .B1(new_n606), .B2(new_n601), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n523), .A2(G92), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT80), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n507), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n535), .A2(G54), .B1(G651), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g193(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G321));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NOR2_X1   g197(.A1(G286), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G299), .B(KEYINPUT81), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n622), .ZN(G297));
  AOI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(new_n622), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n619), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n619), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n481), .A2(G2104), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n481), .A2(G135), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT82), .Z(new_n640));
  OR2_X1    g215(.A1(new_n471), .A2(G111), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(KEYINPUT83), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n641), .B2(KEYINPUT83), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n642), .A2(new_n644), .B1(new_n483), .B2(G123), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G2096), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n637), .A2(new_n638), .A3(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT14), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n655), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(new_n664), .A3(G14), .ZN(G401));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT17), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  OR3_X1    g246(.A1(new_n668), .A2(new_n666), .A3(new_n669), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n666), .A3(new_n669), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n647), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n688), .B(new_n687), .S(new_n680), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT84), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  INV_X1    g270(.A(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n694), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n557), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n701), .B2(G19), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(G1341), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G26), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n481), .A2(G140), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n483), .A2(G128), .ZN(new_n710));
  OR2_X1    g285(.A1(G104), .A2(G2105), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n711), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT91), .A4(new_n712), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n708), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2067), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n704), .A2(G1341), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n705), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n706), .A2(G35), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G162), .B2(new_n706), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT29), .Z(new_n724));
  INV_X1    g299(.A(G2090), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n706), .A2(G32), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT26), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n481), .A2(G141), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n483), .A2(G129), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(new_n706), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n724), .A2(new_n725), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT24), .ZN(new_n740));
  INV_X1    g315(.A(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G160), .B2(new_n706), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G2084), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n726), .A2(new_n738), .A3(new_n739), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n701), .A2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G168), .B2(new_n701), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1966), .ZN(new_n749));
  INV_X1    g324(.A(G28), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(KEYINPUT30), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n750), .B2(KEYINPUT30), .ZN(new_n752));
  OR2_X1    g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  NAND2_X1  g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n751), .A2(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n646), .B2(new_n706), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n706), .A2(G33), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT25), .Z(new_n759));
  INV_X1    g334(.A(G139), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n465), .A2(new_n471), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(new_n471), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n757), .B1(new_n765), .B2(new_n706), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n756), .B1(G2072), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n706), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n706), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n767), .B(new_n771), .C1(G2072), .C2(new_n766), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n721), .A2(new_n746), .A3(new_n749), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n619), .A2(new_n701), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G4), .B2(new_n701), .ZN(new_n775));
  INV_X1    g350(.A(G1348), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n701), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n701), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT93), .B(G1961), .Z(new_n781));
  OAI22_X1  g356(.A1(new_n780), .A2(new_n781), .B1(G2084), .B2(new_n744), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n773), .A2(new_n777), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n701), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT94), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n701), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G288), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT33), .B(G1976), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n795), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G1971), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n701), .A2(G22), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n799), .B(new_n800), .C1(G166), .C2(new_n701), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(G166), .B2(new_n701), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G1971), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n701), .A2(G6), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n592), .A2(new_n595), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n701), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n798), .A2(new_n801), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT87), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n481), .A2(G131), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n483), .A2(G119), .ZN(new_n814));
  OR2_X1    g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT85), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n706), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n706), .A2(G25), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n812), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n821), .A2(new_n812), .A3(new_n822), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n809), .A2(KEYINPUT34), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G1986), .ZN(new_n828));
  NAND2_X1  g403(.A1(G290), .A2(G16), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n701), .A2(G24), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n701), .B1(new_n603), .B2(new_n607), .ZN(new_n832));
  INV_X1    g407(.A(new_n830), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n832), .A2(G1986), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT86), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n831), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n829), .A2(new_n828), .A3(new_n830), .ZN(new_n837));
  OAI21_X1  g412(.A(G1986), .B1(new_n832), .B2(new_n833), .ZN(new_n838));
  AOI21_X1  g413(.A(KEYINPUT86), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n811), .B1(new_n827), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n835), .B1(new_n831), .B2(new_n834), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n837), .A2(KEYINPUT86), .A3(new_n838), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n844), .A2(new_n826), .A3(KEYINPUT87), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n810), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT88), .ZN(new_n848));
  INV_X1    g423(.A(new_n810), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n827), .A2(new_n840), .A3(new_n811), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT87), .B1(new_n844), .B2(new_n826), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT88), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n848), .A2(KEYINPUT36), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n847), .B1(new_n855), .B2(KEYINPUT89), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT89), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n848), .A2(new_n854), .A3(new_n857), .A4(KEYINPUT36), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(KEYINPUT90), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT36), .B1(new_n852), .B2(new_n853), .ZN(new_n860));
  AOI211_X1 g435(.A(KEYINPUT88), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT89), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n847), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT90), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n792), .B1(new_n859), .B2(new_n866), .ZN(G311));
  AOI21_X1  g442(.A(KEYINPUT90), .B1(new_n856), .B2(new_n858), .ZN(new_n868));
  AND4_X1   g443(.A1(KEYINPUT90), .A2(new_n862), .A3(new_n858), .A4(new_n863), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n791), .B1(new_n868), .B2(new_n869), .ZN(G150));
  XOR2_X1   g445(.A(KEYINPUT95), .B(G55), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n535), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(G80), .A2(G543), .ZN(new_n873));
  INV_X1    g448(.A(G67), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n507), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G651), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n523), .A2(G93), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT98), .B(G860), .Z(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT37), .Z(new_n882));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n556), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n878), .A2(new_n883), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n872), .A2(KEYINPUT96), .A3(new_n876), .A4(new_n877), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n556), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT38), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n619), .A2(G559), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT97), .Z(new_n894));
  OAI21_X1  g469(.A(new_n879), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n882), .B1(new_n894), .B2(new_n895), .ZN(G145));
  XNOR2_X1  g471(.A(new_n646), .B(G162), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(G160), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n717), .A2(G164), .ZN(new_n899));
  INV_X1    g474(.A(new_n735), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n715), .B(new_n716), .C1(new_n500), .C2(new_n494), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n904));
  OAI22_X1  g479(.A1(new_n903), .A2(new_n904), .B1(new_n764), .B2(new_n762), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n765), .A3(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n819), .A2(new_n820), .ZN(new_n909));
  INV_X1    g484(.A(new_n634), .ZN(new_n910));
  OR2_X1    g485(.A1(G106), .A2(G2105), .ZN(new_n911));
  INV_X1    g486(.A(G2104), .ZN(new_n912));
  INV_X1    g487(.A(G118), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(G2105), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n483), .A2(G130), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT99), .B1(new_n481), .B2(G142), .ZN(new_n916));
  AND4_X1   g491(.A1(KEYINPUT99), .A2(new_n465), .A3(G142), .A4(new_n471), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n918), .A2(KEYINPUT100), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(KEYINPUT100), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n910), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n910), .B1(new_n919), .B2(new_n920), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n909), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n634), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n926), .A2(new_n820), .A3(new_n819), .A4(new_n921), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n908), .A2(KEYINPUT103), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT103), .B1(new_n908), .B2(new_n928), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n928), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n932), .A2(KEYINPUT101), .A3(new_n907), .A4(new_n905), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n908), .B2(new_n928), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n933), .B2(new_n935), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n898), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n933), .A2(new_n935), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n898), .B1(new_n928), .B2(new_n908), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g520(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n580), .A2(new_n581), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n619), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n577), .A2(new_n582), .A3(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT41), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT41), .B1(new_n948), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n629), .B(new_n888), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n948), .A2(new_n950), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(G290), .B(KEYINPUT104), .ZN(new_n960));
  XNOR2_X1  g535(.A(G166), .B(KEYINPUT105), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n960), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(G288), .B(G305), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n960), .A2(new_n961), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n961), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n956), .B1(new_n955), .B2(new_n958), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n959), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n959), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(G868), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n878), .A2(new_n622), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(G295));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n975), .ZN(G331));
  NAND3_X1  g552(.A1(new_n884), .A2(new_n887), .A3(G286), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G286), .B1(new_n884), .B2(new_n887), .ZN(new_n980));
  OAI21_X1  g555(.A(G301), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n980), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(G171), .A3(new_n978), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n957), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n953), .B2(new_n984), .ZN(new_n986));
  INV_X1    g561(.A(new_n969), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n969), .B(new_n985), .C1(new_n953), .C2(new_n984), .ZN(new_n989));
  INV_X1    g564(.A(G37), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n992));
  AOI21_X1  g567(.A(G37), .B1(new_n986), .B2(new_n987), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n994), .A3(new_n989), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n996), .B(new_n997), .ZN(G397));
  INV_X1    g573(.A(G2067), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n717), .B(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(G126), .B1(new_n473), .B2(new_n474), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G114), .A2(G2104), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1003), .A2(G2105), .B1(new_n491), .B2(new_n489), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n490), .A2(G138), .A3(new_n495), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n499), .B1(new_n1005), .B2(new_n480), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n471), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n466), .A2(new_n467), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n471), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT70), .B1(new_n477), .B2(G2105), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n469), .B(new_n471), .C1(new_n475), .C2(new_n476), .ZN(new_n1013));
  OAI211_X1 g588(.A(G40), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  OR3_X1    g591(.A1(new_n1000), .A2(KEYINPUT107), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT107), .B1(new_n1000), .B2(new_n1016), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1016), .ZN(new_n1019));
  INV_X1    g594(.A(G1996), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n735), .B(new_n1020), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1017), .A2(new_n1018), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n909), .B(new_n812), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1016), .B1(new_n1023), .B2(KEYINPUT108), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(KEYINPUT108), .B2(new_n1023), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(G290), .B(new_n828), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n1016), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1014), .B1(KEYINPUT45), .B2(new_n1008), .ZN(new_n1029));
  INV_X1    g604(.A(G1384), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n494), .B2(new_n500), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT109), .B1(new_n1008), .B2(KEYINPUT45), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1029), .A2(new_n770), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT119), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1040), .A3(new_n1037), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1014), .B1(new_n1042), .B2(new_n1008), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1031), .A2(KEYINPUT50), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1961), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1009), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1048), .A2(new_n1029), .A3(KEYINPUT53), .A4(new_n770), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1039), .A2(new_n1041), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G171), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1038), .A2(KEYINPUT119), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n770), .A2(KEYINPUT120), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n770), .A2(KEYINPUT120), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT53), .B(G40), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1055), .B(new_n468), .C1(G2105), .C2(new_n477), .ZN(new_n1056));
  OAI211_X1 g631(.A(KEYINPUT45), .B(new_n1030), .C1(new_n494), .C2(new_n500), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1048), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1052), .A2(G301), .A3(new_n1041), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1051), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n1063));
  NAND3_X1  g638(.A1(G303), .A2(new_n1063), .A3(G8), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT55), .B1(G166), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1029), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1042), .B(new_n1030), .C1(new_n494), .C2(new_n500), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1044), .A2(new_n1015), .A3(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1068), .A2(new_n799), .B1(new_n1070), .B2(new_n725), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1067), .B1(new_n1071), .B2(new_n1065), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1057), .A2(G40), .A3(G160), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1032), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1971), .B1(new_n1076), .B2(new_n1034), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1045), .A2(G2090), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1073), .B(G8), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G288), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1014), .B2(new_n1031), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT110), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT110), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1084), .B(G8), .C1(new_n1014), .C2(new_n1031), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1081), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n1080), .ZN(new_n1087));
  INV_X1    g662(.A(new_n595), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(new_n696), .A3(new_n590), .A4(new_n591), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  NAND3_X1  g667(.A1(G305), .A2(new_n1092), .A3(G1981), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT49), .B1(new_n805), .B2(new_n696), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1091), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1086), .A2(new_n1087), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1098), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT52), .B1(new_n1100), .B2(new_n1081), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1072), .A2(new_n1079), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G2084), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1043), .A2(new_n1103), .A3(new_n1044), .ZN(new_n1104));
  INV_X1    g679(.A(G1966), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1074), .B2(new_n1009), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(new_n1106), .A3(KEYINPUT118), .ZN(new_n1110));
  AOI21_X1  g685(.A(G286), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT51), .B1(new_n1111), .B2(new_n1065), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1110), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT118), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(G168), .A2(new_n1065), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1104), .A2(new_n1106), .A3(G168), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1065), .A2(KEYINPUT51), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1115), .A2(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1102), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1062), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1052), .A2(G301), .A3(new_n1041), .A4(new_n1049), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT54), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1052), .A2(new_n1124), .A3(new_n1041), .A4(new_n1058), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1039), .A2(new_n1041), .A3(new_n1047), .A4(new_n1058), .ZN(new_n1126));
  AOI21_X1  g701(.A(G301), .B1(new_n1126), .B2(KEYINPUT121), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1123), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT122), .B1(new_n1121), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1125), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1123), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1062), .A4(new_n1120), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1029), .A2(new_n1020), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT58), .B(G1341), .Z(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1014), .B2(new_n1031), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n556), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT59), .B1(new_n1138), .B2(KEYINPUT114), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT114), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1140), .B(new_n556), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1138), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT115), .B(KEYINPUT59), .Z(new_n1143));
  OAI22_X1  g718(.A1(new_n1139), .A2(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1015), .A2(new_n999), .A3(new_n1008), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1070), .B2(G1348), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n949), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n619), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n949), .B(new_n1145), .C1(new_n1070), .C2(G1348), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1147), .B1(new_n1150), .B2(KEYINPUT60), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT112), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n568), .A2(new_n578), .A3(KEYINPUT57), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1152), .B(new_n1154), .C1(new_n576), .C2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n579), .B2(new_n571), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT112), .B1(new_n1157), .B2(new_n1153), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1045), .A2(new_n789), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT56), .B(G2072), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1076), .A2(new_n1034), .A3(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT61), .B1(new_n1162), .B2(KEYINPUT116), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1144), .A2(new_n1151), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1161), .A2(new_n1159), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT117), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n1162), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1156), .A2(new_n1158), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT117), .ZN(new_n1171));
  NOR2_X1   g746(.A1(KEYINPUT116), .A2(KEYINPUT61), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1164), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1162), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1170), .A2(KEYINPUT113), .B1(new_n619), .B2(new_n1146), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT113), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1167), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1175), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1174), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1129), .A2(new_n1134), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1184));
  NOR2_X1   g759(.A1(G288), .A2(G1976), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1184), .A2(new_n1185), .B1(new_n696), .B2(new_n805), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n1183), .A2(new_n1079), .B1(new_n1186), .B2(new_n1100), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1107), .A2(G8), .A3(G168), .ZN(new_n1189));
  OR3_X1    g764(.A1(new_n1102), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1188), .B1(new_n1102), .B2(new_n1189), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1187), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(KEYINPUT62), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1112), .A2(new_n1119), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1102), .A2(new_n1051), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1192), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1028), .B1(new_n1182), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n909), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1022), .A2(new_n812), .A3(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n717), .A2(G2067), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1019), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n1205), .A2(KEYINPUT123), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(KEYINPUT123), .ZN(new_n1207));
  AOI21_X1  g782(.A(KEYINPUT46), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1000), .A2(new_n735), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1208), .B1(new_n1209), .B2(new_n1019), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1019), .A2(KEYINPUT46), .A3(new_n1020), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1210), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT47), .ZN(new_n1216));
  NOR3_X1   g791(.A1(G290), .A2(new_n1016), .A3(G1986), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1217), .B(KEYINPUT125), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(KEYINPUT48), .ZN(new_n1219));
  OR2_X1    g794(.A1(new_n1218), .A2(KEYINPUT48), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1026), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  NAND4_X1  g796(.A1(new_n1206), .A2(new_n1207), .A3(new_n1216), .A4(new_n1221), .ZN(new_n1222));
  OAI21_X1  g797(.A(KEYINPUT126), .B1(new_n1201), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n1224));
  AND4_X1   g799(.A1(new_n1206), .A2(new_n1207), .A3(new_n1216), .A4(new_n1221), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1179), .B1(new_n1164), .B2(new_n1173), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1132), .A2(new_n1062), .A3(new_n1120), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1226), .B1(new_n1227), .B2(KEYINPUT122), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1199), .B1(new_n1228), .B2(new_n1134), .ZN(new_n1229));
  OAI211_X1 g804(.A(new_n1224), .B(new_n1225), .C1(new_n1229), .C2(new_n1028), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1223), .A2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g806(.A1(G401), .A2(G227), .A3(new_n463), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n699), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g808(.A(new_n1234), .B1(new_n940), .B2(new_n943), .ZN(new_n1235));
  AND3_X1   g809(.A1(new_n993), .A2(new_n994), .A3(new_n989), .ZN(new_n1236));
  AOI21_X1  g810(.A(new_n994), .B1(new_n993), .B2(new_n989), .ZN(new_n1237));
  OAI211_X1 g811(.A(new_n1235), .B(KEYINPUT127), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  INV_X1    g812(.A(new_n1238), .ZN(new_n1239));
  AOI21_X1  g813(.A(KEYINPUT127), .B1(new_n996), .B2(new_n1235), .ZN(new_n1240));
  NOR2_X1   g814(.A1(new_n1239), .A2(new_n1240), .ZN(G308));
  NAND2_X1  g815(.A1(new_n996), .A2(new_n1235), .ZN(G225));
endmodule


