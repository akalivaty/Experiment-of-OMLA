//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT65), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n465), .B2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n463), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n466), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OR2_X1    g052(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OR3_X1    g055(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n472), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n476), .B(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(new_n480), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT71), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT72), .Z(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n485), .A2(new_n470), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n485), .A2(KEYINPUT70), .A3(new_n470), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(G136), .B2(new_n497), .ZN(G162));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n474), .A2(new_n475), .A3(new_n466), .A4(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT73), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n478), .A2(G138), .A3(new_n479), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT4), .B1(new_n476), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G138), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n460), .A2(new_n461), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n464), .A2(new_n466), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n505), .A2(new_n506), .B1(new_n508), .B2(new_n513), .ZN(G164));
  NAND2_X1  g089(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n520), .A2(G543), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n522), .A2(G88), .B1(new_n523), .B2(G50), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  AND2_X1   g100(.A1(G75), .A2(G543), .ZN(new_n526));
  AND3_X1   g101(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(G543), .B1(KEYINPUT74), .B2(KEYINPUT5), .ZN(new_n528));
  OAI21_X1  g103(.A(G62), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n526), .B1(new_n529), .B2(KEYINPUT75), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n519), .A2(new_n531), .A3(G62), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n525), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n524), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI211_X1 g110(.A(KEYINPUT76), .B(new_n525), .C1(new_n530), .C2(new_n532), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(G166));
  XOR2_X1   g112(.A(KEYINPUT78), .B(KEYINPUT7), .Z(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n522), .A2(G89), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT77), .B(G51), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n523), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G168));
  AOI22_X1  g121(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n525), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT79), .B(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n520), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n521), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n548), .A2(new_n552), .ZN(G171));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n521), .A2(new_n554), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n525), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G860), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT81), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g140(.A(KEYINPUT82), .B(KEYINPUT8), .Z(new_n566));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(new_n523), .A2(G53), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n527), .A2(new_n528), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(G91), .A2(new_n522), .B1(new_n575), .B2(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n571), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  XNOR2_X1  g153(.A(new_n545), .B(KEYINPUT83), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  AOI22_X1  g155(.A1(new_n522), .A2(G87), .B1(new_n523), .B2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n573), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n523), .B2(G48), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n519), .A2(G86), .A3(new_n520), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n525), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n521), .A2(new_n595), .B1(new_n550), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(G301), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n519), .A2(G92), .A3(new_n520), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n573), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(new_n523), .B2(G54), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT85), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(new_n600), .ZN(G284));
  XOR2_X1   g185(.A(G284), .B(KEYINPUT86), .Z(G321));
  NOR2_X1   g186(.A1(G299), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G286), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  AOI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G280));
  INV_X1    g190(.A(new_n609), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G559), .B2(new_n562), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT87), .Z(G148));
  NAND2_X1  g193(.A1(new_n561), .A2(new_n600), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n616), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n600), .ZN(G323));
  XOR2_X1   g196(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n622));
  XNOR2_X1  g197(.A(G323), .B(new_n622), .ZN(G282));
  NAND2_X1  g198(.A1(new_n497), .A2(G135), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n480), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n486), .B2(G123), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n624), .A2(new_n631), .A3(new_n628), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n632), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT89), .ZN(new_n652));
  INV_X1    g227(.A(G14), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n649), .B2(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n636), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n631), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  AOI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n670), .C2(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT91), .ZN(new_n679));
  XOR2_X1   g254(.A(G1981), .B(G1986), .Z(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT90), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n679), .B(new_n685), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  MUX2_X1   g262(.A(G23), .B(G288), .S(G16), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT33), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1976), .ZN(new_n690));
  NAND2_X1  g265(.A1(G166), .A2(G16), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G16), .B2(G22), .ZN(new_n692));
  INV_X1    g267(.A(G1971), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  MUX2_X1   g270(.A(G6), .B(G305), .S(G16), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT93), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n690), .A2(new_n694), .A3(new_n695), .A4(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT34), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n497), .A2(G131), .ZN(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n706));
  INV_X1    g281(.A(G107), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n480), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n486), .B2(G119), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n704), .B1(new_n711), .B2(new_n703), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT35), .B(G1991), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT92), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT92), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G24), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n598), .B2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(G1986), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n702), .A2(new_n715), .A3(new_n716), .A4(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n717), .A2(G20), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT23), .Z(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G299), .B2(G16), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT98), .ZN(new_n728));
  INV_X1    g303(.A(G1956), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n703), .A2(G35), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G162), .B2(new_n703), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT29), .Z(new_n733));
  INV_X1    g308(.A(G2090), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT99), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g312(.A(KEYINPUT99), .B(new_n730), .C1(new_n733), .C2(new_n734), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n733), .A2(new_n734), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n497), .A2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  NAND3_X1  g317(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n486), .B2(G129), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(new_n703), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n703), .B2(G32), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n703), .A2(G33), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n497), .A2(G139), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT25), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n511), .A2(G127), .ZN(new_n756));
  INV_X1    g331(.A(G115), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n463), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n755), .B1(new_n480), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n752), .B1(new_n760), .B2(G29), .ZN(new_n761));
  INV_X1    g336(.A(G2072), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G171), .A2(new_n717), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G5), .B2(new_n717), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G1966), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n545), .A2(G16), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n717), .A2(G21), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n767), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n768), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n766), .B2(new_n765), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G34), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(G29), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n482), .B2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n703), .A2(G27), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT97), .Z(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G164), .B2(new_n703), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2078), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n772), .A2(new_n774), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT30), .B(G28), .ZN(new_n787));
  OR2_X1    g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  NAND2_X1  g363(.A1(KEYINPUT31), .A2(G11), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n787), .A2(new_n703), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n629), .B2(new_n703), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n751), .A2(new_n763), .A3(new_n786), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n717), .A2(G4), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n609), .B2(new_n717), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G1348), .Z(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n703), .A2(G26), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n497), .A2(G140), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G116), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n480), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n486), .B2(G128), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(G29), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2067), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n717), .A2(G19), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT94), .ZN(new_n810));
  INV_X1    g385(.A(new_n561), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n717), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1341), .Z(new_n813));
  NAND3_X1  g388(.A1(new_n797), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n762), .A2(new_n761), .B1(new_n749), .B2(new_n750), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n791), .A2(new_n792), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n794), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n724), .A2(new_n818), .ZN(G311));
  OR2_X1    g394(.A1(new_n724), .A2(new_n818), .ZN(G150));
  NAND2_X1  g395(.A1(new_n609), .A2(G559), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT38), .Z(new_n822));
  AOI22_X1  g397(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n525), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  INV_X1    g400(.A(G55), .ZN(new_n826));
  OAI22_X1  g401(.A1(new_n521), .A2(new_n825), .B1(new_n550), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n561), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n822), .B(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(new_n562), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n828), .A2(new_n562), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n629), .B(new_n482), .ZN(new_n838));
  XNOR2_X1  g413(.A(G162), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n497), .A2(G142), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n841));
  INV_X1    g416(.A(G118), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n841), .B1(new_n480), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n486), .B2(G130), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(new_n634), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n845), .A2(new_n634), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n710), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n848), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n850), .A2(new_n711), .A3(new_n846), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n760), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n746), .A2(new_n806), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n508), .A2(new_n513), .ZN(new_n856));
  INV_X1    g431(.A(new_n503), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n740), .A2(new_n801), .A3(new_n745), .A4(new_n805), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n855), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n854), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n855), .A2(new_n859), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n503), .B1(new_n508), .B2(new_n513), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n760), .B(new_n853), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n852), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n839), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI211_X1 g446(.A(KEYINPUT103), .B(new_n852), .C1(new_n862), .C2(new_n868), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n862), .A2(new_n868), .A3(new_n852), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT101), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n868), .A2(new_n862), .A3(new_n852), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n869), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n839), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT102), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n869), .B1(new_n875), .B2(new_n877), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n884), .A2(new_n885), .A3(new_n839), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n879), .B(KEYINPUT40), .C1(new_n883), .C2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(KEYINPUT102), .A3(new_n882), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n884), .B2(new_n839), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT40), .B1(new_n891), .B2(new_n879), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n888), .A2(new_n892), .ZN(G395));
  XOR2_X1   g468(.A(G166), .B(G305), .Z(new_n894));
  XNOR2_X1  g469(.A(G288), .B(new_n598), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(KEYINPUT105), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(KEYINPUT105), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n894), .B2(new_n897), .ZN(new_n899));
  XNOR2_X1  g474(.A(G299), .B(new_n608), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(KEYINPUT41), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(KEYINPUT41), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OR3_X1    g479(.A1(new_n900), .A2(new_n902), .A3(KEYINPUT41), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n620), .A2(new_n830), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n561), .B(new_n828), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n616), .B2(G559), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n900), .A3(new_n909), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n899), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  INV_X1    g493(.A(new_n899), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(G868), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n828), .A2(G868), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(G295));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n922), .B2(new_n924), .ZN(new_n927));
  AOI211_X1 g502(.A(KEYINPUT106), .B(new_n923), .C1(new_n921), .C2(G868), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(G331));
  NAND2_X1  g504(.A1(new_n830), .A2(KEYINPUT107), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n908), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G301), .A2(new_n545), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(G286), .B2(G301), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n930), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n900), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n937), .A2(new_n905), .A3(new_n904), .A4(new_n938), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n899), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G37), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n901), .A2(new_n903), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n937), .A2(new_n948), .A3(new_n938), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n899), .B1(new_n941), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n947), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n899), .B1(new_n941), .B2(new_n942), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT43), .B1(new_n945), .B2(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n954), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n946), .A2(new_n947), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n946), .A2(KEYINPUT108), .A3(new_n947), .A4(new_n957), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT43), .B1(new_n945), .B2(new_n950), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n956), .B1(new_n963), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n864), .B2(G1384), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n472), .A2(new_n481), .A3(G40), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n746), .A2(G1996), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n806), .A2(G2067), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n746), .A2(G1996), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n806), .A2(G2067), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n968), .B(KEYINPUT109), .Z(new_n975));
  AOI21_X1  g550(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n711), .A2(new_n713), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n711), .A2(new_n713), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n598), .B(new_n720), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n968), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT73), .B1(new_n500), .B2(new_n502), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT73), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n856), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n989));
  INV_X1    g564(.A(G40), .ZN(new_n990));
  NOR4_X1   g565(.A1(new_n989), .A2(new_n469), .A3(new_n990), .A4(new_n471), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n991), .A3(new_n966), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(G2078), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(G1384), .B1(new_n856), .B2(new_n857), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n967), .B1(new_n996), .B2(KEYINPUT45), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n965), .B1(G164), .B2(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n993), .B1(new_n999), .B2(G2078), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n858), .A2(new_n1002), .A3(new_n987), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n991), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n766), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n995), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(G171), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT123), .Z(new_n1008));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n966), .A2(new_n991), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT121), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n464), .A2(new_n466), .A3(new_n512), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n507), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n510), .A2(new_n474), .A3(new_n466), .A4(new_n475), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1014), .B2(KEYINPUT4), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT45), .B(new_n987), .C1(new_n1015), .C2(new_n503), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT122), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT53), .B1(new_n1017), .B2(G2078), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n1017), .B2(G2078), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1011), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1010), .A2(KEYINPUT121), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1000), .B(new_n1005), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1009), .B1(new_n1022), .B2(G171), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1006), .A2(G171), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n1022), .B2(G171), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1008), .A2(new_n1023), .B1(new_n1009), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1002), .B1(new_n986), .B2(new_n987), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n864), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n991), .A2(new_n780), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1030), .A2(KEYINPUT114), .B1(new_n768), .B2(new_n992), .ZN(new_n1031));
  AND4_X1   g606(.A1(G40), .A2(new_n472), .A3(new_n780), .A4(new_n481), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n505), .A2(new_n506), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n1033), .B2(new_n856), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1003), .B(new_n1032), .C1(new_n1034), .C2(new_n1002), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G168), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g613(.A1(G164), .A2(new_n965), .A3(G1384), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n768), .B1(new_n1039), .B2(new_n1010), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1001), .A2(KEYINPUT114), .A3(new_n1003), .A4(new_n1032), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1037), .A2(new_n1040), .A3(G168), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G8), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT51), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1045), .A3(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1016), .A2(new_n991), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT45), .B1(new_n986), .B2(new_n987), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n693), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1001), .A2(new_n734), .A3(new_n991), .A4(new_n1003), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n535), .B2(new_n536), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT55), .B(G8), .C1(new_n535), .C2(new_n536), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1057), .A3(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n996), .A2(new_n991), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n581), .A2(G1976), .A3(new_n582), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(G8), .A3(new_n1060), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1061), .A2(KEYINPUT110), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(KEYINPUT110), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(KEYINPUT52), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n587), .A2(new_n588), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G1981), .ZN(new_n1066));
  INV_X1    g641(.A(G1981), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n587), .A2(new_n590), .A3(new_n1067), .A4(new_n591), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT49), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1059), .A2(G8), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1068), .A3(KEYINPUT49), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1061), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT111), .B(G1976), .Z(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1071), .A2(new_n1072), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1058), .A2(new_n1064), .A3(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT112), .B(new_n991), .C1(new_n996), .C2(new_n1002), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n986), .A2(new_n1002), .A3(new_n987), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT50), .B1(new_n864), .B2(G1384), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT112), .B1(new_n1081), .B2(new_n991), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1080), .A2(G2090), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1050), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT113), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n991), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(new_n1079), .A3(new_n1078), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1086), .B(new_n1050), .C1(new_n1090), .C2(G2090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(G8), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1057), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1077), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1026), .A2(new_n1047), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT117), .B(G1996), .Z(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT58), .B(G1341), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1059), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n561), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT59), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n729), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G299), .B(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1096), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1105), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1102), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1109), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1090), .A2(new_n729), .B1(new_n1096), .B2(new_n1106), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT116), .B1(new_n1114), .B2(new_n1105), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .A4(KEYINPUT116), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1113), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT118), .B1(new_n1118), .B2(new_n1110), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1108), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1109), .B1(new_n1121), .B2(new_n1116), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1122), .A2(new_n1123), .A3(KEYINPUT61), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1112), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1112), .B(KEYINPUT119), .C1(new_n1119), .C2(new_n1124), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1004), .ZN(new_n1129));
  OAI22_X1  g704(.A1(new_n1129), .A2(G1348), .B1(G2067), .B2(new_n1059), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n608), .A2(KEYINPUT120), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n608), .A2(KEYINPUT120), .ZN(new_n1134));
  OR3_X1    g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1135), .B(new_n1136), .C1(KEYINPUT60), .C2(new_n1131), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1127), .A2(new_n1128), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1113), .B1(new_n1131), .B2(new_n608), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1095), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1044), .A2(new_n1143), .A3(new_n1046), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1024), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1094), .A3(KEYINPUT124), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1047), .A2(KEYINPUT62), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g723(.A(new_n1024), .B(new_n1077), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT124), .B1(new_n1149), .B2(new_n1144), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1142), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1144), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1077), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(new_n1145), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1152), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(KEYINPUT125), .A3(new_n1147), .A4(new_n1146), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1064), .A2(new_n1076), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1068), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1162));
  NOR2_X1   g737(.A1(G288), .A2(G1976), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1160), .A2(new_n1058), .B1(new_n1164), .B2(new_n1070), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n613), .A2(G8), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1052), .A2(G8), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1093), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1155), .A2(new_n1167), .A3(KEYINPUT63), .A4(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT115), .Z(new_n1171));
  AND2_X1   g746(.A1(new_n1094), .A2(new_n1167), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1172), .A2(KEYINPUT63), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1165), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1159), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n983), .B1(new_n1141), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n973), .A2(new_n747), .A3(new_n971), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT46), .B1(new_n969), .B2(G1996), .ZN(new_n1178));
  OR3_X1    g753(.A1(new_n969), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1177), .A2(new_n975), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT47), .Z(new_n1181));
  NAND3_X1  g756(.A1(new_n968), .A2(new_n720), .A3(new_n598), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT48), .Z(new_n1183));
  OAI21_X1  g758(.A(new_n1181), .B1(new_n981), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n975), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n976), .A2(new_n977), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(new_n973), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1187), .A2(KEYINPUT126), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(KEYINPUT126), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1184), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1176), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g766(.A(new_n879), .B1(new_n883), .B2(new_n886), .ZN(new_n1193));
  NOR2_X1   g767(.A1(G227), .A2(new_n458), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n655), .A2(new_n1194), .ZN(new_n1195));
  XOR2_X1   g769(.A(new_n1195), .B(KEYINPUT127), .Z(new_n1196));
  NAND2_X1  g770(.A1(new_n952), .A2(new_n955), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n1193), .A2(new_n1196), .A3(new_n686), .A4(new_n1197), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


