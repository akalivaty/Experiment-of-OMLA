//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n192), .A3(new_n195), .A4(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT0), .B(G128), .Z(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n198), .A2(new_n213), .A3(new_n206), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n207), .A2(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G128), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n209), .A2(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n212), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n191), .A2(G134), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n190), .A2(new_n221), .A3(KEYINPUT65), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(G131), .C1(KEYINPUT65), .C2(new_n221), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n196), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n197), .A2(new_n225), .A3(new_n202), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n204), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT30), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G116), .B(G119), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  XOR2_X1   g045(.A(new_n230), .B(new_n231), .Z(new_n232));
  NAND2_X1  g046(.A1(new_n224), .A2(new_n203), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT30), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n230), .B(new_n231), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n237), .A3(new_n203), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n224), .A2(new_n203), .A3(KEYINPUT67), .A4(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(G101), .ZN(new_n244));
  NOR2_X1   g058(.A1(G237), .A2(G953), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G210), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n244), .B(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n236), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT31), .ZN(new_n249));
  INV_X1    g063(.A(new_n247), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n227), .A2(new_n232), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n242), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n238), .A2(new_n251), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT31), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n236), .A2(new_n257), .A3(new_n242), .A4(new_n247), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n249), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(G472), .A2(G902), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT32), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(KEYINPUT32), .A3(new_n260), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n240), .A2(new_n241), .B1(new_n232), .B2(new_n233), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n254), .B1(new_n266), .B2(new_n251), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n250), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n265), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n240), .A2(new_n241), .B1(new_n227), .B2(new_n232), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT68), .B(new_n254), .C1(new_n272), .C2(new_n251), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n247), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n236), .A2(new_n242), .A3(new_n250), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n254), .B(new_n247), .C1(new_n272), .C2(new_n251), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT29), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n271), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G472), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n263), .B(new_n264), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G221), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT9), .B(G234), .Z(new_n284));
  AOI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(new_n265), .ZN(new_n285));
  INV_X1    g099(.A(G104), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT3), .B1(new_n286), .B2(G107), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n288));
  INV_X1    g102(.A(G107), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(G104), .ZN(new_n290));
  INV_X1    g104(.A(G101), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(G107), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n287), .A2(new_n290), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n289), .A2(G104), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n286), .A2(G107), .ZN(new_n295));
  OAI21_X1  g109(.A(G101), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT80), .B1(new_n220), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n220), .A2(new_n297), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n220), .A2(new_n297), .A3(KEYINPUT80), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n197), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT12), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g118(.A(KEYINPUT12), .B(new_n197), .C1(new_n300), .C2(new_n301), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT81), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n220), .A2(new_n297), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n220), .A2(new_n297), .A3(KEYINPUT10), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n287), .A2(new_n290), .A3(new_n292), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G101), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT4), .A3(new_n293), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n315), .A3(G101), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(new_n202), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n310), .A2(new_n311), .A3(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n197), .B(KEYINPUT79), .Z(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(G110), .B(G140), .Z(new_n322));
  INV_X1    g136(.A(G227), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G953), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n322), .B(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n304), .A2(new_n327), .A3(new_n305), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n307), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n320), .B1(new_n197), .B2(new_n318), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(new_n325), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G469), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n265), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n318), .A2(new_n197), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n321), .A2(new_n335), .A3(new_n325), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n320), .B1(new_n304), .B2(new_n305), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(new_n325), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n333), .B1(new_n338), .B2(new_n265), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n285), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n342));
  INV_X1    g156(.A(G119), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT69), .B1(new_n343), .B2(G128), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n205), .A3(G119), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n344), .A2(new_n346), .B1(new_n343), .B2(G128), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT24), .B(G110), .Z(new_n348));
  AND3_X1   g162(.A1(new_n347), .A2(KEYINPUT70), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT70), .B1(new_n347), .B2(new_n348), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT23), .B1(new_n343), .B2(G128), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n205), .A3(G119), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n343), .A2(G128), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G110), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT16), .B1(new_n359), .B2(G125), .ZN(new_n360));
  INV_X1    g174(.A(G125), .ZN(new_n361));
  OAI211_X1 g175(.A(KEYINPUT72), .B(G140), .C1(new_n361), .C2(KEYINPUT71), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT72), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n359), .B2(G125), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT71), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n359), .A3(G125), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n360), .B1(new_n367), .B2(KEYINPUT16), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n209), .ZN(new_n369));
  AOI211_X1 g183(.A(G146), .B(new_n360), .C1(new_n367), .C2(KEYINPUT16), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n351), .B(new_n358), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G110), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n355), .A2(new_n372), .A3(new_n356), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n347), .B2(new_n348), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT73), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n367), .A2(KEYINPUT16), .ZN(new_n377));
  OAI21_X1  g191(.A(G146), .B1(new_n377), .B2(new_n360), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n361), .A2(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n359), .A2(G125), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT74), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT74), .B1(new_n379), .B2(new_n380), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n209), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n373), .B(KEYINPUT73), .C1(new_n347), .C2(new_n348), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n376), .A2(new_n378), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(G137), .ZN(new_n387));
  INV_X1    g201(.A(G953), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(G221), .A3(G234), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n387), .B(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n371), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n390), .B1(new_n371), .B2(new_n385), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n391), .A2(new_n392), .A3(G902), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n342), .B1(new_n393), .B2(KEYINPUT76), .ZN(new_n394));
  INV_X1    g208(.A(G217), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(G234), .B2(new_n265), .ZN(new_n396));
  INV_X1    g210(.A(new_n392), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n371), .A2(new_n385), .A3(new_n390), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n265), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT76), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT25), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n396), .A2(G902), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT78), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n397), .B2(new_n398), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT77), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n245), .A2(G214), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n207), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n245), .B(G214), .C1(KEYINPUT86), .C2(G143), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G131), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n413), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n367), .A2(G146), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n383), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n416), .A2(new_n417), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT88), .B1(new_n420), .B2(new_n195), .ZN(new_n425));
  OR3_X1    g239(.A1(new_n420), .A2(new_n195), .A3(KEYINPUT88), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n418), .A2(KEYINPUT87), .A3(KEYINPUT18), .A4(G131), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n421), .A2(new_n423), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n381), .B2(new_n382), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n367), .A2(KEYINPUT19), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n209), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT89), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n431), .A2(new_n435), .A3(new_n209), .A4(new_n432), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n378), .A3(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n437), .A2(KEYINPUT90), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n439), .A3(new_n378), .A4(new_n436), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n424), .A2(new_n195), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n419), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n429), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(G113), .B(G122), .Z(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT91), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(new_n286), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n369), .A2(new_n370), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n441), .A2(new_n450), .A3(new_n419), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n418), .A2(KEYINPUT17), .A3(G131), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n429), .A3(new_n447), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n453), .A2(new_n429), .A3(KEYINPUT92), .A4(new_n447), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n444), .A2(new_n448), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G475), .A2(G902), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n412), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G478), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(KEYINPUT15), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G128), .B(G143), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n188), .ZN(new_n466));
  XOR2_X1   g280(.A(new_n466), .B(KEYINPUT94), .Z(new_n467));
  AOI21_X1  g281(.A(new_n188), .B1(new_n465), .B2(KEYINPUT13), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n207), .A2(G128), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n468), .B1(KEYINPUT13), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT93), .A2(G122), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(KEYINPUT93), .A2(G122), .ZN(new_n473));
  OAI21_X1  g287(.A(G116), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G116), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G122), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(G107), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n289), .B1(new_n474), .B2(new_n476), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n467), .B(new_n470), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n476), .B(KEYINPUT14), .ZN(new_n481));
  INV_X1    g295(.A(new_n474), .ZN(new_n482));
  OAI21_X1  g296(.A(G107), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n465), .B(new_n188), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n483), .B(new_n484), .C1(G107), .C2(new_n477), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n284), .A2(G217), .A3(new_n388), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n487), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n464), .B1(new_n491), .B2(new_n265), .ZN(new_n492));
  AOI211_X1 g306(.A(G902), .B(new_n463), .C1(new_n488), .C2(new_n490), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n456), .A2(new_n457), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n437), .A2(KEYINPUT90), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n442), .A3(new_n440), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n447), .B1(new_n497), .B2(new_n429), .ZN(new_n498));
  OAI211_X1 g312(.A(KEYINPUT20), .B(new_n459), .C1(new_n495), .C2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n447), .B1(new_n453), .B2(new_n429), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n456), .B2(new_n457), .ZN(new_n501));
  OAI21_X1  g315(.A(G475), .B1(new_n501), .B2(G902), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n461), .A2(new_n494), .A3(new_n499), .A4(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n232), .A2(new_n314), .A3(new_n316), .ZN(new_n504));
  XNOR2_X1  g318(.A(G110), .B(G122), .ZN(new_n505));
  INV_X1    g319(.A(G113), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n475), .A2(G119), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n230), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n507), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n510), .A2(new_n231), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n297), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n504), .A2(new_n505), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n293), .A2(new_n296), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(new_n515), .A3(new_n512), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n505), .B(KEYINPUT8), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n510), .A2(new_n231), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n230), .A2(KEYINPUT5), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n518), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n516), .B(new_n517), .C1(new_n520), .C2(new_n515), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n220), .A2(new_n361), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n202), .A2(G125), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n388), .A2(G224), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n525), .B(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n504), .A2(new_n513), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT84), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n532));
  INV_X1    g346(.A(new_n505), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  AOI211_X1 g348(.A(KEYINPUT84), .B(new_n505), .C1(new_n504), .C2(new_n513), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT85), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n523), .B2(new_n524), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n523), .A2(new_n538), .A3(new_n524), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n540), .A2(G224), .A3(new_n388), .A4(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n526), .B1(new_n543), .B2(new_n539), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n529), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(G210), .B1(G237), .B2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT6), .A3(new_n514), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(new_n542), .A3(new_n544), .A4(new_n534), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n547), .A3(new_n529), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G214), .B1(G237), .B2(G902), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT82), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n388), .A2(G952), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(G234), .B2(G237), .ZN(new_n558));
  XOR2_X1   g372(.A(KEYINPUT21), .B(G898), .Z(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(G234), .A2(G237), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(G902), .A3(G953), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n558), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n554), .A2(new_n556), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n503), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n282), .A2(new_n341), .A3(new_n411), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G101), .ZN(G3));
  INV_X1    g383(.A(new_n285), .ZN(new_n570));
  AOI211_X1 g384(.A(G469), .B(G902), .C1(new_n329), .C2(new_n331), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n411), .B(new_n570), .C1(new_n571), .C2(new_n339), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(new_n281), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n259), .B2(new_n265), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n259), .A2(new_n265), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n461), .A2(new_n502), .A3(new_n499), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n555), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n547), .B1(new_n552), .B2(new_n529), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(KEYINPUT96), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n549), .A2(new_n586), .A3(new_n553), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n490), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n489), .B1(new_n480), .B2(new_n485), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n491), .A2(KEYINPUT33), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(G478), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n491), .A2(new_n462), .A3(new_n265), .ZN(new_n596));
  NAND2_X1  g410(.A1(G478), .A2(G902), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NOR4_X1   g412(.A1(new_n582), .A2(new_n588), .A3(new_n564), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n580), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT34), .B(G104), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  NOR4_X1   g416(.A1(new_n588), .A2(new_n581), .A3(new_n494), .A4(new_n564), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n580), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  AOI21_X1  g420(.A(G902), .B1(new_n329), .B2(new_n331), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n339), .B1(new_n607), .B2(new_n333), .ZN(new_n608));
  INV_X1    g422(.A(new_n390), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT36), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n371), .A2(new_n385), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n405), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n402), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n608), .A2(new_n615), .A3(new_n285), .ZN(new_n616));
  INV_X1    g430(.A(new_n578), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n576), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n567), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G110), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n619), .B(new_n621), .ZN(G12));
  AND3_X1   g436(.A1(new_n259), .A2(KEYINPUT32), .A3(new_n260), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT32), .B1(new_n259), .B2(new_n260), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n271), .ZN(new_n626));
  INV_X1    g440(.A(new_n275), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n247), .B2(new_n273), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n277), .A2(new_n278), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n268), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n626), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G472), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n588), .B1(new_n625), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n558), .B1(new_n563), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n461), .A2(new_n502), .A3(new_n499), .A4(new_n636), .ZN(new_n637));
  OR3_X1    g451(.A1(new_n637), .A2(KEYINPUT98), .A3(new_n494), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT98), .B1(new_n637), .B2(new_n494), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n633), .A2(new_n616), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  XNOR2_X1  g455(.A(new_n554), .B(KEYINPUT38), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n570), .B1(new_n571), .B2(new_n339), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n635), .B(KEYINPUT39), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n645), .A2(KEYINPUT101), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n648));
  INV_X1    g462(.A(new_n646), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n341), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n644), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT101), .B1(new_n645), .B2(new_n646), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n341), .A2(new_n648), .A3(new_n649), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT40), .ZN(new_n654));
  AOI211_X1 g468(.A(new_n583), .B(new_n643), .C1(new_n651), .C2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n656));
  INV_X1    g470(.A(new_n266), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n265), .B1(new_n657), .B2(new_n247), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n250), .B1(new_n236), .B2(new_n242), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n656), .B1(new_n625), .B2(new_n660), .ZN(new_n661));
  AND4_X1   g475(.A1(new_n656), .A2(new_n263), .A3(new_n264), .A4(new_n660), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n625), .A2(new_n656), .A3(new_n660), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n263), .A2(new_n264), .A3(new_n660), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT99), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT100), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n494), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n581), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n655), .A2(new_n672), .A3(KEYINPUT102), .A4(new_n615), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n674));
  INV_X1    g488(.A(new_n654), .ZN(new_n675));
  AOI21_X1  g489(.A(KEYINPUT40), .B1(new_n652), .B2(new_n653), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n555), .B(new_n642), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n663), .B1(new_n661), .B2(new_n662), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n665), .A2(new_n667), .A3(KEYINPUT100), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n671), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n615), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n674), .B1(new_n677), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n207), .ZN(G45));
  INV_X1    g499(.A(new_n598), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n581), .A2(new_n686), .A3(new_n636), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n581), .A2(new_n686), .A3(KEYINPUT103), .A4(new_n636), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n633), .A2(new_n616), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  AOI21_X1  g506(.A(new_n410), .B1(new_n625), .B2(new_n632), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n607), .A2(new_n333), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n571), .A3(new_n285), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n599), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND3_X1  g512(.A1(new_n693), .A2(new_n603), .A3(new_n695), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  NOR4_X1   g514(.A1(new_n694), .A2(new_n571), .A3(new_n285), .A4(new_n564), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n615), .A2(new_n503), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n633), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  NAND4_X1  g518(.A1(new_n581), .A2(new_n670), .A3(new_n587), .A4(new_n585), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT108), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n585), .A2(new_n587), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n670), .A4(new_n581), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n410), .A2(KEYINPUT106), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n267), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g527(.A(KEYINPUT104), .B(new_n254), .C1(new_n266), .C2(new_n251), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n250), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n249), .A2(new_n258), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n260), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n402), .A2(new_n719), .A3(new_n409), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n259), .A2(new_n265), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT105), .B(G472), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n711), .A2(new_n718), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n402), .A2(new_n719), .A3(new_n409), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n719), .B1(new_n402), .B2(new_n409), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n260), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n249), .A2(new_n258), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n730), .B1(new_n731), .B2(new_n715), .ZN(new_n732));
  INV_X1    g546(.A(new_n722), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n259), .B2(new_n265), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n726), .B1(new_n729), .B2(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n701), .B(new_n710), .C1(new_n725), .C2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR3_X1   g552(.A1(new_n615), .A2(new_n732), .A3(new_n734), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n689), .A2(new_n695), .A3(new_n739), .A4(new_n690), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n588), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n361), .ZN(G27));
  NAND2_X1  g556(.A1(new_n282), .A2(new_n729), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n689), .A2(new_n690), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n549), .A2(new_n570), .A3(new_n555), .A4(new_n553), .ZN(new_n748));
  OAI211_X1 g562(.A(G469), .B(new_n336), .C1(new_n337), .C2(new_n325), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n607), .B2(new_n333), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n333), .A2(new_n265), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT109), .Z(new_n753));
  AOI21_X1  g567(.A(new_n748), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n745), .A2(new_n747), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n411), .A3(new_n282), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n756), .B(new_n744), .C1(new_n757), .C2(new_n746), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n693), .A2(new_n689), .A3(new_n690), .A4(new_n754), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n756), .B1(new_n760), .B2(new_n744), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n755), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  AND2_X1   g577(.A1(new_n638), .A2(new_n639), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n693), .A3(new_n754), .ZN(new_n765));
  XOR2_X1   g579(.A(KEYINPUT111), .B(G134), .Z(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G36));
  NOR2_X1   g581(.A1(new_n581), .A2(new_n598), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT43), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n581), .B2(new_n598), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n579), .A3(new_n614), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n554), .A2(new_n583), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n772), .A2(KEYINPUT44), .A3(new_n579), .A4(new_n614), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n338), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT45), .B(new_n336), .C1(new_n337), .C2(new_n325), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(G469), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n753), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n571), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n753), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n789), .A2(new_n285), .A3(new_n646), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n775), .A2(KEYINPUT112), .A3(new_n776), .A4(new_n777), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n780), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n789), .B2(new_n285), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n787), .A2(new_n788), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(KEYINPUT47), .A3(new_n570), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n746), .A2(new_n282), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n410), .A3(new_n776), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NAND2_X1  g615(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n729), .A2(new_n726), .A3(new_n735), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n558), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n769), .B2(new_n771), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n642), .A2(new_n555), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n804), .A2(new_n695), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n804), .A2(new_n806), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n694), .A2(new_n571), .A3(new_n570), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n776), .B(new_n811), .C1(new_n798), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n694), .A2(new_n571), .ZN(new_n814));
  INV_X1    g628(.A(new_n748), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n558), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n581), .A2(new_n686), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n669), .A2(new_n411), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n739), .A3(new_n772), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n810), .A2(new_n813), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n557), .B1(new_n821), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n582), .A2(new_n598), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n669), .A2(new_n411), .A3(new_n825), .A4(new_n817), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n811), .A2(new_n707), .A3(new_n695), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n823), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n817), .A2(new_n282), .A3(new_n729), .A4(new_n772), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT48), .Z(new_n830));
  NOR2_X1   g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  INV_X1    g646(.A(new_n566), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n580), .A2(new_n833), .A3(new_n825), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n737), .A2(new_n699), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n696), .A2(new_n703), .A3(new_n568), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n492), .B2(new_n493), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n463), .B1(new_n591), .B2(G902), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n491), .A2(new_n265), .A3(new_n464), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT113), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n502), .A3(new_n461), .A4(new_n499), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n572), .A2(new_n579), .A3(new_n566), .A4(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n341), .A2(new_n618), .A3(new_n567), .A4(new_n614), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n838), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n341), .A2(new_n618), .A3(new_n411), .A4(new_n833), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n619), .B(KEYINPUT114), .C1(new_n849), .C2(new_n845), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n747), .A2(new_n739), .A3(new_n754), .ZN(new_n852));
  INV_X1    g666(.A(new_n844), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n637), .A2(new_n583), .A3(new_n554), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n616), .A2(new_n282), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n852), .A2(new_n765), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n837), .A2(new_n762), .A3(new_n851), .A4(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n640), .B(new_n691), .C1(new_n588), .C2(new_n740), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n614), .B1(new_n751), .B2(new_n753), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n636), .B(new_n860), .C1(new_n661), .C2(new_n662), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n710), .A2(new_n570), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT52), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n741), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n633), .A2(new_n616), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n747), .B2(new_n764), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n285), .B1(new_n706), .B2(new_n709), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n665), .A2(new_n667), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n636), .A4(new_n860), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(new_n867), .A3(new_n868), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n832), .B1(new_n858), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n864), .A2(new_n872), .ZN(new_n875));
  INV_X1    g689(.A(new_n836), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n814), .A2(new_n570), .A3(new_n565), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n802), .B2(new_n803), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n693), .A2(new_n695), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n878), .A2(new_n710), .B1(new_n879), .B2(new_n603), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n851), .A2(new_n876), .A3(new_n834), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n744), .B1(new_n757), .B2(new_n746), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT110), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n758), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n856), .B1(new_n884), .B2(new_n755), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n881), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n874), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT115), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n887), .B1(new_n874), .B2(new_n886), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI211_X1 g705(.A(KEYINPUT115), .B(new_n887), .C1(new_n874), .C2(new_n886), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n831), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT116), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(G952), .A2(G953), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n831), .B(KEYINPUT116), .C1(new_n891), .C2(new_n892), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n680), .A2(new_n285), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n814), .B(KEYINPUT49), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n900), .A2(new_n556), .A3(new_n643), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n899), .A2(new_n729), .A3(new_n768), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(G75));
  XOR2_X1   g717(.A(new_n545), .B(KEYINPUT55), .Z(new_n904));
  AOI21_X1  g718(.A(new_n265), .B1(new_n874), .B2(new_n886), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT118), .B1(new_n905), .B2(G210), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n537), .B(KEYINPUT117), .Z(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n906), .B2(new_n907), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n907), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n908), .ZN(new_n914));
  INV_X1    g728(.A(new_n904), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n388), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n912), .A2(new_n917), .A3(new_n919), .ZN(G51));
  INV_X1    g734(.A(new_n890), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n922), .A3(new_n888), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n874), .A2(new_n886), .A3(KEYINPUT119), .A4(new_n887), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n753), .B(KEYINPUT57), .Z(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n332), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n905), .A2(G469), .A3(new_n782), .A4(new_n783), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n918), .B1(new_n927), .B2(new_n928), .ZN(G54));
  NAND3_X1  g743(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n458), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n458), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n918), .ZN(G60));
  NAND3_X1  g747(.A1(new_n921), .A2(KEYINPUT115), .A3(new_n888), .ZN(new_n934));
  INV_X1    g748(.A(new_n892), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n597), .B(KEYINPUT59), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n594), .A3(new_n593), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n593), .A2(new_n594), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n923), .A2(new_n939), .A3(new_n924), .A4(new_n936), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n938), .A2(new_n919), .A3(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(new_n874), .A2(new_n886), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n395), .A2(new_n265), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n407), .A2(new_n408), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n918), .B1(new_n946), .B2(new_n612), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n951), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n949), .A2(new_n950), .A3(new_n953), .A4(new_n954), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  INV_X1    g772(.A(G224), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n560), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n881), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n909), .B1(G898), .B2(new_n388), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  OAI21_X1  g777(.A(G953), .B1(new_n323), .B2(new_n634), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n965));
  NAND2_X1  g779(.A1(G900), .A2(G953), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n229), .A2(new_n235), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n431), .A2(new_n432), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n790), .A2(new_n282), .A3(new_n710), .A4(new_n729), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n792), .A2(new_n970), .A3(new_n800), .ZN(new_n971));
  INV_X1    g785(.A(new_n859), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n762), .A2(new_n765), .A3(new_n972), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n966), .B(new_n969), .C1(new_n974), .C2(G953), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n673), .A2(new_n683), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n845), .B1(new_n582), .B2(new_n598), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n693), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n979), .A2(new_n653), .A3(new_n652), .A4(new_n776), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n792), .A2(new_n800), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n673), .A2(new_n683), .A3(new_n982), .A4(new_n972), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n977), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT123), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT123), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n977), .A2(new_n981), .A3(new_n986), .A4(new_n983), .ZN(new_n987));
  AOI21_X1  g801(.A(G953), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n969), .B(KEYINPUT122), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n965), .B(new_n975), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(G72));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n985), .A2(new_n881), .A3(new_n987), .ZN(new_n994));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n993), .B1(new_n997), .B2(new_n659), .ZN(new_n998));
  INV_X1    g812(.A(new_n659), .ZN(new_n999));
  AOI211_X1 g813(.A(KEYINPUT125), .B(new_n999), .C1(new_n994), .C2(new_n996), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n942), .A2(new_n275), .A3(new_n999), .A4(new_n996), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n275), .B(KEYINPUT126), .Z(new_n1002));
  INV_X1    g816(.A(new_n881), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n971), .A2(new_n1003), .A3(new_n973), .ZN(new_n1004));
  INV_X1    g818(.A(new_n996), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1006), .A2(KEYINPUT127), .A3(new_n919), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT127), .B1(new_n1006), .B2(new_n919), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1001), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n998), .A2(new_n1000), .A3(new_n1009), .ZN(G57));
endmodule


