//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  AOI21_X1  g003(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n190));
  OAI21_X1  g004(.A(G131), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n190), .ZN(new_n192));
  INV_X1    g006(.A(G131), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(new_n188), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  OR2_X1    g009(.A1(new_n195), .A2(KEYINPUT17), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT75), .B(G125), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT16), .ZN(new_n201));
  OR3_X1    g015(.A1(new_n199), .A2(KEYINPUT16), .A3(G140), .ZN(new_n202));
  AOI21_X1  g016(.A(G146), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(G146), .A3(new_n202), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT17), .B(G131), .C1(new_n189), .C2(new_n190), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n196), .A2(new_n204), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT91), .B1(new_n200), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n208), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT91), .ZN(new_n212));
  OR2_X1    g026(.A1(KEYINPUT75), .A2(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT75), .A2(G125), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n197), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n212), .B(G146), .C1(new_n215), .C2(new_n198), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n209), .A2(new_n211), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT90), .A2(KEYINPUT18), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n191), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n192), .B(new_n188), .C1(new_n193), .C2(new_n218), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n207), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G113), .B(G122), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n207), .A2(new_n225), .A3(new_n221), .ZN(new_n228));
  AOI21_X1  g042(.A(G902), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G475), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT20), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT19), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n210), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n208), .B(new_n235), .C1(new_n200), .C2(new_n234), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n205), .A2(new_n195), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n221), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT92), .B1(new_n238), .B2(new_n226), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT92), .ZN(new_n240));
  AOI211_X1 g054(.A(new_n240), .B(new_n225), .C1(new_n221), .C2(new_n237), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(G475), .B1(new_n242), .B2(new_n228), .ZN(new_n243));
  INV_X1    g057(.A(G902), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n233), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n226), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n240), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n238), .A2(KEYINPUT92), .A3(new_n226), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n228), .A3(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(new_n233), .A3(new_n230), .A4(new_n244), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n232), .B1(new_n245), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n230), .A3(new_n244), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT20), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n250), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT93), .A3(new_n232), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G107), .ZN(new_n260));
  INV_X1    g074(.A(G122), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G116), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n262), .B2(KEYINPUT14), .ZN(new_n263));
  XNOR2_X1  g077(.A(G116), .B(G122), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G128), .B(G143), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT13), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n270), .B(G134), .C1(new_n271), .C2(G128), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n266), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n266), .B(G134), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n273), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT94), .B(G107), .Z(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(new_n264), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n269), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT9), .B(G234), .Z(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G217), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n281), .A2(new_n282), .A3(G953), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n279), .B(new_n283), .Z(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n244), .ZN(new_n285));
  INV_X1    g099(.A(G478), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n286), .A2(KEYINPUT15), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n285), .B(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n259), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT3), .B1(new_n224), .B2(G107), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(new_n260), .A3(G104), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n224), .A2(G107), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT82), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(G101), .ZN(new_n297));
  INV_X1    g111(.A(G101), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n291), .A2(new_n293), .A3(new_n298), .A4(new_n294), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT4), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT4), .A4(G101), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n208), .A2(G143), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n271), .A2(G146), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT0), .A4(G128), .ZN(new_n306));
  XNOR2_X1  g120(.A(G143), .B(G146), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT0), .B(G128), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g125(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n304), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n307), .B1(new_n314), .B2(G128), .ZN(new_n315));
  AND2_X1   g129(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n316));
  NOR2_X1   g130(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n317));
  OAI21_X1  g131(.A(G128), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n304), .A2(new_n305), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT67), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n312), .A2(new_n313), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n307), .A3(G128), .ZN(new_n324));
  INV_X1    g138(.A(G128), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n316), .A2(new_n317), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(new_n304), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n322), .B(new_n324), .C1(new_n327), .C2(new_n307), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n260), .A2(G104), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n224), .A2(G107), .ZN(new_n331));
  OAI21_X1  g145(.A(G101), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n299), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n299), .A2(new_n332), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT1), .B1(new_n271), .B2(G146), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT83), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n304), .A2(new_n338), .A3(KEYINPUT1), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(G128), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n319), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n335), .B1(new_n341), .B2(new_n324), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n342), .A2(KEYINPUT84), .A3(KEYINPUT10), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n325), .B1(new_n336), .B2(KEYINPUT83), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n307), .B1(new_n345), .B2(new_n339), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n333), .B1(new_n346), .B2(new_n320), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n311), .B(new_n334), .C1(new_n343), .C2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT11), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n267), .B2(G137), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n267), .A2(G137), .ZN(new_n353));
  INV_X1    g167(.A(G137), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT11), .A3(G134), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G131), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n352), .A2(new_n355), .A3(new_n193), .A4(new_n353), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT84), .B1(new_n342), .B2(KEYINPUT10), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n347), .A2(new_n344), .A3(new_n348), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n359), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n363), .A2(new_n364), .A3(new_n311), .A4(new_n334), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G110), .B(G140), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT80), .ZN(new_n368));
  INV_X1    g182(.A(G227), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G953), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n368), .B(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n314), .A2(G128), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n319), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n335), .A3(new_n324), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n364), .B1(new_n347), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT12), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n365), .A2(new_n380), .A3(new_n371), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n366), .A2(KEYINPUT86), .A3(new_n372), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G469), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n244), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n244), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n365), .A2(new_n371), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT85), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT85), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n365), .A2(new_n390), .A3(new_n371), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n360), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n365), .A2(new_n380), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n371), .A2(KEYINPUT81), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n371), .A2(KEYINPUT81), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n392), .A2(G469), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n385), .A2(new_n387), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G221), .B1(new_n281), .B2(G902), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g215(.A(G110), .B(G122), .Z(new_n402));
  XOR2_X1   g216(.A(KEYINPUT2), .B(G113), .Z(new_n403));
  INV_X1    g217(.A(G119), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G116), .ZN(new_n405));
  INV_X1    g219(.A(G116), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G119), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT66), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n407), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT2), .B(G113), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT66), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n301), .B2(new_n302), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT5), .ZN(new_n417));
  OAI21_X1  g231(.A(G113), .B1(new_n405), .B2(KEYINPUT5), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n408), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(new_n335), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n402), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n413), .A2(new_n414), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n422), .B2(new_n303), .ZN(new_n423));
  INV_X1    g237(.A(new_n402), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT6), .ZN(new_n426));
  OR3_X1    g240(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n424), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n199), .B1(new_n315), .B2(new_n320), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n199), .B2(new_n309), .ZN(new_n429));
  INV_X1    g243(.A(G953), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G224), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n426), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n418), .B(KEYINPUT88), .Z(new_n434));
  OAI21_X1  g248(.A(new_n408), .B1(new_n434), .B2(new_n417), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n333), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n419), .A2(new_n333), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT8), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(new_n424), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n436), .B(new_n439), .C1(new_n438), .C2(new_n424), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n431), .A2(KEYINPUT7), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n429), .B(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n442), .A3(new_n425), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n433), .A2(new_n244), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(KEYINPUT89), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n446), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n433), .A2(new_n244), .A3(new_n448), .A4(new_n443), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n430), .A2(G952), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(G234), .B2(G237), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(G898), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT95), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI211_X1 g269(.A(new_n244), .B(new_n430), .C1(G234), .C2(G237), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n452), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n459), .B(KEYINPUT87), .Z(new_n460));
  NAND3_X1  g274(.A1(new_n450), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n290), .A2(new_n401), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT96), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n404), .A2(G128), .ZN(new_n467));
  NAND2_X1  g281(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G110), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n325), .A2(G119), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n404), .A2(G128), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n471), .A2(new_n472), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT76), .ZN(new_n477));
  INV_X1    g291(.A(new_n475), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT74), .B(KEYINPUT23), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n479), .B2(new_n467), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT76), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n472), .A4(new_n474), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT73), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT73), .B1(new_n404), .B2(G128), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n473), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT24), .B(G110), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n477), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n211), .A3(new_n205), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT77), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n480), .A2(new_n474), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G110), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n486), .A2(new_n487), .ZN(new_n494));
  INV_X1    g308(.A(new_n205), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n493), .B(new_n494), .C1(new_n495), .C2(new_n203), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT77), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n489), .A2(new_n497), .A3(new_n211), .A4(new_n205), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n430), .A2(G221), .A3(G234), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT78), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT22), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(G137), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n503), .B(new_n354), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n506), .A2(new_n496), .A3(new_n491), .A4(new_n498), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT79), .B(KEYINPUT25), .C1(new_n508), .C2(G902), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n282), .B1(G234), .B2(new_n244), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n505), .B2(new_n507), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT79), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n509), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n508), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n510), .A2(G902), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT64), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n267), .B2(G137), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n354), .A2(KEYINPUT64), .A3(G134), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n353), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G131), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n358), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n321), .B2(new_n328), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n309), .B1(new_n357), .B2(new_n358), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n526), .A2(new_n422), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(KEYINPUT28), .ZN(new_n529));
  INV_X1    g343(.A(new_n525), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n329), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n415), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n310), .A2(new_n359), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n524), .B(new_n358), .C1(new_n315), .C2(new_n320), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n422), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT69), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT69), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n538), .A3(new_n422), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n532), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n529), .B1(new_n540), .B2(KEYINPUT28), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n187), .A2(G210), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT27), .Z(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT26), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(new_n298), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n322), .B1(new_n377), .B2(new_n324), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n315), .A2(new_n320), .A3(KEYINPUT67), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n530), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT30), .A3(new_n533), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT30), .B1(new_n533), .B2(new_n534), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n553), .A3(new_n422), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT68), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT68), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n551), .A2(new_n553), .A3(new_n556), .A4(new_n422), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n555), .A2(new_n532), .A3(new_n545), .A4(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT31), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n547), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G472), .A2(G902), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT70), .Z(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(KEYINPUT32), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT32), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n552), .B1(new_n531), .B2(KEYINPUT30), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n556), .B1(new_n568), .B2(new_n422), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT30), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n526), .A2(new_n570), .A3(new_n527), .ZN(new_n571));
  NOR4_X1   g385(.A1(new_n571), .A2(KEYINPUT68), .A3(new_n415), .A4(new_n552), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n573), .A2(KEYINPUT31), .A3(new_n532), .A4(new_n545), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n558), .A2(new_n559), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n546), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n567), .B1(new_n576), .B2(new_n564), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n566), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n422), .B1(new_n526), .B2(new_n527), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n532), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n529), .B1(new_n580), .B2(KEYINPUT28), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n581), .A2(KEYINPUT71), .A3(KEYINPUT29), .A4(new_n545), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n415), .B1(new_n550), .B2(new_n533), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT28), .B1(new_n583), .B2(new_n528), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT28), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n532), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n584), .A2(KEYINPUT29), .A3(new_n586), .A4(new_n545), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT71), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n582), .A2(new_n589), .A3(new_n244), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT72), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT29), .B1(new_n541), .B2(new_n545), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n569), .A2(new_n572), .A3(new_n528), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n592), .B1(new_n545), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT72), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n582), .A2(new_n589), .A3(new_n595), .A4(new_n244), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n591), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G472), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n519), .B1(new_n578), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n465), .A2(new_n466), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT97), .B(G101), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G3));
  NAND2_X1  g416(.A1(new_n562), .A2(new_n244), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT98), .ZN(new_n604));
  OR3_X1    g418(.A1(new_n576), .A2(KEYINPUT98), .A3(G902), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(G472), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n562), .A2(new_n565), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n609));
  INV_X1    g423(.A(new_n519), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n608), .A2(new_n609), .A3(new_n401), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n401), .A2(new_n606), .A3(new_n607), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT99), .B1(new_n612), .B2(new_n519), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n284), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n279), .B(new_n283), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT33), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n616), .A2(G478), .A3(new_n244), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT100), .B(G478), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n285), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n259), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n444), .A2(new_n445), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n444), .A2(new_n445), .ZN(new_n625));
  INV_X1    g439(.A(new_n459), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n458), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n614), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n231), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n256), .A2(KEYINPUT101), .A3(new_n250), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n250), .A2(KEYINPUT101), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n289), .A4(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n628), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n614), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT103), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT35), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n260), .ZN(G9));
  INV_X1    g456(.A(KEYINPUT36), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n504), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT104), .Z(new_n645));
  INV_X1    g459(.A(new_n499), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n644), .B(KEYINPUT104), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n499), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n649), .A3(new_n517), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n515), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n465), .A2(new_n466), .A3(new_n608), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT37), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n472), .ZN(G12));
  AND3_X1   g468(.A1(new_n399), .A2(new_n400), .A3(new_n627), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n598), .A2(new_n577), .A3(new_n566), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n452), .B1(new_n456), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n637), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n655), .A2(new_n656), .A3(new_n651), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT105), .ZN(new_n661));
  INV_X1    g475(.A(new_n651), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n578), .B2(new_n598), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n659), .A4(new_n655), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  AND3_X1   g481(.A1(new_n447), .A2(KEYINPUT38), .A3(new_n449), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT38), .B1(new_n447), .B2(new_n449), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n259), .A2(new_n459), .A3(new_n289), .A4(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n658), .B(KEYINPUT39), .Z(new_n672));
  AND2_X1   g486(.A1(new_n401), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n555), .A2(new_n532), .A3(new_n557), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n545), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n244), .B1(new_n545), .B2(new_n580), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n566), .A2(new_n577), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n662), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n675), .B(new_n683), .C1(new_n674), .C2(new_n673), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  INV_X1    g499(.A(new_n658), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT93), .B1(new_n257), .B2(new_n232), .ZN(new_n687));
  AOI211_X1 g501(.A(new_n253), .B(new_n231), .C1(new_n256), .C2(new_n250), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n622), .B(new_n686), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n663), .A2(new_n655), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  AOI21_X1  g506(.A(KEYINPUT86), .B1(new_n366), .B2(new_n372), .ZN(new_n693));
  AOI211_X1 g507(.A(new_n374), .B(new_n371), .C1(new_n360), .C2(new_n365), .ZN(new_n694));
  INV_X1    g508(.A(new_n381), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(KEYINPUT106), .A2(G469), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n696), .A2(G902), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n697), .B1(new_n383), .B2(new_n244), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n400), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n599), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n629), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT107), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(G15));
  NAND3_X1  g522(.A1(new_n599), .A2(new_n703), .A3(new_n638), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  NAND3_X1  g524(.A1(new_n663), .A2(new_n458), .A3(new_n627), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n703), .A2(new_n290), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n404), .ZN(G21));
  OAI211_X1 g528(.A(new_n289), .B(new_n627), .C1(new_n687), .C2(new_n688), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n259), .A2(KEYINPUT108), .A3(new_n289), .A4(new_n627), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n576), .B2(G902), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n581), .A2(new_n545), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n560), .B2(new_n561), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n565), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n610), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n702), .A2(new_n457), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NAND3_X1  g542(.A1(new_n720), .A2(new_n651), .A3(new_n723), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT109), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n720), .A2(new_n651), .A3(new_n723), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n701), .A2(new_n400), .A3(new_n627), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n690), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  AOI21_X1  g550(.A(new_n395), .B1(new_n365), .B2(new_n380), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n394), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n738), .B1(new_n737), .B2(new_n394), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n392), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n385), .B(new_n387), .C1(new_n741), .C2(new_n384), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n400), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n450), .A2(new_n626), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n599), .A3(new_n690), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  NAND3_X1  g564(.A1(new_n746), .A2(new_n599), .A3(new_n659), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NAND2_X1  g566(.A1(new_n622), .A2(KEYINPUT114), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n619), .A2(new_n754), .A3(new_n621), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n687), .A2(new_n688), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT115), .B1(new_n757), .B2(KEYINPUT43), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n254), .A2(KEYINPUT43), .A3(new_n258), .A4(new_n622), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n760), .B(new_n761), .C1(new_n259), .C2(new_n756), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n608), .A2(new_n662), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n385), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n392), .A2(new_n397), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g588(.A(KEYINPUT45), .B(new_n392), .C1(new_n739), .C2(new_n740), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(G469), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(KEYINPUT46), .A3(new_n387), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n771), .B1(new_n777), .B2(KEYINPUT111), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n384), .B1(new_n772), .B2(new_n773), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n386), .B1(new_n779), .B2(new_n775), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT46), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n780), .B2(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n776), .A2(new_n387), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(KEYINPUT112), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n778), .A2(new_n782), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n400), .A3(new_n672), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT113), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n768), .A2(new_n769), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n770), .A2(new_n744), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n788), .A2(new_n794), .A3(new_n400), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n794), .B1(new_n788), .B2(new_n400), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n656), .A2(new_n610), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n690), .A3(new_n744), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n801));
  NOR2_X1   g615(.A1(G952), .A2(G953), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n689), .B1(new_n730), .B2(new_n732), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n746), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n597), .A2(G472), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n566), .A2(new_n577), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n651), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n808), .A2(new_n289), .A3(new_n658), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n401), .A3(new_n810), .A4(new_n744), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n749), .A2(new_n805), .A3(new_n751), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n725), .A2(new_n726), .B1(new_n704), .B2(new_n629), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n259), .A2(KEYINPUT117), .A3(new_n288), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT117), .B1(new_n259), .B2(new_n288), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n623), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n611), .A2(new_n613), .A3(new_n462), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n709), .B1(new_n711), .B2(new_n712), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n813), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n652), .A2(new_n600), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n812), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n743), .A2(new_n658), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n719), .A2(new_n683), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT118), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n399), .A2(new_n400), .A3(new_n627), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n808), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n827), .A2(new_n690), .B1(new_n804), .B2(new_n734), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n682), .B1(new_n717), .B2(new_n718), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n830), .A3(new_n823), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n666), .A2(new_n825), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n735), .A2(new_n691), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n665), .B2(new_n661), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n830), .A2(new_n719), .A3(new_n683), .A4(new_n823), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n830), .B1(new_n829), .B2(new_n823), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n835), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n833), .A2(new_n840), .A3(KEYINPUT119), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT119), .B1(new_n833), .B2(new_n840), .ZN(new_n842));
  OAI211_X1 g656(.A(KEYINPUT53), .B(new_n822), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n749), .A2(new_n751), .A3(new_n805), .A4(new_n811), .ZN(new_n845));
  INV_X1    g659(.A(new_n820), .ZN(new_n846));
  INV_X1    g660(.A(new_n821), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n833), .A2(new_n840), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n803), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n844), .B(new_n822), .C1(new_n841), .C2(new_n842), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT53), .B1(new_n848), .B2(new_n849), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT54), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n763), .A2(new_n452), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n724), .ZN(new_n857));
  INV_X1    g671(.A(new_n734), .ZN(new_n858));
  OAI211_X1 g672(.A(G952), .B(new_n430), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n702), .A2(new_n745), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n856), .A2(new_n599), .A3(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(KEYINPUT48), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(KEYINPUT48), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n681), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n860), .A2(new_n452), .A3(new_n610), .A4(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(new_n623), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n857), .A2(new_n745), .ZN(new_n868));
  INV_X1    g682(.A(new_n701), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n400), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n797), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT51), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n856), .A2(new_n733), .A3(new_n860), .ZN(new_n873));
  OR3_X1    g687(.A1(new_n866), .A2(new_n259), .A3(new_n622), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n698), .B1(new_n696), .B2(G902), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n383), .A2(new_n244), .A3(new_n697), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n626), .A3(new_n400), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n670), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n701), .A2(KEYINPUT121), .A3(new_n626), .A4(new_n400), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n763), .A2(new_n883), .A3(new_n452), .A4(new_n724), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT50), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n876), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n864), .B(new_n867), .C1(new_n872), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n886), .B2(new_n887), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n856), .A2(KEYINPUT50), .A3(new_n724), .A4(new_n883), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n884), .A2(new_n885), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(KEYINPUT122), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n795), .B2(new_n796), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n777), .A2(KEYINPUT111), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(new_n385), .A3(new_n782), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n787), .A2(new_n784), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n400), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT47), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n788), .A2(new_n794), .A3(new_n400), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(KEYINPUT120), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n870), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n897), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n868), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n895), .A2(new_n876), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT51), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT123), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n908), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n889), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n802), .B1(new_n855), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n610), .A2(new_n400), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n259), .B(new_n916), .C1(new_n621), .C2(new_n619), .ZN(new_n917));
  INV_X1    g731(.A(new_n670), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n918), .A2(new_n460), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n701), .B(KEYINPUT49), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n917), .A2(new_n865), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n801), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n889), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n875), .B1(new_n891), .B2(new_n894), .ZN(new_n925));
  AOI211_X1 g739(.A(KEYINPUT123), .B(KEYINPUT51), .C1(new_n925), .C2(new_n907), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n912), .B1(new_n908), .B2(new_n909), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n928), .A2(new_n851), .A3(new_n854), .ZN(new_n929));
  OAI211_X1 g743(.A(KEYINPUT124), .B(new_n921), .C1(new_n929), .C2(new_n802), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n923), .A2(new_n930), .ZN(G75));
  AND2_X1   g745(.A1(new_n852), .A2(new_n853), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(G210), .A3(G902), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n426), .A2(new_n427), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n432), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n933), .B2(new_n934), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n430), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  AND2_X1   g755(.A1(new_n932), .A2(G902), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n775), .A3(new_n779), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n386), .B(KEYINPUT57), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n852), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(new_n854), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n383), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n943), .B2(new_n947), .ZN(G54));
  NAND4_X1  g762(.A1(new_n942), .A2(KEYINPUT58), .A3(G475), .A4(new_n249), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n932), .A2(KEYINPUT58), .A3(G902), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n228), .B(new_n242), .C1(new_n950), .C2(new_n230), .ZN(new_n951));
  INV_X1    g765(.A(new_n940), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(G60));
  NAND2_X1  g767(.A1(new_n616), .A2(new_n618), .ZN(new_n954));
  XNOR2_X1  g768(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n286), .A2(new_n244), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n954), .B1(new_n855), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n954), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n960), .B(new_n957), .C1(new_n945), .C2(new_n854), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n959), .A2(new_n952), .A3(new_n961), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  AOI21_X1  g778(.A(new_n516), .B1(new_n932), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n647), .A2(new_n649), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n852), .A2(new_n853), .A3(new_n966), .A4(new_n964), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n952), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n967), .A2(KEYINPUT126), .A3(new_n952), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(KEYINPUT61), .B(new_n970), .C1(new_n965), .C2(new_n968), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G66));
  AOI21_X1  g788(.A(new_n430), .B1(new_n454), .B2(G224), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n846), .A2(new_n847), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n430), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n935), .B1(G898), .B2(new_n430), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT127), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n977), .B(new_n979), .ZN(G69));
  AND2_X1   g794(.A1(new_n792), .A2(new_n799), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n790), .A2(new_n599), .A3(new_n719), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n835), .A2(new_n749), .A3(new_n751), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n984), .A2(G953), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n235), .B1(new_n200), .B2(new_n234), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n568), .B(new_n986), .Z(new_n987));
  AND2_X1   g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n657), .B2(G227), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n816), .A2(new_n599), .A3(new_n673), .A4(new_n744), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n835), .A2(new_n684), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT62), .Z(new_n992));
  NAND3_X1  g806(.A1(new_n981), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n987), .B1(new_n993), .B2(new_n430), .ZN(new_n994));
  OAI21_X1  g808(.A(G953), .B1(new_n369), .B2(new_n657), .ZN(new_n995));
  AOI22_X1  g809(.A1(new_n988), .A2(new_n989), .B1(new_n994), .B2(new_n995), .ZN(G72));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n993), .B2(new_n976), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n940), .B1(new_n999), .B2(new_n678), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n998), .B1(new_n984), .B2(new_n976), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n676), .A2(new_n545), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n678), .B(new_n1002), .C1(new_n843), .C2(new_n850), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n998), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n1000), .A2(new_n1003), .A3(new_n1005), .ZN(G57));
endmodule


