//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(G1gat), .B2(new_n203), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n207), .B(new_n208), .Z(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  OR3_X1    g009(.A1(new_n210), .A2(KEYINPUT88), .A3(KEYINPUT15), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n213));
  XOR2_X1   g012(.A(KEYINPUT14), .B(G29gat), .Z(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(G36gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT15), .B1(new_n210), .B2(KEYINPUT88), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT89), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n222), .A2(KEYINPUT17), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(KEYINPUT17), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n209), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT91), .ZN(new_n227));
  INV_X1    g026(.A(new_n222), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(new_n209), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n225), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT18), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n222), .B(new_n209), .Z(new_n233));
  XOR2_X1   g032(.A(new_n227), .B(KEYINPUT13), .Z(new_n234));
  AOI22_X1  g033(.A1(new_n231), .A2(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT11), .B(G169gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n222), .B(KEYINPUT17), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n229), .B1(new_n242), .B2(new_n209), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT18), .A3(new_n227), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n235), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n241), .B1(new_n235), .B2(new_n244), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G8gat), .B(G36gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(G64gat), .B(G92gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G211gat), .A2(G218gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(G211gat), .A2(G218gat), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT74), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT73), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT22), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(G197gat), .A2(G204gat), .ZN(new_n259));
  AND2_X1   g058(.A1(G197gat), .A2(G204gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n256), .B1(new_n252), .B2(new_n257), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n254), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n252), .ZN(new_n266));
  INV_X1    g065(.A(new_n262), .ZN(new_n267));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .A4(new_n258), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G226gat), .A2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT26), .ZN(new_n275));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(G169gat), .B2(G176gat), .ZN(new_n278));
  AND2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n275), .B(new_n276), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G183gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT27), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G183gat), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(KEYINPUT28), .A3(new_n285), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n280), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT25), .ZN(new_n292));
  AND2_X1   g091(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n293), .A2(new_n285), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  OR2_X1    g093(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(G190gat), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n294), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n274), .ZN(new_n302));
  NAND2_X1  g101(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(KEYINPUT23), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n273), .A2(KEYINPUT64), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT64), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G169gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n292), .B1(new_n300), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n292), .B1(new_n311), .B2(KEYINPUT23), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n294), .A2(new_n297), .A3(new_n299), .A4(new_n312), .ZN(new_n313));
  AOI211_X1 g112(.A(KEYINPUT76), .B(new_n291), .C1(new_n310), .C2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(new_n313), .ZN(new_n316));
  INV_X1    g115(.A(new_n280), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT28), .B1(new_n289), .B2(new_n285), .ZN(new_n318));
  AND4_X1   g117(.A1(KEYINPUT28), .A2(new_n282), .A3(new_n284), .A4(new_n285), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n315), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(KEYINPUT66), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n291), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n316), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n272), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n272), .A2(new_n322), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g129(.A1(new_n328), .A2(new_n329), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n270), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n270), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n322), .A2(new_n327), .A3(new_n271), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n326), .A2(new_n271), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n251), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n328), .A2(new_n329), .ZN(new_n338));
  INV_X1    g137(.A(new_n321), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n316), .A2(new_n315), .A3(new_n320), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n272), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n328), .A2(new_n329), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n333), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n271), .A2(new_n327), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n335), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n270), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n348), .A3(new_n250), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n332), .A2(new_n336), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n250), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n355));
  INV_X1    g154(.A(G134gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G127gat), .ZN(new_n357));
  INV_X1    g156(.A(G127gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G134gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT67), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G113gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G120gat), .ZN(new_n365));
  INV_X1    g164(.A(G120gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G113gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT1), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n355), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n367), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT1), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n372), .A2(KEYINPUT68), .A3(new_n361), .A4(new_n362), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n366), .A2(KEYINPUT69), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT69), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G120gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n377), .A3(G113gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n365), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(KEYINPUT70), .A3(new_n365), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n357), .A2(new_n359), .A3(new_n371), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G148gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G141gat), .ZN(new_n386));
  INV_X1    g185(.A(G141gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G148gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G155gat), .B(G162gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT2), .ZN(new_n392));
  AND4_X1   g191(.A1(KEYINPUT77), .A2(new_n389), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n386), .B2(new_n388), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n390), .B1(new_n395), .B2(new_n392), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n374), .A2(new_n384), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT78), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n374), .A2(new_n384), .A3(new_n397), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n374), .A2(new_n384), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n387), .A2(G148gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n385), .A2(G141gat), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT77), .B(new_n392), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n390), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n395), .A2(new_n390), .A3(new_n392), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n399), .A2(new_n401), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n354), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n415), .A3(new_n401), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n409), .A2(KEYINPUT3), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT3), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n407), .A2(new_n418), .A3(new_n408), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n413), .B1(new_n420), .B2(new_n402), .ZN(new_n421));
  INV_X1    g220(.A(new_n398), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT4), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n416), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n414), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n399), .A2(new_n401), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT4), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n422), .A2(KEYINPUT4), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n427), .A2(new_n429), .A3(new_n354), .A4(new_n421), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G1gat), .B(G29gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT0), .ZN(new_n433));
  XNOR2_X1  g232(.A(G57gat), .B(G85gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n431), .A2(KEYINPUT83), .A3(new_n436), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n350), .A2(new_n353), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT84), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT40), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n428), .B1(new_n426), .B2(KEYINPUT4), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n420), .A2(new_n402), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n412), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT39), .B1(new_n411), .B2(new_n413), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n436), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n449), .A2(new_n444), .A3(new_n451), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n442), .B(new_n443), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n452), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT84), .B1(new_n455), .B2(new_n441), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(G50gat), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G228gat), .A2(G233gat), .ZN(new_n462));
  OAI22_X1  g261(.A1(new_n261), .A2(new_n262), .B1(new_n253), .B2(new_n254), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n253), .A2(new_n254), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n267), .A2(new_n464), .A3(new_n268), .A4(new_n258), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n327), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n397), .B1(new_n466), .B2(new_n418), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n270), .B1(new_n327), .B2(new_n419), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n419), .A2(new_n327), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n333), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT29), .B1(new_n263), .B2(new_n269), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n409), .B1(new_n472), .B2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g272(.A(new_n462), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n461), .B1(new_n476), .B2(G22gat), .ZN(new_n477));
  INV_X1    g276(.A(G22gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n469), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT80), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n469), .A2(new_n475), .A3(KEYINPUT80), .A4(new_n478), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT81), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT81), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n477), .A2(new_n481), .A3(new_n485), .A4(new_n482), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n479), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n478), .B1(new_n469), .B2(new_n475), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n461), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n344), .A2(new_n348), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n251), .B1(new_n492), .B2(KEYINPUT37), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n351), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT38), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n270), .B1(new_n342), .B2(new_n343), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n494), .B1(new_n347), .B2(new_n333), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT38), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n499), .B(new_n251), .C1(KEYINPUT37), .C2(new_n492), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n496), .A2(new_n349), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n425), .A2(new_n430), .A3(new_n435), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n439), .A2(new_n502), .A3(new_n503), .A4(new_n440), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n431), .A2(KEYINPUT6), .A3(new_n436), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT85), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n505), .A2(KEYINPUT85), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n491), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n457), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n374), .A2(new_n384), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n326), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n402), .A2(new_n316), .A3(new_n323), .A4(new_n325), .ZN(new_n514));
  AND2_X1   g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT32), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT71), .B(KEYINPUT33), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G15gat), .B(G43gat), .Z(new_n520));
  XNOR2_X1  g319(.A(G71gat), .B(G99gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n522), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n516), .B(KEYINPUT32), .C1(new_n518), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT34), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n513), .A2(new_n514), .ZN(new_n528));
  OAI211_X1 g327(.A(KEYINPUT72), .B(new_n527), .C1(new_n528), .C2(new_n515), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n515), .B1(new_n513), .B2(new_n514), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT34), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n523), .A2(new_n532), .A3(new_n529), .A4(new_n525), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT36), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n535), .B2(new_n537), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n491), .B(KEYINPUT82), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n437), .A2(new_n502), .A3(new_n503), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n353), .A2(new_n350), .B1(new_n545), .B2(new_n505), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n543), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n511), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n350), .A2(new_n353), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n487), .A2(new_n490), .B1(new_n534), .B2(new_n536), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n552));
  NAND4_X1  g351(.A1(new_n508), .A2(new_n550), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT87), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555));
  AOI211_X1 g354(.A(new_n554), .B(new_n555), .C1(new_n546), .C2(new_n551), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n545), .A2(new_n505), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT87), .B1(new_n558), .B2(KEYINPUT35), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n553), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n247), .B1(new_n549), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562));
  AND2_X1   g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(G57gat), .A2(G64gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(G57gat), .A2(G64gat), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n567), .B(new_n568), .C1(new_n563), .C2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n566), .B(new_n569), .C1(new_n570), .C2(new_n563), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n563), .B(new_n564), .C1(new_n569), .C2(new_n570), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n562), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n569), .B1(new_n570), .B2(new_n563), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n565), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(KEYINPUT93), .A3(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT94), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT95), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G183gat), .B(G211gat), .Z(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  OAI21_X1  g386(.A(new_n209), .B1(new_n579), .B2(new_n580), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT96), .ZN(new_n589));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n589), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n587), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT7), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n602), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n600), .A2(new_n605), .A3(new_n609), .A4(new_n601), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n242), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT99), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n242), .A2(new_n615), .A3(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n608), .A2(new_n610), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n228), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G190gat), .B(G218gat), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n624), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n617), .A2(new_n629), .A3(new_n622), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n628), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n629), .B1(new_n617), .B2(new_n622), .ZN(new_n633));
  AOI211_X1 g432(.A(new_n624), .B(new_n621), .C1(new_n614), .C2(new_n616), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n597), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  AOI21_X1  g439(.A(new_n611), .B1(new_n574), .B2(new_n577), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n620), .A2(new_n572), .A3(new_n573), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT100), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n640), .B1(new_n646), .B2(KEYINPUT101), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(KEYINPUT101), .B2(new_n646), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n641), .B2(new_n642), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n645), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n640), .ZN(new_n655));
  INV_X1    g454(.A(new_n646), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n655), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n637), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n561), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n557), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n660), .A2(new_n550), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n202), .B2(new_n665), .ZN(new_n668));
  MUX2_X1   g467(.A(new_n667), .B(new_n668), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g468(.A(new_n538), .ZN(new_n670));
  AOI21_X1  g469(.A(G15gat), .B1(new_n661), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n542), .A2(G15gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT102), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n661), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n660), .A2(new_n544), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NOR2_X1   g476(.A1(new_n597), .A2(new_n658), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n636), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n561), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(G29gat), .A3(new_n557), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT45), .Z(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n560), .A2(KEYINPUT103), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n686), .B(new_n553), .C1(new_n556), .C2(new_n559), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n685), .A2(new_n687), .B1(new_n511), .B2(new_n548), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n688), .B2(new_n636), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n549), .A2(new_n560), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n631), .A2(new_n635), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(KEYINPUT44), .A3(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n679), .A2(new_n247), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n557), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n683), .A2(new_n696), .ZN(G1328gat));
  OAI21_X1  g496(.A(G36gat), .B1(new_n695), .B2(new_n550), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n681), .A2(G36gat), .A3(new_n550), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1329gat));
  NOR3_X1   g500(.A1(new_n681), .A2(G43gat), .A3(new_n538), .ZN(new_n702));
  INV_X1    g501(.A(new_n695), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n542), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n704), .B2(G43gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g505(.A(new_n491), .ZN(new_n707));
  OAI21_X1  g506(.A(G50gat), .B1(new_n695), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n681), .A2(G50gat), .A3(new_n544), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT48), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n709), .B1(new_n708), .B2(new_n712), .ZN(new_n714));
  INV_X1    g513(.A(new_n544), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n703), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n710), .B1(new_n716), .B2(G50gat), .ZN(new_n717));
  OAI22_X1  g516(.A1(new_n713), .A2(new_n714), .B1(new_n717), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g517(.A1(new_n558), .A2(KEYINPUT35), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n554), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n558), .A2(KEYINPUT87), .A3(KEYINPUT35), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n686), .B1(new_n722), .B2(new_n553), .ZN(new_n723));
  INV_X1    g522(.A(new_n687), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n549), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n245), .A2(new_n246), .ZN(new_n726));
  INV_X1    g525(.A(new_n658), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n637), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n662), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g531(.A1(new_n729), .A2(new_n550), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  AND2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n733), .B2(new_n734), .ZN(G1333gat));
  NAND3_X1  g536(.A1(new_n730), .A2(G71gat), .A3(new_n542), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n538), .B(KEYINPUT105), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n729), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(G71gat), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n730), .A2(new_n715), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g543(.A1(new_n597), .A2(new_n726), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n725), .A2(KEYINPUT51), .A3(new_n691), .A4(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n685), .A2(new_n687), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n636), .B1(new_n751), .B2(new_n549), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT51), .B1(new_n752), .B2(new_n745), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n753), .A2(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(KEYINPUT108), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n662), .A2(new_n603), .A3(new_n658), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n597), .A2(new_n726), .A3(new_n727), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n689), .A2(new_n692), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT106), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n689), .A2(new_n761), .A3(new_n692), .A4(new_n758), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n760), .A2(new_n662), .A3(new_n762), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n756), .A2(new_n757), .B1(new_n603), .B2(new_n763), .ZN(G1336gat));
  INV_X1    g563(.A(new_n550), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n760), .A2(new_n765), .A3(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G92gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n727), .A2(new_n550), .A3(G92gat), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n725), .A2(new_n691), .A3(new_n745), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n770), .A2(KEYINPUT109), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT109), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n746), .B(new_n747), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n769), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n767), .B1(new_n776), .B2(KEYINPUT110), .ZN(new_n777));
  INV_X1    g576(.A(new_n773), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n753), .A2(KEYINPUT109), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n778), .B(new_n779), .C1(new_n748), .C2(new_n749), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n780), .A2(KEYINPUT110), .A3(new_n768), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT52), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G92gat), .B1(new_n759), .B2(new_n550), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n784));
  OAI211_X1 g583(.A(new_n783), .B(new_n784), .C1(new_n756), .C2(new_n769), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1337gat));
  XNOR2_X1  g585(.A(KEYINPUT112), .B(G99gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n670), .A2(new_n658), .A3(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n760), .A2(new_n542), .A3(new_n762), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n756), .A2(new_n788), .B1(new_n789), .B2(new_n787), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n693), .A2(new_n491), .A3(new_n758), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n707), .A2(new_n727), .A3(G106gat), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n794), .A2(new_n795), .B1(new_n756), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n760), .A2(new_n715), .A3(new_n762), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n799), .B1(new_n780), .B2(new_n796), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n798), .A2(new_n799), .B1(new_n801), .B2(new_n802), .ZN(G1339gat));
  INV_X1    g602(.A(new_n597), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n650), .A2(new_n645), .A3(new_n651), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n650), .A2(KEYINPUT114), .A3(new_n645), .A4(new_n651), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n807), .A2(new_n653), .A3(KEYINPUT54), .A4(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n640), .B1(new_n652), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n809), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT55), .B1(new_n809), .B2(new_n811), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n653), .B2(new_n648), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n726), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n235), .A2(new_n241), .A3(new_n244), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n243), .A2(new_n227), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n233), .A2(new_n234), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n239), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n658), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n691), .B1(new_n820), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n816), .A2(new_n818), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n636), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n804), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n597), .A2(new_n247), .A3(new_n636), .A4(new_n727), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n557), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n551), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT116), .Z(new_n835));
  NAND4_X1  g634(.A1(new_n835), .A2(new_n364), .A3(new_n550), .A4(new_n726), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n715), .B1(new_n831), .B2(new_n832), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n662), .A2(new_n550), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n538), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n247), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(G1340gat));
  OAI21_X1  g644(.A(G120gat), .B1(new_n841), .B2(new_n727), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n835), .A2(new_n550), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n658), .A2(new_n375), .A3(new_n377), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT118), .ZN(G1341gat));
  NAND3_X1  g649(.A1(new_n840), .A2(G127gat), .A3(new_n597), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT119), .Z(new_n852));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n550), .A3(new_n597), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n358), .B2(new_n853), .ZN(G1342gat));
  NOR2_X1   g653(.A1(new_n636), .A2(new_n765), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n835), .A2(new_n356), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n841), .B2(new_n636), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G1343gat));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n707), .B1(new_n831), .B2(new_n832), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n542), .A2(new_n838), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n247), .B1(new_n829), .B2(KEYINPUT121), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n819), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n827), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT122), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n868), .A2(new_n870), .B1(new_n658), .B2(new_n826), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n873), .A2(new_n636), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n830), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n597), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n832), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n715), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n247), .B(new_n867), .C1(new_n881), .C2(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n862), .B1(new_n882), .B2(new_n387), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n542), .A2(new_n707), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n833), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n765), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n387), .A3(new_n726), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n882), .B2(new_n387), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n883), .A2(new_n888), .A3(KEYINPUT58), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  OAI221_X1 g689(.A(new_n887), .B1(new_n862), .B2(new_n890), .C1(new_n882), .C2(new_n387), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1344gat));
  NAND3_X1  g691(.A1(new_n886), .A2(new_n385), .A3(new_n658), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n866), .A2(new_n658), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n636), .B1(new_n874), .B2(new_n875), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n871), .A2(new_n875), .A3(new_n827), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n878), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n880), .B1(new_n898), .B2(new_n804), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n864), .B1(new_n899), .B2(new_n544), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n863), .A2(KEYINPUT124), .A3(KEYINPUT57), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT124), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n895), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n385), .B1(new_n904), .B2(KEYINPUT125), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n831), .A2(new_n832), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(KEYINPUT57), .A3(new_n491), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n863), .A2(KEYINPUT124), .A3(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n881), .B2(new_n864), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n906), .B1(new_n913), .B2(new_n895), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n894), .B1(new_n905), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n867), .B1(new_n881), .B2(KEYINPUT57), .ZN(new_n916));
  AOI211_X1 g715(.A(KEYINPUT59), .B(new_n385), .C1(new_n916), .C2(new_n658), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n893), .B1(new_n915), .B2(new_n917), .ZN(G1345gat));
  INV_X1    g717(.A(G155gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n886), .A2(new_n919), .A3(new_n597), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n916), .A2(new_n597), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n919), .ZN(G1346gat));
  AND2_X1   g721(.A1(new_n916), .A2(new_n691), .ZN(new_n923));
  INV_X1    g722(.A(G162gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n855), .A2(new_n924), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n923), .A2(new_n924), .B1(new_n885), .B2(new_n925), .ZN(G1347gat));
  AOI21_X1  g725(.A(new_n662), .B1(new_n831), .B2(new_n832), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n765), .A2(new_n551), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT126), .Z(new_n929));
  AND2_X1   g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n930), .A2(new_n305), .A3(new_n307), .A4(new_n726), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n765), .A2(new_n557), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n739), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n837), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n934), .A2(new_n726), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(new_n273), .ZN(G1348gat));
  AOI21_X1  g735(.A(G176gat), .B1(new_n930), .B2(new_n658), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n727), .B1(new_n302), .B2(new_n303), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n934), .B2(new_n938), .ZN(G1349gat));
  AOI21_X1  g738(.A(new_n281), .B1(new_n934), .B2(new_n597), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n597), .A2(new_n289), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n930), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g742(.A1(new_n930), .A2(new_n285), .A3(new_n691), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n934), .A2(new_n691), .ZN(new_n945));
  NOR2_X1   g744(.A1(KEYINPUT127), .A2(KEYINPUT61), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n285), .B1(KEYINPUT127), .B2(KEYINPUT61), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  AND3_X1   g749(.A1(new_n927), .A2(new_n765), .A3(new_n884), .ZN(new_n951));
  AOI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n726), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n900), .A2(new_n903), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n542), .A2(new_n932), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n726), .A2(G197gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  INV_X1    g756(.A(G204gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n951), .A2(new_n958), .A3(new_n658), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  AND2_X1   g759(.A1(new_n955), .A2(new_n658), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n958), .ZN(G1353gat));
  INV_X1    g761(.A(G211gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n951), .A2(new_n963), .A3(new_n597), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n953), .A2(new_n597), .A3(new_n954), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  INV_X1    g767(.A(G218gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n969), .A3(new_n691), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n955), .A2(new_n691), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n969), .ZN(G1355gat));
endmodule


