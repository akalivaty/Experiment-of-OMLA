//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT20), .Z(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT90), .ZN(new_n205));
  AOI21_X1  g004(.A(G1gat), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT16), .B1(new_n207), .B2(KEYINPUT90), .ZN(new_n208));
  INV_X1    g007(.A(G15gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G22gat), .ZN(new_n210));
  INV_X1    g009(.A(G22gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G15gat), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(G8gat), .B1(new_n206), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n212), .A3(new_n205), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  INV_X1    g015(.A(G8gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n204), .A2(new_n208), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(G71gat), .A2(G78gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT94), .ZN(new_n222));
  NAND2_X1  g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(G71gat), .A2(G78gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G71gat), .A2(G78gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT94), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n225), .A2(KEYINPUT9), .ZN(new_n228));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n224), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G64gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT95), .B1(new_n231), .B2(G57gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT95), .ZN(new_n233));
  INV_X1    g032(.A(G57gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(G64gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(G57gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n225), .A2(KEYINPUT9), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n230), .A2(new_n240), .A3(KEYINPUT21), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n220), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G211gat), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n230), .A2(new_n240), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT21), .ZN(new_n245));
  INV_X1    g044(.A(G211gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n220), .A2(new_n246), .A3(new_n241), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n243), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n245), .B1(new_n243), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n203), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n247), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n244), .A2(KEYINPUT21), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n243), .A2(new_n245), .A3(new_n247), .ZN(new_n254));
  INV_X1    g053(.A(new_n203), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G231gat), .A2(G233gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(KEYINPUT96), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT19), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT97), .B(G183gat), .Z(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n250), .A2(new_n256), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n250), .B2(new_n256), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G134gat), .B(G162gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(G99gat), .A2(G106gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT8), .ZN(new_n267));
  NAND2_X1  g066(.A1(G85gat), .A2(G92gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT7), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G85gat), .ZN(new_n271));
  INV_X1    g070(.A(G92gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n267), .A2(new_n270), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G99gat), .B(G106gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(KEYINPUT8), .A2(new_n266), .B1(new_n271), .B2(new_n272), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n279), .A2(new_n276), .A3(new_n270), .A4(new_n274), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G50gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G43gat), .ZN(new_n283));
  INV_X1    g082(.A(G43gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G50gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT15), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT14), .ZN(new_n288));
  INV_X1    g087(.A(G29gat), .ZN(new_n289));
  INV_X1    g088(.A(G36gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT89), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI211_X1 g093(.A(KEYINPUT89), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G29gat), .A2(G36gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n287), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT17), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT15), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n284), .A2(G50gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n282), .A2(G43gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n291), .A2(new_n293), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n296), .A4(new_n286), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n298), .A2(new_n299), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n299), .B1(new_n298), .B2(new_n305), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n281), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT98), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n298), .A2(new_n305), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n278), .A2(new_n280), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT41), .ZN(new_n315));
  INV_X1    g114(.A(G232gat), .ZN(new_n316));
  INV_X1    g115(.A(G233gat), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n311), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  AOI211_X1 g119(.A(KEYINPUT98), .B(new_n318), .C1(new_n312), .C2(new_n313), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n308), .B(new_n310), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n281), .B1(new_n298), .B2(new_n305), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT98), .B1(new_n324), .B2(new_n318), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n314), .A2(new_n311), .A3(new_n319), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n310), .B1(new_n327), .B2(new_n308), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n265), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G190gat), .B(G218gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n308), .B1(new_n320), .B2(new_n321), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n309), .ZN(new_n332));
  INV_X1    g131(.A(new_n265), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n322), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n330), .B1(new_n329), .B2(new_n334), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n264), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G197gat), .ZN(new_n339));
  INV_X1    g138(.A(G204gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G197gat), .A2(G204gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT22), .ZN(new_n343));
  NAND2_X1  g142(.A1(G211gat), .A2(G218gat), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(G211gat), .A2(G218gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G211gat), .A2(G218gat), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT70), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n349));
  INV_X1    g148(.A(G218gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n246), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n349), .B1(new_n351), .B2(new_n344), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n345), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n354));
  NOR2_X1   g153(.A1(G197gat), .A2(G204gat), .ZN(new_n355));
  AND2_X1   g154(.A1(G197gat), .A2(G204gat), .ZN(new_n356));
  OAI22_X1  g155(.A1(new_n355), .A2(new_n356), .B1(new_n346), .B2(KEYINPUT22), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT70), .B1(new_n346), .B2(new_n347), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n349), .A3(new_n344), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n353), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(KEYINPUT79), .B(new_n345), .C1(new_n348), .C2(new_n352), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367));
  INV_X1    g166(.A(G155gat), .ZN(new_n368));
  INV_X1    g167(.A(G162gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT2), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT73), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT73), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT2), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G141gat), .B(G148gat), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n367), .B(new_n370), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n368), .A3(new_n369), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n367), .ZN(new_n379));
  INV_X1    g178(.A(G148gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G141gat), .ZN(new_n381));
  INV_X1    g180(.A(G141gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G148gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n377), .A2(KEYINPUT75), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT75), .B1(new_n377), .B2(new_n385), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n353), .A2(new_n360), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n378), .A2(new_n367), .B1(new_n381), .B2(new_n383), .ZN(new_n390));
  INV_X1    g189(.A(new_n367), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT73), .B(KEYINPUT2), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n384), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n393), .B2(new_n370), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n394), .B2(new_n365), .ZN(new_n395));
  OAI22_X1  g194(.A1(new_n366), .A2(new_n388), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G228gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(new_n317), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT80), .B1(new_n395), .B2(new_n389), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n377), .A2(new_n365), .A3(new_n385), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n363), .ZN(new_n403));
  INV_X1    g202(.A(new_n389), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n377), .A2(new_n385), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT29), .B1(new_n353), .B2(new_n360), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(KEYINPUT3), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n398), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n400), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n403), .A2(new_n405), .A3(new_n404), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n405), .B1(new_n403), .B2(new_n404), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n411), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(KEYINPUT81), .A3(new_n416), .ZN(new_n417));
  AOI221_X4 g216(.A(G22gat), .B1(new_n396), .B2(new_n399), .C1(new_n412), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n412), .A2(new_n417), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n396), .A2(new_n399), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n211), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT82), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT81), .B1(new_n415), .B2(new_n416), .ZN(new_n423));
  NOR4_X1   g222(.A1(new_n411), .A2(new_n413), .A3(new_n414), .A4(new_n400), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G22gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n419), .A2(new_n211), .A3(new_n420), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT31), .B(G50gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n422), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT69), .B(G71gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(G99gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G15gat), .B(G43gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G227gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(new_n317), .ZN(new_n441));
  INV_X1    g240(.A(G190gat), .ZN(new_n442));
  AND2_X1   g241(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT28), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT27), .B(G183gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT28), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n442), .ZN(new_n449));
  OR3_X1    g248(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(G169gat), .A2(G176gat), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G183gat), .A2(G190gat), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n446), .A2(new_n449), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G134gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G127gat), .ZN(new_n457));
  INV_X1    g256(.A(G127gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G134gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G113gat), .B(G120gat), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(KEYINPUT1), .ZN(new_n462));
  INV_X1    g261(.A(G120gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(G113gat), .ZN(new_n464));
  INV_X1    g263(.A(G113gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G120gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G127gat), .B(G134gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT1), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n454), .ZN(new_n473));
  NAND3_X1  g272(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT66), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n479));
  INV_X1    g278(.A(G169gat), .ZN(new_n480));
  INV_X1    g279(.A(G176gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n451), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n486));
  INV_X1    g285(.A(new_n451), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(KEYINPUT65), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n478), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n487), .B1(new_n473), .B2(new_n474), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n482), .A2(new_n483), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n455), .B(new_n471), .C1(new_n489), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n473), .A2(new_n474), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n451), .A3(new_n493), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n490), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n478), .A2(new_n485), .A3(new_n488), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n471), .B1(new_n501), .B2(new_n455), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n441), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n441), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n455), .B1(new_n489), .B2(new_n494), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n462), .A2(new_n470), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n506), .B1(new_n509), .B2(new_n495), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT67), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n439), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n510), .A2(KEYINPUT67), .ZN(new_n516));
  AOI211_X1 g315(.A(new_n504), .B(new_n506), .C1(new_n509), .C2(new_n495), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT32), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n509), .A2(new_n506), .A3(new_n495), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT34), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT34), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n509), .A2(new_n521), .A3(new_n506), .A4(new_n495), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n512), .A2(KEYINPUT32), .A3(new_n523), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n515), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n514), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n525), .A2(new_n526), .B1(new_n528), .B2(new_n438), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n426), .A2(new_n427), .A3(new_n428), .A4(new_n432), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n434), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g332(.A1(G226gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n507), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n533), .B1(new_n507), .B2(new_n535), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n507), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n501), .A2(KEYINPUT71), .A3(new_n455), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT29), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n538), .B(new_n404), .C1(new_n535), .C2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n541), .A3(new_n535), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n507), .A2(new_n363), .A3(new_n534), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n389), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G8gat), .B(G36gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(new_n231), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(new_n272), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n543), .A2(new_n546), .A3(new_n550), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(KEYINPUT30), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n547), .A2(new_n555), .A3(new_n551), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n408), .A2(new_n508), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT4), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT78), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n559), .B(new_n471), .C1(new_n386), .C2(new_n387), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n394), .A2(new_n471), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT78), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT4), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n408), .A2(KEYINPUT3), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n462), .A2(new_n470), .A3(KEYINPUT74), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT74), .B1(new_n462), .B2(new_n470), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n566), .B(new_n402), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT5), .ZN(new_n571));
  NAND2_X1  g370(.A1(G225gat), .A2(G233gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT76), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n408), .B1(new_n567), .B2(new_n568), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n575), .B2(new_n562), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n574), .B1(new_n576), .B2(new_n571), .ZN(new_n577));
  INV_X1    g376(.A(new_n572), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT74), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n508), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n462), .A2(new_n470), .A3(KEYINPUT74), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n394), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n578), .B1(new_n582), .B2(new_n558), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n388), .A2(KEYINPUT4), .A3(new_n471), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n578), .B1(new_n562), .B2(new_n559), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n569), .A3(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n585), .A2(KEYINPUT77), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT77), .B1(new_n585), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n573), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT0), .B(G57gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G85gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G1gat), .B(G29gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT6), .ZN(new_n597));
  INV_X1    g396(.A(new_n595), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n598), .B(new_n573), .C1(new_n589), .C2(new_n590), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n591), .A2(KEYINPUT6), .A3(new_n595), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n557), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT35), .B1(new_n532), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n554), .A2(new_n556), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(new_n597), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT76), .B1(new_n583), .B2(KEYINPUT5), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n576), .A2(new_n574), .A3(new_n571), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n588), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT77), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n585), .A2(KEYINPUT77), .A3(new_n588), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n598), .B1(new_n612), .B2(new_n573), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n601), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n604), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n434), .A2(new_n530), .A3(new_n531), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT87), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n434), .A2(new_n530), .A3(KEYINPUT87), .A4(new_n531), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n603), .B1(new_n621), .B2(KEYINPUT35), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n434), .A2(new_n531), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT83), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT83), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n434), .A2(new_n625), .A3(new_n531), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n616), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n530), .B(KEYINPUT36), .ZN(new_n628));
  INV_X1    g427(.A(new_n623), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n544), .A2(new_n404), .A3(new_n545), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n538), .B1(new_n535), .B2(new_n542), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n630), .B(KEYINPUT86), .C1(new_n631), .C2(new_n404), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n632), .B(KEYINPUT37), .C1(KEYINPUT86), .C2(new_n630), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n551), .B1(new_n547), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n600), .A2(new_n601), .A3(new_n637), .A4(new_n552), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n543), .A2(KEYINPUT37), .A3(new_n546), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n634), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n629), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n575), .A2(new_n572), .A3(new_n562), .ZN(new_n642));
  OAI211_X1 g441(.A(KEYINPUT39), .B(new_n642), .C1(new_n570), .C2(new_n572), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n572), .B1(new_n565), .B2(new_n569), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n595), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(KEYINPUT40), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n596), .A2(new_n556), .A3(new_n554), .A4(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT40), .B1(new_n643), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT84), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT85), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n554), .A2(new_n556), .A3(new_n647), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT84), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n649), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT85), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n652), .A2(new_n654), .A3(new_n655), .A4(new_n596), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n627), .B(new_n628), .C1(new_n641), .C2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n338), .B1(new_n622), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G113gat), .B(G141gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G169gat), .B(G197gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT12), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n214), .A2(new_n219), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n312), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT91), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT91), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n667), .A2(new_n670), .A3(new_n312), .ZN(new_n671));
  AND4_X1   g470(.A1(new_n304), .A2(new_n303), .A3(new_n296), .A4(new_n286), .ZN(new_n672));
  INV_X1    g471(.A(new_n297), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n286), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT17), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n298), .A2(new_n299), .A3(new_n305), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n669), .A2(new_n671), .B1(new_n678), .B2(new_n220), .ZN(new_n679));
  NAND2_X1  g478(.A1(G229gat), .A2(G233gat), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT18), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n666), .B1(new_n681), .B2(KEYINPUT93), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n220), .B1(new_n306), .B2(new_n307), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n667), .A2(new_n670), .A3(new_n312), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n670), .B1(new_n667), .B2(new_n312), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n683), .B(new_n680), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT18), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n680), .B(KEYINPUT13), .Z(new_n689));
  NOR2_X1   g488(.A1(new_n684), .A2(new_n685), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n672), .A2(new_n675), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT92), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n220), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT92), .B1(new_n667), .B2(new_n312), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n689), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n669), .A2(new_n671), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n697), .A2(KEYINPUT18), .A3(new_n680), .A4(new_n683), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n688), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n688), .A2(new_n696), .A3(new_n698), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT93), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n688), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n703), .A3(new_n666), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n277), .A2(KEYINPUT99), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n244), .A2(new_n313), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n230), .A2(new_n240), .A3(new_n707), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n281), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(G230gat), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n317), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT10), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n708), .A2(new_n716), .A3(new_n710), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n244), .A2(new_n313), .A3(KEYINPUT10), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n714), .ZN(new_n720));
  XNOR2_X1  g519(.A(G120gat), .B(G148gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(new_n481), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(new_n340), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n715), .A2(new_n720), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n711), .A2(new_n714), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n725), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT100), .B(new_n723), .C1(new_n727), .C2(new_n726), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n706), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n659), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n614), .A2(new_n615), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n207), .ZN(G1324gat));
  NOR2_X1   g538(.A1(new_n735), .A2(new_n604), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n740), .A2(new_n741), .A3(G8gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(KEYINPUT102), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT101), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT16), .B(G8gat), .Z(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n742), .B1(new_n740), .B2(new_n746), .ZN(G1325gat));
  INV_X1    g546(.A(new_n530), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n209), .B1(new_n735), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n628), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n659), .A2(G15gat), .A3(new_n734), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT103), .ZN(G1326gat));
  NAND2_X1  g552(.A1(new_n624), .A2(new_n626), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n735), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT43), .B(G22gat), .Z(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1327gat));
  NAND2_X1  g556(.A1(new_n622), .A2(new_n658), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n337), .A2(new_n335), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n264), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n734), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n289), .A3(new_n736), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n758), .A2(new_n767), .A3(new_n759), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n762), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT104), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n767), .B1(new_n758), .B2(new_n759), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n332), .A2(new_n333), .A3(new_n322), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n333), .B1(new_n332), .B2(new_n322), .ZN(new_n775));
  INV_X1    g574(.A(new_n330), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n336), .ZN(new_n778));
  AOI211_X1 g577(.A(KEYINPUT44), .B(new_n778), .C1(new_n622), .C2(new_n658), .ZN(new_n779));
  OAI211_X1 g578(.A(KEYINPUT104), .B(new_n770), .C1(new_n773), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n737), .B1(new_n772), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n765), .B1(new_n781), .B2(new_n289), .ZN(G1328gat));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n290), .A3(new_n557), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT46), .Z(new_n784));
  AOI21_X1  g583(.A(new_n604), .B1(new_n772), .B2(new_n780), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n290), .ZN(G1329gat));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n770), .ZN(new_n787));
  OAI21_X1  g586(.A(G43gat), .B1(new_n787), .B2(new_n628), .ZN(new_n788));
  INV_X1    g587(.A(new_n763), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n789), .A2(G43gat), .A3(new_n748), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n791), .A3(KEYINPUT47), .ZN(new_n792));
  INV_X1    g591(.A(new_n780), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n750), .B1(new_n771), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n794), .B2(G43gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n792), .B1(new_n795), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g595(.A(G50gat), .B1(new_n787), .B2(new_n629), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n789), .A2(G50gat), .A3(new_n754), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n799), .A3(KEYINPUT48), .ZN(new_n800));
  INV_X1    g599(.A(new_n754), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n771), .B2(new_n793), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n798), .B1(new_n802), .B2(G50gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n803), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g603(.A(new_n732), .B1(new_n622), .B2(new_n658), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n338), .A2(new_n705), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n736), .B(KEYINPUT105), .Z(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(new_n234), .ZN(G1332gat));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n604), .ZN(new_n811));
  NOR2_X1   g610(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n812));
  AND2_X1   g611(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n811), .B2(new_n812), .ZN(G1333gat));
  INV_X1    g614(.A(new_n807), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(G71gat), .A3(new_n750), .ZN(new_n817));
  OR3_X1    g616(.A1(new_n807), .A2(KEYINPUT106), .A3(new_n748), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT106), .B1(new_n807), .B2(new_n748), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n817), .B1(new_n820), .B2(G71gat), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g621(.A1(new_n816), .A2(new_n801), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g623(.A1(new_n264), .A2(new_n705), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n758), .A2(new_n759), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n758), .A2(KEYINPUT51), .A3(new_n759), .A4(new_n825), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n732), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(G85gat), .B1(new_n830), .B2(new_n736), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n733), .B(new_n825), .C1(new_n773), .C2(new_n779), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n832), .A2(new_n271), .A3(new_n737), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n831), .A2(new_n833), .ZN(G1336gat));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n557), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n272), .ZN(new_n836));
  OR3_X1    g635(.A1(new_n832), .A2(new_n272), .A3(new_n604), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT107), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT52), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n838), .A2(KEYINPUT52), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n836), .A2(new_n837), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(G92gat), .B1(new_n830), .B2(new_n557), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n832), .A2(new_n272), .A3(new_n604), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n838), .B(KEYINPUT52), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n841), .A2(new_n844), .ZN(G1337gat));
  INV_X1    g644(.A(G99gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n846), .A3(new_n530), .ZN(new_n847));
  OAI21_X1  g646(.A(G99gat), .B1(new_n832), .B2(new_n628), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1338gat));
  NAND2_X1  g648(.A1(new_n828), .A2(new_n829), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n629), .A2(G106gat), .A3(new_n732), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT109), .Z(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT110), .ZN(new_n854));
  XNOR2_X1  g653(.A(KEYINPUT108), .B(G106gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n832), .B2(new_n754), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n857), .A3(new_n852), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT53), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n855), .B1(new_n832), .B2(new_n629), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT53), .B1(new_n850), .B2(new_n851), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(G1339gat));
  NAND3_X1  g663(.A1(new_n806), .A2(KEYINPUT111), .A3(new_n732), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n778), .A2(new_n706), .A3(new_n264), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n733), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n717), .A2(new_n713), .A3(new_n718), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n727), .B2(KEYINPUT112), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n717), .A2(new_n872), .A3(new_n713), .A4(new_n718), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(KEYINPUT54), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n724), .B1(new_n727), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(KEYINPUT55), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT55), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n720), .A2(new_n872), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n870), .ZN(new_n881));
  INV_X1    g680(.A(new_n876), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n705), .A2(new_n725), .A3(new_n877), .A4(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n664), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n690), .A2(new_n695), .A3(new_n689), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n680), .B1(new_n697), .B2(new_n683), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n688), .A2(new_n696), .A3(new_n665), .A4(new_n698), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n732), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n759), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n877), .B(new_n883), .C1(new_n777), .C2(new_n336), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT113), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT113), .B1(new_n888), .B2(new_n889), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n725), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT114), .ZN(new_n900));
  INV_X1    g699(.A(new_n725), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT113), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n890), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT113), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n881), .A2(new_n878), .A3(new_n882), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT55), .B1(new_n874), .B2(new_n876), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n759), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT114), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n900), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n869), .B1(new_n912), .B2(new_n761), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n913), .A2(new_n801), .A3(new_n748), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n737), .A2(new_n557), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G113gat), .B1(new_n916), .B2(new_n706), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n808), .A2(new_n557), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n912), .A2(new_n761), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n868), .A3(new_n865), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n619), .A2(new_n620), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n705), .A2(new_n465), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT115), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n917), .B1(new_n925), .B2(new_n927), .ZN(G1340gat));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n463), .A3(new_n733), .ZN(new_n929));
  OAI21_X1  g728(.A(G120gat), .B1(new_n916), .B2(new_n732), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1341gat));
  AOI21_X1  g730(.A(G127gat), .B1(new_n924), .B2(new_n264), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n458), .A3(new_n761), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(G1342gat));
  NAND3_X1  g733(.A1(new_n924), .A2(new_n456), .A3(new_n759), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT56), .Z(new_n936));
  OAI21_X1  g735(.A(G134gat), .B1(new_n916), .B2(new_n778), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1343gat));
  NAND2_X1  g737(.A1(new_n915), .A2(new_n628), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT57), .B1(new_n920), .B2(new_n623), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT57), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n913), .A2(new_n942), .A3(new_n754), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n705), .B(new_n940), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G141gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n628), .A2(new_n623), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n921), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n382), .A3(new_n705), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT116), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT116), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n945), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT58), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n950), .A2(KEYINPUT58), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1344gat));
  NAND3_X1  g756(.A1(new_n947), .A2(new_n380), .A3(new_n733), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n941), .A2(new_n943), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(new_n939), .ZN(new_n960));
  AOI211_X1 g759(.A(KEYINPUT59), .B(new_n380), .C1(new_n960), .C2(new_n733), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT59), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT118), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n893), .B2(new_n899), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n901), .B1(new_n700), .B2(new_n704), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n891), .B1(new_n908), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n909), .B(KEYINPUT118), .C1(new_n966), .C2(new_n759), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n761), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT117), .B1(new_n806), .B2(new_n732), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT117), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n867), .A2(new_n970), .A3(new_n733), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n801), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT119), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n974), .A2(new_n975), .A3(new_n942), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n754), .B1(new_n968), .B2(new_n972), .ZN(new_n977));
  OAI21_X1  g776(.A(KEYINPUT119), .B1(new_n977), .B2(KEYINPUT57), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n920), .A2(KEYINPUT57), .A3(new_n623), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n733), .A3(new_n940), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n962), .B1(new_n981), .B2(G148gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n958), .B1(new_n961), .B2(new_n982), .ZN(G1345gat));
  AOI21_X1  g782(.A(G155gat), .B1(new_n947), .B2(new_n264), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n761), .A2(new_n368), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n984), .B1(new_n960), .B2(new_n985), .ZN(G1346gat));
  AOI21_X1  g785(.A(G162gat), .B1(new_n947), .B2(new_n759), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n778), .A2(new_n369), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n987), .B1(new_n960), .B2(new_n988), .ZN(G1347gat));
  AND2_X1   g788(.A1(new_n808), .A2(new_n557), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n914), .A2(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(G169gat), .B1(new_n992), .B2(new_n706), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n920), .A2(KEYINPUT120), .A3(new_n737), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT120), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n995), .B1(new_n913), .B2(new_n736), .ZN(new_n996));
  AOI211_X1 g795(.A(new_n604), .B(new_n923), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n997), .A2(new_n480), .A3(new_n705), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n993), .A2(new_n998), .ZN(G1348gat));
  NOR3_X1   g798(.A1(new_n992), .A2(new_n481), .A3(new_n732), .ZN(new_n1000));
  AOI21_X1  g799(.A(G176gat), .B1(new_n997), .B2(new_n733), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1349gat));
  AOI21_X1  g801(.A(new_n923), .B1(new_n994), .B2(new_n996), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n1003), .A2(new_n447), .A3(new_n557), .A4(new_n264), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n914), .A2(new_n264), .A3(new_n990), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(G183gat), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(KEYINPUT121), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT121), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1004), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n1008), .A2(KEYINPUT60), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g810(.A(KEYINPUT60), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1011), .A2(new_n1012), .ZN(G1350gat));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n442), .A3(new_n759), .ZN(new_n1014));
  XNOR2_X1  g813(.A(new_n1014), .B(KEYINPUT122), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n442), .B1(new_n991), .B2(new_n759), .ZN(new_n1016));
  XOR2_X1   g815(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n1017));
  NAND2_X1  g816(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OR2_X1    g817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1015), .A2(new_n1018), .A3(new_n1019), .ZN(G1351gat));
  NAND2_X1  g819(.A1(new_n994), .A2(new_n996), .ZN(new_n1021));
  INV_X1    g820(.A(new_n946), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1021), .A2(new_n557), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1023), .A2(KEYINPUT124), .ZN(new_n1024));
  INV_X1    g823(.A(KEYINPUT124), .ZN(new_n1025));
  NAND4_X1  g824(.A1(new_n1021), .A2(new_n1025), .A3(new_n557), .A4(new_n1022), .ZN(new_n1026));
  NAND4_X1  g825(.A1(new_n1024), .A2(new_n339), .A3(new_n705), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g826(.A(KEYINPUT125), .ZN(new_n1028));
  AND2_X1   g827(.A1(new_n990), .A2(new_n628), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n980), .A2(new_n705), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1030), .A2(G197gat), .ZN(new_n1031));
  AND3_X1   g830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1028), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1033));
  NOR2_X1   g832(.A1(new_n1032), .A2(new_n1033), .ZN(G1352gat));
  NOR3_X1   g833(.A1(new_n1023), .A2(G204gat), .A3(new_n732), .ZN(new_n1035));
  INV_X1    g834(.A(KEYINPUT62), .ZN(new_n1036));
  OR2_X1    g835(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  AND3_X1   g837(.A1(new_n980), .A2(new_n733), .A3(new_n1029), .ZN(new_n1039));
  OAI211_X1 g838(.A(new_n1037), .B(new_n1038), .C1(new_n340), .C2(new_n1039), .ZN(G1353gat));
  NAND3_X1  g839(.A1(new_n980), .A2(new_n264), .A3(new_n1029), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1041), .A2(KEYINPUT126), .ZN(new_n1042));
  INV_X1    g841(.A(KEYINPUT126), .ZN(new_n1043));
  NAND4_X1  g842(.A1(new_n980), .A2(new_n1043), .A3(new_n264), .A4(new_n1029), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n1042), .A2(G211gat), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g844(.A(KEYINPUT63), .ZN(new_n1046));
  NAND2_X1  g845(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g846(.A1(new_n1042), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n1044), .ZN(new_n1048));
  NAND2_X1  g847(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g848(.A1(new_n1024), .A2(new_n246), .A3(new_n264), .A4(new_n1026), .ZN(new_n1050));
  NAND2_X1  g849(.A1(new_n1049), .A2(new_n1050), .ZN(G1354gat));
  AND4_X1   g850(.A1(G218gat), .A2(new_n980), .A3(new_n759), .A4(new_n1029), .ZN(new_n1052));
  NAND3_X1  g851(.A1(new_n1024), .A2(new_n759), .A3(new_n1026), .ZN(new_n1053));
  NAND2_X1  g852(.A1(new_n1053), .A2(new_n350), .ZN(new_n1054));
  INV_X1    g853(.A(KEYINPUT127), .ZN(new_n1055));
  NAND2_X1  g854(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g855(.A1(new_n1053), .A2(KEYINPUT127), .A3(new_n350), .ZN(new_n1057));
  AOI21_X1  g856(.A(new_n1052), .B1(new_n1056), .B2(new_n1057), .ZN(G1355gat));
endmodule


