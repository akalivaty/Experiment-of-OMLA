//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT64), .Z(new_n213));
  AOI211_X1 g0013(.A(new_n211), .B(new_n213), .C1(G77), .C2(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G116), .ZN(new_n217));
  INV_X1    g0017(.A(G270), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n203), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n206), .B(new_n224), .C1(new_n227), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n216), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT65), .B(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G270), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G222), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n250), .B(new_n252), .C1(new_n253), .C2(new_n251), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(G1), .B(G13), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n254), .B(new_n258), .C1(G77), .C2(new_n250), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n261), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n259), .B(new_n264), .C1(new_n208), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G169), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(G20), .B1(new_n229), .B2(G50), .ZN(new_n269));
  INV_X1    g0069(.A(G150), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n226), .A2(G33), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n269), .B1(new_n270), .B2(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n225), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n207), .ZN(new_n281));
  INV_X1    g0081(.A(new_n277), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n260), .A2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n278), .B(new_n281), .C1(new_n207), .C2(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n268), .B(new_n285), .C1(G179), .C2(new_n266), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n285), .B(KEYINPUT9), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n266), .A2(G200), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n266), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n288), .A2(KEYINPUT68), .A3(new_n289), .A4(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n292), .A2(KEYINPUT10), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(KEYINPUT10), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n287), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT67), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G238), .A2(G1698), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n250), .B(new_n297), .C1(new_n216), .C2(G1698), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n258), .C1(G107), .C2(new_n250), .ZN(new_n299));
  INV_X1    g0099(.A(new_n265), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G244), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n264), .A3(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n302), .A2(new_n290), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(G200), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n282), .A2(G77), .A3(new_n283), .ZN(new_n305));
  INV_X1    g0105(.A(new_n273), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n306), .A2(new_n271), .B1(G20), .B2(G77), .ZN(new_n307));
  XOR2_X1   g0107(.A(KEYINPUT15), .B(G87), .Z(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n307), .B1(new_n274), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G77), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n310), .A2(new_n277), .B1(new_n311), .B2(new_n280), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n305), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n302), .A2(G179), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n302), .A2(new_n267), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT75), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT3), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT71), .B1(new_n320), .B2(G33), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(new_n255), .A3(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n253), .A2(new_n251), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n208), .A2(G1698), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G87), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n258), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n264), .B1(new_n265), .B2(new_n216), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n290), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n257), .B1(new_n328), .B2(new_n329), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n332), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n334), .A2(KEYINPUT74), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT74), .B1(new_n334), .B2(new_n337), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n324), .A2(new_n325), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT7), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(new_n226), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n321), .B2(new_n323), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT7), .B1(new_n346), .B2(G20), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(G68), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n215), .A2(new_n209), .ZN(new_n349));
  OAI21_X1  g0149(.A(G20), .B1(new_n349), .B2(new_n228), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n271), .A2(G159), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n348), .A2(KEYINPUT16), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n343), .A2(KEYINPUT72), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT7), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n250), .B2(G20), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n325), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(new_n226), .A3(new_n356), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n209), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n355), .B1(new_n364), .B2(new_n352), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n354), .A2(new_n277), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n284), .A2(new_n306), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n280), .B2(new_n306), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n340), .A2(new_n341), .A3(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n366), .A2(new_n368), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT74), .ZN(new_n372));
  AOI21_X1  g0172(.A(G200), .B1(new_n331), .B2(new_n333), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n336), .A2(G190), .A3(new_n332), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n334), .A2(KEYINPUT74), .A3(new_n337), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT17), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n319), .B1(new_n370), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n341), .B1(new_n340), .B2(new_n369), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n371), .A2(new_n377), .A3(KEYINPUT17), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(KEYINPUT75), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n336), .A2(new_n332), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G179), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n267), .B2(new_n383), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n369), .A2(KEYINPUT18), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n369), .A2(new_n385), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n387), .A3(new_n390), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n379), .A2(new_n382), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  OAI221_X1 g0195(.A(new_n295), .B1(new_n296), .B2(new_n318), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT69), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n265), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT69), .B1(new_n257), .B2(new_n261), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(G238), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G97), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n255), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(G226), .A2(G1698), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n216), .B2(G1698), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n405), .B1(new_n407), .B2(new_n250), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n264), .B1(new_n408), .B2(new_n257), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n397), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n399), .A2(new_n210), .A3(new_n401), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n412), .A2(new_n409), .A3(KEYINPUT13), .ZN(new_n413));
  OAI21_X1  g0213(.A(G169), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n403), .A2(new_n410), .A3(new_n397), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT13), .B1(new_n412), .B2(new_n409), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(G179), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(G169), .C1(new_n411), .C2(new_n413), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n272), .A2(new_n207), .B1(new_n226), .B2(G68), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n274), .A2(new_n311), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n277), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g0224(.A(new_n424), .B(KEYINPUT11), .Z(new_n425));
  INV_X1    g0225(.A(KEYINPUT12), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n280), .B2(new_n209), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n279), .A2(KEYINPUT12), .A3(G68), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n427), .A2(new_n428), .B1(new_n284), .B2(new_n209), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G200), .B1(new_n411), .B2(new_n413), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n416), .A2(new_n417), .A3(G190), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT70), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT70), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n432), .A2(new_n430), .A3(new_n436), .A4(new_n433), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n421), .A2(new_n431), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n318), .A2(new_n296), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n392), .A2(new_n393), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n380), .A2(KEYINPUT75), .A3(new_n381), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT75), .B1(new_n380), .B2(new_n381), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n438), .B(new_n439), .C1(new_n443), .C2(KEYINPUT76), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n396), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G257), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n251), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n221), .A2(G1698), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n324), .A2(new_n325), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n362), .A2(G303), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n258), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT5), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(G41), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n256), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n455), .A2(new_n456), .A3(new_n458), .A4(G274), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n455), .A2(new_n458), .A3(new_n456), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n461), .A2(new_n257), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n462), .B2(G270), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n452), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n280), .A2(new_n217), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n260), .A2(G33), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n282), .A2(G116), .A3(new_n279), .A4(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n276), .A2(new_n225), .B1(G20), .B2(new_n217), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n469), .B(new_n226), .C1(G33), .C2(new_n404), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n468), .A2(KEYINPUT20), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT20), .B1(new_n468), .B2(new_n470), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n465), .B(new_n467), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n464), .A2(KEYINPUT21), .A3(G169), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT21), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(G169), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n257), .B1(new_n449), .B2(new_n450), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n461), .A2(new_n257), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n459), .B1(new_n478), .B2(new_n218), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n475), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G179), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n477), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n473), .ZN(new_n485));
  INV_X1    g0285(.A(new_n473), .ZN(new_n486));
  OAI21_X1  g0286(.A(G200), .B1(new_n477), .B2(new_n479), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n487), .C1(new_n464), .C2(new_n290), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n482), .A2(KEYINPUT82), .A3(new_n485), .A4(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n488), .A2(new_n474), .A3(new_n481), .A4(new_n485), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n459), .B1(new_n478), .B2(new_n446), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT4), .B1(new_n346), .B2(G244), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n361), .A2(new_n325), .A3(G250), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n251), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(new_n361), .A3(new_n325), .A4(G244), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n469), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n496), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n495), .B1(new_n503), .B2(new_n257), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G169), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n324), .A2(G244), .A3(new_n325), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n499), .ZN(new_n507));
  INV_X1    g0307(.A(new_n498), .ZN(new_n508));
  INV_X1    g0308(.A(new_n502), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n494), .B1(new_n510), .B2(new_n258), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G179), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n279), .A2(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n360), .A2(new_n363), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G107), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n272), .A2(new_n311), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT77), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT77), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n521));
  AOI211_X1 g0321(.A(new_n404), .B(G107), .C1(new_n519), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n220), .A2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n404), .A2(G107), .ZN(new_n524));
  AND4_X1   g0324(.A1(new_n523), .A2(new_n519), .A3(new_n521), .A4(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n515), .B(new_n517), .C1(new_n526), .C2(new_n226), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n513), .B1(new_n527), .B2(new_n277), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n282), .A2(new_n279), .A3(new_n466), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G97), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n505), .A2(new_n512), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n511), .A2(new_n335), .ZN(new_n533));
  INV_X1    g0333(.A(new_n513), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n220), .B1(new_n360), .B2(new_n363), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n518), .A2(KEYINPUT77), .ZN(new_n537));
  OAI211_X1 g0337(.A(G97), .B(new_n220), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n523), .A2(new_n519), .A3(new_n521), .A4(new_n524), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n226), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n535), .A2(new_n540), .A3(new_n516), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n531), .B(new_n534), .C1(new_n541), .C2(new_n282), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT78), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n517), .B1(new_n526), .B2(new_n226), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n277), .B1(new_n545), .B2(new_n535), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(KEYINPUT78), .A3(new_n531), .A4(new_n534), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n533), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT80), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n504), .A2(new_n549), .A3(new_n290), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT80), .B1(new_n511), .B2(G190), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n532), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G87), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n529), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n308), .A2(new_n279), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n346), .A2(new_n226), .A3(G68), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n274), .B2(new_n404), .ZN(new_n559));
  AOI21_X1  g0359(.A(G20), .B1(new_n405), .B2(KEYINPUT19), .ZN(new_n560));
  NOR3_X1   g0360(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n557), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n555), .B(new_n556), .C1(new_n562), .C2(new_n277), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G244), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n210), .B2(G1698), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n322), .B1(KEYINPUT3), .B2(new_n255), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n320), .A2(KEYINPUT71), .A3(G33), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n325), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n255), .A2(new_n217), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT81), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT81), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n568), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n258), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G250), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n458), .A2(new_n576), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n577), .B(new_n258), .C1(G274), .C2(new_n458), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(G200), .A3(new_n579), .ZN(new_n580));
  AOI211_X1 g0380(.A(KEYINPUT81), .B(new_n569), .C1(new_n346), .C2(new_n565), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n573), .B1(new_n568), .B2(new_n570), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n578), .B1(new_n583), .B2(new_n258), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n563), .B(new_n580), .C1(new_n584), .C2(new_n290), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n562), .A2(new_n277), .ZN(new_n586));
  INV_X1    g0386(.A(new_n556), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n530), .A2(new_n308), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n575), .A2(new_n267), .A3(new_n579), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n584), .C2(G179), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT22), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n593), .A2(new_n554), .A3(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n324), .A2(new_n325), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n220), .A2(G20), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT23), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n554), .A2(G20), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n361), .A3(new_n325), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n593), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n569), .A2(new_n226), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n595), .A2(new_n598), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT24), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n346), .A2(new_n594), .B1(new_n593), .B2(new_n600), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT24), .A3(new_n598), .A4(new_n602), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n607), .A3(new_n277), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n530), .A2(G107), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n279), .A2(G107), .ZN(new_n610));
  XNOR2_X1  g0410(.A(KEYINPUT83), .B(KEYINPUT25), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n461), .A2(G264), .A3(new_n257), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n576), .A2(new_n251), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n446), .A2(G1698), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n324), .A2(new_n325), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G33), .A2(G294), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n614), .B1(new_n619), .B2(new_n258), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n459), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n267), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n483), .A3(new_n459), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n613), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(new_n258), .ZN(new_n625));
  INV_X1    g0425(.A(new_n614), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(G190), .A3(new_n459), .A4(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n608), .A2(new_n627), .A3(new_n609), .A4(new_n612), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n335), .B1(new_n620), .B2(new_n459), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n592), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n445), .A2(new_n493), .A3(new_n553), .A4(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n532), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT26), .B1(new_n633), .B2(new_n592), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n548), .A2(new_n552), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n628), .A2(new_n629), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n613), .A2(new_n622), .A3(new_n623), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n482), .A2(new_n637), .A3(new_n485), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n635), .A2(new_n633), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n591), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n563), .A2(new_n580), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n575), .A2(new_n579), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n641), .A2(KEYINPUT84), .B1(G190), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT84), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n563), .A2(new_n580), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n640), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n634), .B1(new_n639), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n645), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n505), .A2(new_n512), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n650), .A2(new_n544), .A3(new_n547), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n651), .A3(new_n591), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n591), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n445), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n435), .A2(new_n437), .ZN(new_n656));
  INV_X1    g0456(.A(new_n317), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n421), .A2(new_n431), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n379), .A2(new_n382), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n391), .A2(new_n386), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n293), .A2(new_n294), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n287), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n655), .A2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n260), .A2(new_n226), .A3(G13), .ZN(new_n668));
  OR3_X1    g0468(.A1(new_n668), .A2(KEYINPUT85), .A3(KEYINPUT27), .ZN(new_n669));
  INV_X1    g0469(.A(G213), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n668), .B2(KEYINPUT27), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT85), .B1(new_n668), .B2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT86), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n493), .B1(new_n486), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n482), .A2(new_n485), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n473), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT87), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n613), .A2(new_n679), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n637), .B1(new_n687), .B2(new_n630), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n624), .A2(new_n680), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n679), .B1(new_n482), .B2(new_n485), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n689), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT88), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(KEYINPUT88), .A3(new_n689), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n691), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n204), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G1), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n561), .A2(new_n217), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n703), .A2(new_n704), .B1(new_n230), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n654), .A2(new_n707), .A3(new_n680), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n635), .A2(new_n633), .A3(new_n638), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT92), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(new_n636), .A4(new_n646), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT26), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n532), .A2(new_n713), .A3(new_n585), .A4(new_n591), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n591), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(KEYINPUT26), .B2(new_n652), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT92), .B1(new_n639), .B2(new_n647), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n707), .B1(new_n718), .B2(new_n680), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n631), .A2(new_n493), .A3(new_n553), .A4(new_n680), .ZN(new_n720));
  XOR2_X1   g0520(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n721));
  AOI21_X1  g0521(.A(G179), .B1(new_n620), .B2(new_n459), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n584), .A2(new_n722), .A3(new_n464), .A4(new_n504), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n642), .A2(new_n484), .A3(new_n511), .A4(new_n620), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g0526(.A(KEYINPUT90), .B(KEYINPUT30), .Z(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n511), .A2(new_n620), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n452), .A2(new_n463), .A3(G179), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n579), .B2(new_n575), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n728), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n679), .B(new_n721), .C1(new_n726), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT91), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n726), .B2(new_n732), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n729), .A2(new_n731), .A3(KEYINPUT30), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n724), .A2(new_n727), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT91), .A4(new_n723), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n679), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n720), .B(new_n733), .C1(new_n740), .C2(KEYINPUT31), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n709), .A2(new_n719), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n706), .B1(new_n743), .B2(G1), .ZN(G364));
  INV_X1    g0544(.A(G13), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n703), .B1(G45), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n686), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G330), .B2(new_n685), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n290), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n483), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n226), .A2(G179), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G190), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n752), .A2(G294), .B1(new_n756), .B2(G329), .ZN(new_n757));
  INV_X1    g0557(.A(G322), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n226), .A2(new_n483), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT95), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(KEYINPUT95), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n760), .A2(new_n761), .A3(new_n750), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n757), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G190), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G317), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(KEYINPUT33), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(KEYINPUT33), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n764), .A2(new_n290), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n250), .B1(new_n770), .B2(G326), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n760), .A2(new_n761), .A3(new_n754), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n763), .B(new_n772), .C1(G311), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n753), .A2(new_n290), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(G303), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n753), .A2(G190), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT96), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n775), .B1(new_n776), .B2(new_n777), .C1(new_n778), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n777), .A2(new_n220), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n765), .A2(G68), .B1(new_n752), .B2(G97), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT97), .Z(new_n787));
  AOI211_X1 g0587(.A(new_n785), .B(new_n787), .C1(G77), .C2(new_n774), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n755), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  INV_X1    g0591(.A(new_n783), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n792), .A2(G87), .B1(G50), .B2(new_n770), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n788), .A2(new_n250), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n762), .A2(new_n215), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n784), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n225), .B1(G20), .B2(new_n267), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n681), .A2(new_n683), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n700), .A2(new_n362), .ZN(new_n803));
  XNOR2_X1  g0603(.A(G355), .B(KEYINPUT93), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n346), .A2(new_n700), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n457), .B2(new_n231), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT94), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n457), .B2(new_n248), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(KEYINPUT94), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n805), .B1(G116), .B2(new_n204), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n801), .A2(new_n797), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n798), .A2(new_n802), .A3(new_n814), .A4(new_n747), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n749), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n654), .A2(new_n680), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n679), .A2(new_n314), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n313), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n317), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n657), .A2(new_n680), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT99), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT99), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n680), .B(new_n827), .C1(new_n648), .C2(new_n653), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(new_n742), .ZN(new_n832));
  INV_X1    g0632(.A(new_n747), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n762), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(G143), .B1(G150), .B2(new_n765), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  INV_X1    g0637(.A(new_n770), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(new_n837), .B2(new_n838), .C1(new_n789), .C2(new_n773), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT34), .ZN(new_n840));
  INV_X1    g0640(.A(new_n752), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n841), .A2(new_n215), .B1(new_n842), .B2(new_n755), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n342), .B(new_n843), .C1(new_n792), .C2(G50), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n840), .B(new_n844), .C1(new_n209), .C2(new_n777), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n774), .A2(G116), .B1(G303), .B2(new_n770), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n776), .B2(new_n766), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT98), .Z(new_n848));
  AOI211_X1 g0648(.A(new_n250), .B(new_n848), .C1(G107), .C2(new_n792), .ZN(new_n849));
  INV_X1    g0649(.A(G311), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n554), .B2(new_n777), .C1(new_n850), .C2(new_n755), .ZN(new_n851));
  INV_X1    g0651(.A(G294), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n762), .A2(new_n852), .B1(new_n841), .B2(new_n404), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n845), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n797), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n797), .A2(new_n799), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n311), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n828), .A2(new_n799), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n855), .A2(new_n747), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n834), .A2(new_n859), .ZN(G384));
  INV_X1    g0660(.A(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n354), .A2(new_n277), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT16), .B1(new_n348), .B2(new_n353), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n368), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n677), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n443), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n371), .A2(new_n377), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n369), .A2(new_n865), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n389), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n864), .B1(new_n385), .B2(new_n865), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n873), .A2(new_n869), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n874), .B2(new_n870), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT38), .B1(new_n868), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n870), .B1(new_n873), .B2(new_n869), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n869), .A2(new_n389), .A3(new_n871), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n878), .B1(new_n879), .B2(new_n870), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n877), .B(new_n880), .C1(new_n443), .C2(new_n867), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n861), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n866), .B1(new_n661), .B2(new_n440), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n877), .B1(new_n883), .B2(new_n880), .ZN(new_n884));
  OAI211_X1 g0684(.A(KEYINPUT38), .B(new_n875), .C1(new_n394), .C2(new_n866), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(KEYINPUT101), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n659), .A2(new_n656), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n680), .A2(new_n430), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n887), .A2(KEYINPUT100), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT100), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n438), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n888), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n438), .B2(new_n890), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n822), .B2(new_n830), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n882), .A2(new_n886), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n869), .A2(new_n389), .A3(new_n871), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(new_n870), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n370), .A2(new_n378), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n871), .B1(new_n899), .B2(new_n663), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n877), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n885), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n421), .A2(new_n431), .A3(new_n680), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT102), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n391), .A2(new_n386), .A3(new_n677), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n896), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n445), .B1(new_n709), .B2(new_n719), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n666), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n910), .B(new_n912), .Z(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n893), .A2(new_n891), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n438), .A2(new_n890), .A3(new_n892), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n828), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n739), .A2(KEYINPUT103), .ZN(new_n918));
  INV_X1    g0718(.A(new_n721), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT103), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n735), .A2(new_n920), .A3(new_n679), .A4(new_n738), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT104), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n679), .A4(new_n738), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n720), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n923), .B1(new_n922), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n917), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n902), .A2(KEYINPUT40), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n922), .A2(new_n925), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT104), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n922), .A2(new_n925), .A3(new_n923), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n882), .A2(new_n934), .A3(new_n917), .A4(new_n886), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n445), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n936), .ZN(new_n939));
  INV_X1    g0739(.A(new_n930), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(G330), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(new_n445), .A3(G330), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n938), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n914), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n914), .A2(new_n945), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(new_n260), .C2(new_n746), .ZN(new_n948));
  INV_X1    g0748(.A(new_n526), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n217), .B1(new_n949), .B2(KEYINPUT35), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n227), .C1(KEYINPUT35), .C2(new_n949), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  OAI21_X1  g0752(.A(G77), .B1(new_n215), .B2(new_n209), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n230), .A2(new_n953), .B1(G50), .B2(new_n209), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n745), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n948), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT105), .Z(G367));
  NOR2_X1   g0757(.A1(new_n680), .A2(new_n563), .ZN(new_n958));
  MUX2_X1   g0758(.A(new_n647), .B(new_n591), .S(new_n958), .Z(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n801), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n770), .A2(G143), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n961), .B1(new_n311), .B2(new_n777), .C1(new_n766), .C2(new_n789), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n250), .B1(new_n773), .B2(new_n207), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n752), .A2(G68), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n837), .B2(new_n755), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n215), .B2(new_n783), .C1(new_n270), .C2(new_n762), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n792), .A2(G116), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT46), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n969), .B(new_n342), .C1(new_n778), .C2(new_n762), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n773), .A2(new_n776), .B1(new_n841), .B2(new_n220), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G311), .B2(new_n770), .ZN(new_n972));
  XOR2_X1   g0772(.A(KEYINPUT109), .B(G317), .Z(new_n973));
  NAND2_X1  g0773(.A1(new_n756), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n777), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(G97), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n765), .A2(G294), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n972), .A2(new_n974), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n967), .B1(new_n970), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT47), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n797), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n813), .B1(new_n204), .B2(new_n309), .C1(new_n240), .C2(new_n807), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n747), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT108), .Z(new_n984));
  NAND3_X1  g0784(.A1(new_n960), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n701), .B(KEYINPUT41), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n544), .A2(new_n547), .A3(new_n679), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n553), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n651), .A2(new_n679), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n698), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT44), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n698), .B2(new_n991), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n698), .A2(new_n994), .A3(new_n991), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT45), .ZN(new_n999));
  INV_X1    g0799(.A(new_n997), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n995), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n993), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n691), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n993), .A2(new_n691), .A3(new_n998), .A4(new_n1001), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n690), .B(new_n692), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n686), .B(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n743), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n987), .B1(new_n1008), .B2(new_n743), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n260), .B1(new_n746), .B2(G45), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT106), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1003), .A2(new_n1013), .A3(new_n991), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n710), .A2(new_n690), .A3(new_n692), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT42), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n991), .A2(new_n624), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n679), .B1(new_n1017), .B2(new_n633), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n959), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1014), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n991), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n691), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT106), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1026), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n985), .B1(new_n1012), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(KEYINPUT110), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT110), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n1035), .A2(new_n1026), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1034), .B1(new_n1036), .B2(new_n985), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1033), .A2(new_n1037), .ZN(G387));
  OR2_X1    g0838(.A1(new_n1007), .A2(new_n743), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1007), .A2(new_n743), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n701), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n976), .B1(new_n270), .B2(new_n755), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n342), .B(new_n1043), .C1(G68), .C2(new_n774), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n835), .A2(G50), .B1(new_n308), .B2(new_n752), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n770), .A2(G159), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n792), .A2(G77), .B1(new_n306), .B2(new_n765), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n774), .A2(G303), .B1(G322), .B2(new_n770), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n850), .B2(new_n766), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n835), .B2(new_n973), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT48), .Z(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n776), .B2(new_n841), .C1(new_n852), .C2(new_n783), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT49), .Z(new_n1054));
  AOI21_X1  g0854(.A(new_n346), .B1(G326), .B2(new_n756), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n217), .B2(new_n777), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1048), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n797), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n807), .B1(new_n236), .B2(G45), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n704), .B2(new_n803), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n273), .A2(G50), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n209), .A2(new_n311), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1063), .A2(G45), .A3(new_n1064), .A4(new_n704), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1060), .A2(new_n1065), .B1(G107), .B2(new_n204), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n833), .B1(new_n1066), .B2(new_n813), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n801), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1058), .B(new_n1067), .C1(new_n690), .C2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1041), .A2(new_n1042), .A3(new_n1069), .ZN(G393));
  OAI22_X1  g0870(.A1(new_n783), .A2(new_n209), .B1(new_n554), .B2(new_n777), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n774), .A2(new_n306), .B1(G50), .B2(new_n765), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1071), .B1(new_n1073), .B2(KEYINPUT113), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n789), .A2(new_n762), .B1(new_n838), .B2(new_n270), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n756), .A2(G143), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n346), .B1(new_n841), .B2(new_n311), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT113), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n1072), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1074), .A2(new_n1077), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n765), .A2(G303), .B1(G322), .B2(new_n756), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n217), .B2(new_n841), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n835), .A2(G311), .B1(G317), .B2(new_n770), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(G294), .C2(new_n774), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1087), .B(new_n362), .C1(new_n776), .C2(new_n783), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1082), .B1(new_n1088), .B2(new_n785), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n797), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n244), .A2(new_n806), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1091), .B(new_n813), .C1(new_n404), .C2(new_n204), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n747), .A3(new_n1092), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1093), .A2(KEYINPUT114), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(KEYINPUT114), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n991), .C2(new_n1068), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n702), .B1(new_n1098), .B2(new_n1040), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1097), .B1(new_n1099), .B2(new_n1008), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n1010), .B2(new_n1098), .ZN(G390));
  NAND3_X1  g0901(.A1(new_n718), .A2(new_n680), .A3(new_n827), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n822), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n888), .B1(new_n887), .B2(KEYINPUT100), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n887), .A2(KEYINPUT100), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n916), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n907), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n902), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n904), .A2(new_n905), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n830), .A2(new_n822), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1106), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1108), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT115), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n742), .A2(new_n1115), .A3(new_n827), .A4(new_n1106), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1106), .A2(G330), .A3(new_n741), .A4(new_n827), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(KEYINPUT115), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1109), .A2(new_n1114), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT116), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n917), .C1(new_n926), .C2(new_n927), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT116), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1109), .A2(new_n1114), .A3(new_n1126), .A4(new_n1119), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1121), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n943), .A2(new_n911), .A3(new_n666), .ZN(new_n1129));
  OAI211_X1 g0929(.A(G330), .B(new_n827), .C1(new_n926), .C2(new_n927), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n894), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1103), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(new_n1119), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1106), .B1(new_n742), .B2(new_n827), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1111), .B1(new_n1124), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1129), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n702), .B1(new_n1128), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1136), .A2(new_n1121), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1110), .A2(new_n799), .ZN(new_n1140));
  INV_X1    g0940(.A(G125), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n250), .B1(new_n755), .B2(new_n1141), .C1(new_n207), .C2(new_n777), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT118), .Z(new_n1143));
  AOI22_X1  g0943(.A1(new_n835), .A2(G132), .B1(G159), .B2(new_n752), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n1144), .C1(new_n1145), .C2(new_n838), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT54), .B(G143), .Z(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n773), .A2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n783), .A2(KEYINPUT53), .A3(new_n270), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT53), .B1(new_n783), .B2(new_n270), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n837), .B2(new_n766), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1146), .A2(new_n1149), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n792), .A2(G87), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n756), .A2(G294), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G68), .A2(new_n975), .B1(new_n752), .B2(G77), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n770), .A2(G283), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n766), .A2(new_n220), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n773), .A2(new_n404), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n362), .B1(new_n762), .B2(new_n217), .ZN(new_n1161));
  NOR4_X1   g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n797), .B1(new_n1153), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1140), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n856), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n747), .B1(new_n306), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT117), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1138), .A2(new_n1139), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1128), .A2(new_n1010), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(G378));
  XNOR2_X1  g0970(.A(new_n295), .B(KEYINPUT122), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n865), .A2(new_n285), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AND4_X1   g0980(.A1(G330), .A2(new_n910), .A3(new_n939), .A4(new_n940), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n910), .B1(new_n937), .B2(G330), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n910), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n941), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n937), .A2(G330), .A3(new_n910), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n1179), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1129), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1139), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n701), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT123), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1185), .A2(new_n1179), .A3(new_n1186), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1179), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1139), .A2(new_n1189), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1183), .A2(KEYINPUT123), .A3(new_n1187), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1191), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1195), .A2(new_n1011), .A3(new_n1197), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1179), .A2(new_n800), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1145), .A2(new_n762), .B1(new_n773), .B2(new_n837), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n792), .A2(new_n1147), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1204), .B2(KEYINPUT120), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(KEYINPUT120), .B2(new_n1204), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G150), .B2(new_n752), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n1141), .B2(new_n838), .C1(new_n842), .C2(new_n766), .ZN(new_n1208));
  XOR2_X1   g1008(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1209));
  XNOR2_X1  g1009(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n255), .B1(new_n777), .B2(new_n789), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G124), .B2(new_n756), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n256), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G41), .B1(new_n346), .B2(G33), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(G50), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n774), .A2(new_n308), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n346), .B1(new_n770), .B2(G116), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n765), .A2(G97), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n964), .A4(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n783), .A2(new_n311), .B1(new_n220), .B2(new_n762), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n777), .A2(new_n215), .B1(new_n755), .B2(new_n776), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(new_n1219), .A2(new_n1220), .A3(G41), .A4(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1222), .B(new_n1223), .Z(new_n1224));
  OAI21_X1  g1024(.A(new_n797), .B1(new_n1215), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1165), .A2(G50), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(new_n1202), .A2(new_n833), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1201), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1200), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(G375));
  AND2_X1   g1032(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1129), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1137), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(new_n987), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT124), .Z(new_n1237));
  NOR2_X1   g1037(.A1(new_n1233), .A2(new_n1010), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n856), .A2(new_n209), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n894), .A2(new_n799), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n777), .A2(new_n215), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n841), .A2(new_n207), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(G150), .C2(new_n774), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n837), .B2(new_n762), .C1(new_n789), .C2(new_n783), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n838), .A2(new_n842), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n766), .A2(new_n1148), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n346), .B1(new_n1145), .B2(new_n755), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n777), .A2(new_n311), .B1(new_n755), .B2(new_n778), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n835), .B2(G283), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n220), .B2(new_n773), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n766), .A2(new_n217), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n783), .A2(new_n404), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n362), .B1(new_n841), .B2(new_n309), .C1(new_n838), .C2(new_n852), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n797), .B1(new_n1248), .B2(new_n1255), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1240), .A2(new_n747), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1238), .B1(new_n1239), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1237), .A2(new_n1258), .ZN(G381));
  INV_X1    g1059(.A(G378), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1231), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(G387), .A2(G384), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(G381), .A2(G390), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(G407));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(G343), .C2(new_n1261), .ZN(G409));
  OAI21_X1  g1067(.A(G378), .B1(new_n1200), .B2(new_n1230), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n678), .A2(G213), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1195), .A2(new_n986), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1183), .A2(new_n1011), .A3(new_n1187), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1260), .A2(new_n1270), .A3(new_n1229), .A4(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1268), .A2(new_n1269), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1235), .A2(KEYINPUT60), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1234), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n701), .A3(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(G384), .A3(new_n1258), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1277), .B2(new_n1258), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n678), .A2(G213), .A3(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1279), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1277), .A2(new_n1258), .ZN(new_n1284));
  INV_X1    g1084(.A(G384), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1281), .B1(new_n1286), .B2(new_n1278), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1273), .A2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1268), .A2(new_n1290), .A3(new_n1269), .A4(new_n1272), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT63), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1004), .A2(new_n1011), .A3(new_n1005), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1100), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1032), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT125), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(G390), .A2(new_n1036), .A3(new_n985), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT125), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1032), .A2(new_n1297), .A3(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1299), .A2(new_n1300), .A3(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(new_n816), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1297), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1032), .A2(new_n1297), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(new_n1304), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1303), .A2(new_n1304), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT126), .B1(new_n1308), .B2(KEYINPUT61), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1302), .A2(new_n1300), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1301), .B1(new_n1032), .B2(new_n1297), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1304), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1309), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1293), .A2(new_n1295), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1314), .A2(KEYINPUT127), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1314), .A2(KEYINPUT127), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1289), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1316), .B1(new_n1291), .B2(KEYINPUT62), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1320), .B(new_n1321), .C1(new_n1323), .C2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1319), .A2(new_n1325), .ZN(G405));
  INV_X1    g1126(.A(new_n1268), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1290), .B1(new_n1262), .B2(new_n1327), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1261), .B(new_n1268), .C1(new_n1280), .C2(new_n1279), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1314), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1328), .A2(new_n1308), .A3(new_n1329), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(G402));
endmodule


