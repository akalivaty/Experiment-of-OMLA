

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U553 ( .A(n656), .B(KEYINPUT91), .ZN(n694) );
  NOR2_X2 U554 ( .A1(n603), .A2(n710), .ZN(n651) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n711) );
  XOR2_X1 U556 ( .A(n759), .B(KEYINPUT105), .Z(n516) );
  AND2_X1 U557 ( .A1(n762), .A2(n761), .ZN(n517) );
  NOR2_X1 U558 ( .A1(n969), .A2(n632), .ZN(n633) );
  INV_X1 U559 ( .A(KEYINPUT97), .ZN(n641) );
  XNOR2_X1 U560 ( .A(n642), .B(n641), .ZN(n645) );
  NAND2_X1 U561 ( .A1(n645), .A2(n644), .ZN(n646) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n648) );
  XNOR2_X1 U563 ( .A(n649), .B(n648), .ZN(n655) );
  NAND2_X1 U564 ( .A1(n655), .A2(n654), .ZN(n682) );
  NOR2_X1 U565 ( .A1(G1966), .A2(n742), .ZN(n684) );
  NAND2_X1 U566 ( .A1(G160), .A2(G40), .ZN(n710) );
  NOR2_X1 U567 ( .A1(n518), .A2(G2105), .ZN(n519) );
  AND2_X1 U568 ( .A1(n760), .A2(n516), .ZN(n761) );
  NOR2_X1 U569 ( .A1(G651), .A2(n593), .ZN(n779) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n876) );
  NAND2_X1 U571 ( .A1(n876), .A2(G113), .ZN(n522) );
  INV_X1 U572 ( .A(G2104), .ZN(n518) );
  XNOR2_X2 U573 ( .A(n519), .B(KEYINPUT64), .ZN(n880) );
  NAND2_X1 U574 ( .A1(n880), .A2(G101), .ZN(n520) );
  XOR2_X1 U575 ( .A(n520), .B(KEYINPUT23), .Z(n521) );
  NAND2_X1 U576 ( .A1(n522), .A2(n521), .ZN(n527) );
  AND2_X1 U577 ( .A1(n518), .A2(G2105), .ZN(n875) );
  NAND2_X1 U578 ( .A1(G125), .A2(n875), .ZN(n525) );
  NOR2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X2 U580 ( .A(KEYINPUT17), .B(n523), .Z(n883) );
  NAND2_X1 U581 ( .A1(G137), .A2(n883), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X2 U583 ( .A1(n527), .A2(n526), .ZN(G160) );
  NAND2_X1 U584 ( .A1(G138), .A2(n883), .ZN(n529) );
  NAND2_X1 U585 ( .A1(G102), .A2(n880), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G126), .A2(n875), .ZN(n531) );
  NAND2_X1 U588 ( .A1(G114), .A2(n876), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U590 ( .A1(n533), .A2(n532), .ZN(G164) );
  XNOR2_X1 U591 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U592 ( .A(G651), .ZN(n537) );
  NOR2_X1 U593 ( .A1(G543), .A2(n537), .ZN(n534) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n534), .Z(n778) );
  NAND2_X1 U595 ( .A1(G60), .A2(n778), .ZN(n536) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n783) );
  NAND2_X1 U597 ( .A1(G85), .A2(n783), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n541) );
  XOR2_X1 U599 ( .A(G543), .B(KEYINPUT0), .Z(n593) );
  NOR2_X1 U600 ( .A1(n593), .A2(n537), .ZN(n787) );
  NAND2_X1 U601 ( .A1(G72), .A2(n787), .ZN(n539) );
  NAND2_X1 U602 ( .A1(G47), .A2(n779), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U604 ( .A1(n541), .A2(n540), .ZN(G290) );
  NAND2_X1 U605 ( .A1(G78), .A2(n787), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(KEYINPUT68), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G65), .A2(n778), .ZN(n544) );
  NAND2_X1 U608 ( .A1(G91), .A2(n783), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U610 ( .A1(G53), .A2(n779), .ZN(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT69), .B(n545), .ZN(n546) );
  NOR2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U614 ( .A(KEYINPUT70), .B(n550), .Z(n793) );
  INV_X1 U615 ( .A(n793), .ZN(G299) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U617 ( .A1(G123), .A2(n875), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(KEYINPUT18), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G111), .A2(n876), .ZN(n553) );
  NAND2_X1 U620 ( .A1(G135), .A2(n883), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U622 ( .A1(G99), .A2(n880), .ZN(n554) );
  XNOR2_X1 U623 ( .A(KEYINPUT77), .B(n554), .ZN(n555) );
  NOR2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n927) );
  XNOR2_X1 U626 ( .A(G2096), .B(n927), .ZN(n559) );
  OR2_X1 U627 ( .A1(G2100), .A2(n559), .ZN(G156) );
  NAND2_X1 U628 ( .A1(n778), .A2(G64), .ZN(n560) );
  XNOR2_X1 U629 ( .A(KEYINPUT65), .B(n560), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n787), .A2(G77), .ZN(n561) );
  XNOR2_X1 U631 ( .A(n561), .B(KEYINPUT66), .ZN(n563) );
  NAND2_X1 U632 ( .A1(G90), .A2(n783), .ZN(n562) );
  NAND2_X1 U633 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U634 ( .A(KEYINPUT67), .B(n564), .Z(n565) );
  XNOR2_X1 U635 ( .A(n565), .B(KEYINPUT9), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G52), .A2(n779), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U638 ( .A1(n569), .A2(n568), .ZN(G171) );
  INV_X1 U639 ( .A(G171), .ZN(G301) );
  INV_X1 U640 ( .A(G132), .ZN(G219) );
  INV_X1 U641 ( .A(G57), .ZN(G237) );
  NAND2_X1 U642 ( .A1(G89), .A2(n783), .ZN(n570) );
  XOR2_X1 U643 ( .A(KEYINPUT75), .B(n570), .Z(n571) );
  XNOR2_X1 U644 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U645 ( .A1(G76), .A2(n787), .ZN(n572) );
  NAND2_X1 U646 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U647 ( .A(n574), .B(KEYINPUT5), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G63), .A2(n778), .ZN(n576) );
  NAND2_X1 U649 ( .A1(G51), .A2(n779), .ZN(n575) );
  NAND2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U651 ( .A(KEYINPUT6), .B(n577), .Z(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U653 ( .A(n580), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U654 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U655 ( .A1(n787), .A2(G75), .ZN(n583) );
  NAND2_X1 U656 ( .A1(G88), .A2(n783), .ZN(n581) );
  XOR2_X1 U657 ( .A(KEYINPUT83), .B(n581), .Z(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G62), .A2(n778), .ZN(n585) );
  NAND2_X1 U660 ( .A1(G50), .A2(n779), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U662 ( .A1(n587), .A2(n586), .ZN(G166) );
  XNOR2_X1 U663 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  NAND2_X1 U664 ( .A1(G651), .A2(G74), .ZN(n588) );
  XOR2_X1 U665 ( .A(KEYINPUT81), .B(n588), .Z(n590) );
  NAND2_X1 U666 ( .A1(n779), .A2(G49), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U668 ( .A(KEYINPUT82), .B(n591), .ZN(n592) );
  NOR2_X1 U669 ( .A1(n778), .A2(n592), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n593), .A2(G87), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(G288) );
  NAND2_X1 U672 ( .A1(G61), .A2(n778), .ZN(n597) );
  NAND2_X1 U673 ( .A1(G48), .A2(n779), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G73), .A2(n787), .ZN(n598) );
  XOR2_X1 U676 ( .A(KEYINPUT2), .B(n598), .Z(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n783), .A2(G86), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(G305) );
  INV_X1 U680 ( .A(n711), .ZN(n603) );
  INV_X1 U681 ( .A(n651), .ZN(n664) );
  NAND2_X1 U682 ( .A1(G1956), .A2(n664), .ZN(n604) );
  XNOR2_X1 U683 ( .A(KEYINPUT95), .B(n604), .ZN(n608) );
  XOR2_X1 U684 ( .A(KEYINPUT27), .B(KEYINPUT94), .Z(n606) );
  NAND2_X1 U685 ( .A1(n651), .A2(G2072), .ZN(n605) );
  XOR2_X1 U686 ( .A(n606), .B(n605), .Z(n607) );
  NOR2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n643) );
  NOR2_X1 U688 ( .A1(n643), .A2(n793), .ZN(n609) );
  XOR2_X1 U689 ( .A(n609), .B(KEYINPUT28), .Z(n647) );
  NAND2_X1 U690 ( .A1(G54), .A2(n779), .ZN(n610) );
  XNOR2_X1 U691 ( .A(n610), .B(KEYINPUT74), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G79), .A2(n787), .ZN(n612) );
  NAND2_X1 U693 ( .A1(G92), .A2(n783), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U695 ( .A1(G66), .A2(n778), .ZN(n613) );
  XNOR2_X1 U696 ( .A(KEYINPUT73), .B(n613), .ZN(n614) );
  NOR2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U699 ( .A(KEYINPUT15), .B(n618), .Z(n766) );
  INV_X1 U700 ( .A(n766), .ZN(n967) );
  NAND2_X1 U701 ( .A1(G56), .A2(n778), .ZN(n619) );
  XOR2_X1 U702 ( .A(KEYINPUT14), .B(n619), .Z(n626) );
  NAND2_X1 U703 ( .A1(G81), .A2(n783), .ZN(n620) );
  XNOR2_X1 U704 ( .A(n620), .B(KEYINPUT12), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n621), .B(KEYINPUT72), .ZN(n623) );
  NAND2_X1 U706 ( .A1(G68), .A2(n787), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U708 ( .A(KEYINPUT13), .B(n624), .Z(n625) );
  NOR2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n779), .A2(G43), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n969) );
  AND2_X1 U712 ( .A1(n651), .A2(G1996), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n629), .B(KEYINPUT26), .ZN(n631) );
  AND2_X1 U714 ( .A1(n664), .A2(G1341), .ZN(n630) );
  OR2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n632) );
  OR2_X1 U716 ( .A1(n967), .A2(n633), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n967), .A2(n633), .ZN(n638) );
  INV_X1 U718 ( .A(G2067), .ZN(n842) );
  NOR2_X1 U719 ( .A1(n664), .A2(n842), .ZN(n634) );
  XOR2_X1 U720 ( .A(n634), .B(KEYINPUT96), .Z(n636) );
  NAND2_X1 U721 ( .A1(n664), .A2(G1348), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n793), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n649) );
  NOR2_X1 U727 ( .A1(n651), .A2(G1961), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n650), .B(KEYINPUT93), .ZN(n653) );
  XNOR2_X1 U729 ( .A(G2078), .B(KEYINPUT25), .ZN(n948) );
  NAND2_X1 U730 ( .A1(n651), .A2(n948), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n669) );
  NAND2_X1 U732 ( .A1(n669), .A2(G171), .ZN(n654) );
  INV_X1 U733 ( .A(G8), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n664), .A2(G8), .ZN(n656) );
  INV_X1 U735 ( .A(n694), .ZN(n742) );
  NOR2_X1 U736 ( .A1(G1971), .A2(n742), .ZN(n657) );
  XOR2_X1 U737 ( .A(KEYINPUT99), .B(n657), .Z(n659) );
  NOR2_X1 U738 ( .A1(G2090), .A2(n664), .ZN(n658) );
  NOR2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n660), .A2(G303), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n661), .B(KEYINPUT100), .ZN(n662) );
  OR2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n674) );
  AND2_X1 U743 ( .A1(n682), .A2(n674), .ZN(n673) );
  NOR2_X1 U744 ( .A1(G2084), .A2(n664), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n684), .A2(n685), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G8), .A2(n665), .ZN(n666) );
  XNOR2_X1 U747 ( .A(n666), .B(KEYINPUT30), .ZN(n667) );
  NOR2_X1 U748 ( .A1(G168), .A2(n667), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n668), .B(KEYINPUT98), .ZN(n671) );
  NOR2_X1 U750 ( .A1(n669), .A2(G171), .ZN(n670) );
  NOR2_X1 U751 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U752 ( .A(KEYINPUT31), .B(n672), .Z(n681) );
  NAND2_X1 U753 ( .A1(n673), .A2(n681), .ZN(n678) );
  INV_X1 U754 ( .A(n674), .ZN(n676) );
  AND2_X1 U755 ( .A1(G286), .A2(G8), .ZN(n675) );
  OR2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U757 ( .A1(n678), .A2(n677), .ZN(n680) );
  XOR2_X1 U758 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n679) );
  XNOR2_X1 U759 ( .A(n680), .B(n679), .ZN(n689) );
  AND2_X1 U760 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U761 ( .A1(n684), .A2(n683), .ZN(n687) );
  NAND2_X1 U762 ( .A1(G8), .A2(n685), .ZN(n686) );
  NAND2_X1 U763 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U764 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U765 ( .A(KEYINPUT102), .B(n690), .Z(n734) );
  NOR2_X1 U766 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NOR2_X1 U767 ( .A1(G1971), .A2(G303), .ZN(n691) );
  NOR2_X1 U768 ( .A1(n974), .A2(n691), .ZN(n692) );
  XNOR2_X1 U769 ( .A(n692), .B(KEYINPUT103), .ZN(n693) );
  NOR2_X1 U770 ( .A1(n734), .A2(n693), .ZN(n696) );
  NAND2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n975) );
  NAND2_X1 U772 ( .A1(n975), .A2(n694), .ZN(n695) );
  NOR2_X1 U773 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U774 ( .A1(KEYINPUT33), .A2(n697), .ZN(n700) );
  NAND2_X1 U775 ( .A1(n974), .A2(KEYINPUT33), .ZN(n698) );
  NOR2_X1 U776 ( .A1(n742), .A2(n698), .ZN(n699) );
  NOR2_X1 U777 ( .A1(n700), .A2(n699), .ZN(n732) );
  XOR2_X1 U778 ( .A(G1981), .B(G305), .Z(n983) );
  NAND2_X1 U779 ( .A1(G140), .A2(n883), .ZN(n702) );
  NAND2_X1 U780 ( .A1(G104), .A2(n880), .ZN(n701) );
  NAND2_X1 U781 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U782 ( .A(KEYINPUT34), .B(n703), .ZN(n708) );
  NAND2_X1 U783 ( .A1(G128), .A2(n875), .ZN(n705) );
  NAND2_X1 U784 ( .A1(G116), .A2(n876), .ZN(n704) );
  NAND2_X1 U785 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U786 ( .A(KEYINPUT35), .B(n706), .Z(n707) );
  NOR2_X1 U787 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U788 ( .A(KEYINPUT36), .B(n709), .ZN(n893) );
  XOR2_X1 U789 ( .A(n842), .B(KEYINPUT37), .Z(n748) );
  NOR2_X1 U790 ( .A1(n893), .A2(n748), .ZN(n926) );
  NOR2_X1 U791 ( .A1(n711), .A2(n710), .ZN(n758) );
  NAND2_X1 U792 ( .A1(n926), .A2(n758), .ZN(n754) );
  NAND2_X1 U793 ( .A1(G119), .A2(n875), .ZN(n713) );
  NAND2_X1 U794 ( .A1(G107), .A2(n876), .ZN(n712) );
  NAND2_X1 U795 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U796 ( .A1(G131), .A2(n883), .ZN(n715) );
  NAND2_X1 U797 ( .A1(G95), .A2(n880), .ZN(n714) );
  NAND2_X1 U798 ( .A1(n715), .A2(n714), .ZN(n716) );
  OR2_X1 U799 ( .A1(n717), .A2(n716), .ZN(n863) );
  NAND2_X1 U800 ( .A1(G1991), .A2(n863), .ZN(n727) );
  NAND2_X1 U801 ( .A1(G129), .A2(n875), .ZN(n719) );
  NAND2_X1 U802 ( .A1(G117), .A2(n876), .ZN(n718) );
  NAND2_X1 U803 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U804 ( .A1(G105), .A2(n880), .ZN(n720) );
  XOR2_X1 U805 ( .A(KEYINPUT38), .B(n720), .Z(n721) );
  NOR2_X1 U806 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U807 ( .A(n723), .B(KEYINPUT90), .ZN(n725) );
  NAND2_X1 U808 ( .A1(G141), .A2(n883), .ZN(n724) );
  NAND2_X1 U809 ( .A1(n725), .A2(n724), .ZN(n892) );
  NAND2_X1 U810 ( .A1(G1996), .A2(n892), .ZN(n726) );
  NAND2_X1 U811 ( .A1(n727), .A2(n726), .ZN(n941) );
  INV_X1 U812 ( .A(n941), .ZN(n728) );
  XOR2_X1 U813 ( .A(G1986), .B(G290), .Z(n972) );
  NAND2_X1 U814 ( .A1(n728), .A2(n972), .ZN(n729) );
  NAND2_X1 U815 ( .A1(n758), .A2(n729), .ZN(n730) );
  NAND2_X1 U816 ( .A1(n754), .A2(n730), .ZN(n745) );
  INV_X1 U817 ( .A(n745), .ZN(n737) );
  AND2_X1 U818 ( .A1(n983), .A2(n737), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n762) );
  NOR2_X1 U820 ( .A1(G2090), .A2(G303), .ZN(n733) );
  NAND2_X1 U821 ( .A1(G8), .A2(n733), .ZN(n736) );
  INV_X1 U822 ( .A(n734), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n739) );
  AND2_X1 U824 ( .A1(n742), .A2(n737), .ZN(n738) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n747) );
  NOR2_X1 U826 ( .A1(G1981), .A2(G305), .ZN(n740) );
  XOR2_X1 U827 ( .A(n740), .B(KEYINPUT24), .Z(n741) );
  NOR2_X1 U828 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U829 ( .A(n743), .B(KEYINPUT92), .Z(n744) );
  OR2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U831 ( .A1(n747), .A2(n746), .ZN(n760) );
  NAND2_X1 U832 ( .A1(n893), .A2(n748), .ZN(n931) );
  NOR2_X1 U833 ( .A1(G1996), .A2(n892), .ZN(n934) );
  NOR2_X1 U834 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U835 ( .A1(G1991), .A2(n863), .ZN(n749) );
  XNOR2_X1 U836 ( .A(KEYINPUT104), .B(n749), .ZN(n930) );
  NOR2_X1 U837 ( .A1(n750), .A2(n930), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n751), .A2(n941), .ZN(n752) );
  NOR2_X1 U839 ( .A1(n934), .A2(n752), .ZN(n753) );
  XNOR2_X1 U840 ( .A(n753), .B(KEYINPUT39), .ZN(n755) );
  NAND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n931), .A2(n756), .ZN(n757) );
  NAND2_X1 U843 ( .A1(n758), .A2(n757), .ZN(n759) );
  INV_X1 U844 ( .A(KEYINPUT40), .ZN(n763) );
  XNOR2_X1 U845 ( .A(n517), .B(n763), .ZN(G329) );
  NAND2_X1 U846 ( .A1(G7), .A2(G661), .ZN(n764) );
  XOR2_X1 U847 ( .A(n764), .B(KEYINPUT10), .Z(n918) );
  NAND2_X1 U848 ( .A1(n918), .A2(G567), .ZN(n765) );
  XOR2_X1 U849 ( .A(KEYINPUT11), .B(n765), .Z(G234) );
  INV_X1 U850 ( .A(G860), .ZN(n772) );
  OR2_X1 U851 ( .A1(n969), .A2(n772), .ZN(G153) );
  NAND2_X1 U852 ( .A1(G868), .A2(G301), .ZN(n768) );
  INV_X1 U853 ( .A(G868), .ZN(n802) );
  NAND2_X1 U854 ( .A1(n766), .A2(n802), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(G284) );
  XOR2_X1 U856 ( .A(KEYINPUT76), .B(G868), .Z(n769) );
  NOR2_X1 U857 ( .A1(G286), .A2(n769), .ZN(n771) );
  NOR2_X1 U858 ( .A1(G299), .A2(G868), .ZN(n770) );
  NOR2_X1 U859 ( .A1(n771), .A2(n770), .ZN(G297) );
  NAND2_X1 U860 ( .A1(n772), .A2(G559), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n773), .A2(n967), .ZN(n774) );
  XNOR2_X1 U862 ( .A(n774), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U863 ( .A1(G868), .A2(n969), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G868), .A2(n967), .ZN(n775) );
  NOR2_X1 U865 ( .A1(G559), .A2(n775), .ZN(n776) );
  NOR2_X1 U866 ( .A1(n777), .A2(n776), .ZN(G282) );
  NAND2_X1 U867 ( .A1(G67), .A2(n778), .ZN(n781) );
  NAND2_X1 U868 ( .A1(G55), .A2(n779), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U870 ( .A(KEYINPUT80), .B(n782), .ZN(n786) );
  NAND2_X1 U871 ( .A1(G93), .A2(n783), .ZN(n784) );
  XNOR2_X1 U872 ( .A(KEYINPUT79), .B(n784), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n787), .A2(G80), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n803) );
  XNOR2_X1 U876 ( .A(n969), .B(KEYINPUT78), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n967), .A2(G559), .ZN(n790) );
  XNOR2_X1 U878 ( .A(n791), .B(n790), .ZN(n800) );
  NOR2_X1 U879 ( .A1(n800), .A2(G860), .ZN(n792) );
  XOR2_X1 U880 ( .A(n803), .B(n792), .Z(G145) );
  XOR2_X1 U881 ( .A(n793), .B(n803), .Z(n799) );
  XNOR2_X1 U882 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n795) );
  XNOR2_X1 U883 ( .A(G288), .B(G166), .ZN(n794) );
  XNOR2_X1 U884 ( .A(n795), .B(n794), .ZN(n796) );
  XOR2_X1 U885 ( .A(n796), .B(G305), .Z(n797) );
  XNOR2_X1 U886 ( .A(G290), .B(n797), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n799), .B(n798), .ZN(n896) );
  XOR2_X1 U888 ( .A(n896), .B(n800), .Z(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n805) );
  NOR2_X1 U890 ( .A1(G868), .A2(n803), .ZN(n804) );
  NOR2_X1 U891 ( .A1(n805), .A2(n804), .ZN(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n806) );
  XOR2_X1 U893 ( .A(KEYINPUT20), .B(n806), .Z(n807) );
  NAND2_X1 U894 ( .A1(G2090), .A2(n807), .ZN(n808) );
  XNOR2_X1 U895 ( .A(KEYINPUT21), .B(n808), .ZN(n809) );
  NAND2_X1 U896 ( .A1(n809), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U897 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NAND2_X1 U898 ( .A1(G120), .A2(G69), .ZN(n810) );
  XNOR2_X1 U899 ( .A(KEYINPUT86), .B(n810), .ZN(n811) );
  NOR2_X1 U900 ( .A1(G237), .A2(n811), .ZN(n812) );
  NAND2_X1 U901 ( .A1(G108), .A2(n812), .ZN(n826) );
  NAND2_X1 U902 ( .A1(G567), .A2(n826), .ZN(n813) );
  XNOR2_X1 U903 ( .A(n813), .B(KEYINPUT87), .ZN(n819) );
  NOR2_X1 U904 ( .A1(G219), .A2(G220), .ZN(n814) );
  XOR2_X1 U905 ( .A(KEYINPUT85), .B(n814), .Z(n815) );
  XNOR2_X1 U906 ( .A(KEYINPUT22), .B(n815), .ZN(n816) );
  NAND2_X1 U907 ( .A1(n816), .A2(G96), .ZN(n817) );
  OR2_X1 U908 ( .A1(G218), .A2(n817), .ZN(n827) );
  AND2_X1 U909 ( .A1(G2106), .A2(n827), .ZN(n818) );
  NOR2_X1 U910 ( .A1(n819), .A2(n818), .ZN(G319) );
  INV_X1 U911 ( .A(G319), .ZN(n822) );
  NAND2_X1 U912 ( .A1(G661), .A2(G483), .ZN(n820) );
  XNOR2_X1 U913 ( .A(KEYINPUT88), .B(n820), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n918), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U918 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(G188) );
  XOR2_X1 U921 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  XNOR2_X1 U922 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  NOR2_X1 U926 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XOR2_X1 U928 ( .A(KEYINPUT112), .B(G1986), .Z(n829) );
  XNOR2_X1 U929 ( .A(G1956), .B(G1971), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U931 ( .A(n830), .B(G2474), .Z(n833) );
  INV_X1 U932 ( .A(G1996), .ZN(n831) );
  XOR2_X1 U933 ( .A(n831), .B(G1991), .Z(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U935 ( .A(G1961), .B(G1966), .Z(n835) );
  XNOR2_X1 U936 ( .A(G1981), .B(G1976), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U938 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U939 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(G229) );
  XOR2_X1 U941 ( .A(KEYINPUT109), .B(G2678), .Z(n841) );
  XNOR2_X1 U942 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n846) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2090), .Z(n844) );
  XOR2_X1 U945 ( .A(n842), .B(G2072), .Z(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U947 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2096), .B(G2100), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n850) );
  XOR2_X1 U950 ( .A(G2078), .B(G2084), .Z(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(G227) );
  NAND2_X1 U952 ( .A1(n880), .A2(G100), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n851), .B(KEYINPUT114), .ZN(n854) );
  NAND2_X1 U954 ( .A1(G136), .A2(n883), .ZN(n852) );
  XOR2_X1 U955 ( .A(KEYINPUT113), .B(n852), .Z(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n875), .A2(G124), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G112), .A2(n876), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U961 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U962 ( .A(KEYINPUT118), .B(KEYINPUT116), .Z(n861) );
  XNOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n865) );
  XNOR2_X1 U966 ( .A(G164), .B(G160), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n890) );
  NAND2_X1 U968 ( .A1(G130), .A2(n875), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G118), .A2(n876), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G142), .A2(n883), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G106), .A2(n880), .ZN(n868) );
  NAND2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U974 ( .A(KEYINPUT115), .B(n870), .ZN(n871) );
  XNOR2_X1 U975 ( .A(KEYINPUT45), .B(n871), .ZN(n872) );
  NOR2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n927), .B(n874), .ZN(n888) );
  NAND2_X1 U978 ( .A1(G127), .A2(n875), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G115), .A2(n876), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n879), .B(KEYINPUT47), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G103), .A2(n880), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G139), .A2(n883), .ZN(n884) );
  XNOR2_X1 U985 ( .A(KEYINPUT117), .B(n884), .ZN(n885) );
  NOR2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n919) );
  XNOR2_X1 U987 ( .A(G162), .B(n919), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(n890), .B(n889), .Z(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n894) );
  XOR2_X1 U991 ( .A(n894), .B(n893), .Z(n895) );
  NOR2_X1 U992 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n969), .B(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(G301), .B(n967), .Z(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n899), .B(G286), .ZN(n900) );
  NOR2_X1 U997 ( .A1(G37), .A2(n900), .ZN(G397) );
  XNOR2_X1 U998 ( .A(G2427), .B(KEYINPUT107), .ZN(n910) );
  XOR2_X1 U999 ( .A(G2443), .B(G2438), .Z(n902) );
  XNOR2_X1 U1000 ( .A(KEYINPUT106), .B(G2454), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1002 ( .A(G2430), .B(G2435), .Z(n904) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U1006 ( .A(G2451), .B(G2446), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n911), .A2(G14), .ZN(n917) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n917), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n917), .ZN(G401) );
  INV_X1 U1018 ( .A(n918), .ZN(G223) );
  XOR2_X1 U1019 ( .A(G2072), .B(n919), .Z(n920) );
  XNOR2_X1 U1020 ( .A(KEYINPUT120), .B(n920), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(G2078), .B(G164), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(KEYINPUT121), .B(n921), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1024 ( .A(KEYINPUT50), .B(n924), .Z(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n939) );
  XNOR2_X1 U1026 ( .A(G160), .B(G2084), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n937) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT51), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n942), .ZN(n943) );
  XOR2_X1 U1037 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n963) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n963), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n958) );
  XOR2_X1 U1041 ( .A(G32), .B(G1996), .Z(n945) );
  NAND2_X1 U1042 ( .A1(n945), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G2072), .B(G33), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(G1991), .B(G25), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n952) );
  XOR2_X1 U1046 ( .A(n948), .B(G27), .Z(n950) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G26), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1051 ( .A(KEYINPUT53), .B(n955), .Z(n956) );
  XNOR2_X1 U1052 ( .A(n956), .B(KEYINPUT123), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1058 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n966), .ZN(n1020) );
  INV_X1 U1061 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1062 ( .A(n1016), .B(KEYINPUT56), .Z(n993) );
  XNOR2_X1 U1063 ( .A(G1348), .B(KEYINPUT124), .ZN(n968) );
  XOR2_X1 U1064 ( .A(n968), .B(n967), .Z(n971) );
  XNOR2_X1 U1065 ( .A(G1341), .B(n969), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n991) );
  XOR2_X1 U1067 ( .A(G299), .B(G1956), .Z(n981) );
  XOR2_X1 U1068 ( .A(G303), .B(G1971), .Z(n973) );
  NAND2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n979) );
  INV_X1 U1070 ( .A(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1072 ( .A(KEYINPUT125), .B(n977), .Z(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(KEYINPUT126), .ZN(n989) );
  XOR2_X1 U1076 ( .A(G301), .B(G1961), .Z(n987) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n985), .B(KEYINPUT57), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n1018) );
  XNOR2_X1 U1084 ( .A(KEYINPUT127), .B(G1961), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(n994), .B(G5), .ZN(n1011) );
  XOR2_X1 U1086 ( .A(G1348), .B(KEYINPUT59), .Z(n995) );
  XNOR2_X1 U1087 ( .A(G4), .B(n995), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(G20), .B(G1956), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G1981), .B(G6), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(n1002), .B(KEYINPUT60), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G1976), .B(G23), .ZN(n1004) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1003) );
  NOR2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XOR2_X1 U1098 ( .A(G1986), .B(G24), .Z(n1005) );
  NAND2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(G21), .B(G1966), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1023), .ZN(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

