

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U324 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U325 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U326 ( .A(n400), .B(G36GAT), .ZN(n401) );
  XNOR2_X1 U327 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U328 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n470) );
  XNOR2_X1 U329 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U330 ( .A(n471), .B(n470), .ZN(n517) );
  XOR2_X1 U331 ( .A(n411), .B(n410), .Z(n506) );
  XNOR2_X1 U332 ( .A(n452), .B(G190GAT), .ZN(n453) );
  XNOR2_X1 U333 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U334 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XNOR2_X1 U335 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  XOR2_X1 U336 ( .A(G43GAT), .B(G29GAT), .Z(n293) );
  XNOR2_X1 U337 ( .A(KEYINPUT70), .B(G50GAT), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U339 ( .A(n294), .B(KEYINPUT8), .Z(n296) );
  XNOR2_X1 U340 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n333) );
  XOR2_X1 U342 ( .A(KEYINPUT64), .B(KEYINPUT77), .Z(n298) );
  XNOR2_X1 U343 ( .A(KEYINPUT9), .B(KEYINPUT66), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n333), .B(n299), .ZN(n308) );
  XOR2_X1 U346 ( .A(G92GAT), .B(G85GAT), .Z(n301) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G106GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n346) );
  XOR2_X1 U349 ( .A(G190GAT), .B(G134GAT), .Z(n309) );
  XOR2_X1 U350 ( .A(n346), .B(n309), .Z(n303) );
  NAND2_X1 U351 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U353 ( .A(n304), .B(KEYINPUT11), .Z(n306) );
  XOR2_X1 U354 ( .A(G218GAT), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U355 ( .A(n415), .B(KEYINPUT10), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n557) );
  XOR2_X1 U358 ( .A(KEYINPUT78), .B(n557), .Z(n542) );
  XOR2_X1 U359 ( .A(G120GAT), .B(G71GAT), .Z(n354) );
  XNOR2_X1 U360 ( .A(n309), .B(n354), .ZN(n312) );
  XOR2_X1 U361 ( .A(G127GAT), .B(KEYINPUT0), .Z(n311) );
  XNOR2_X1 U362 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n438) );
  XNOR2_X1 U364 ( .A(n312), .B(n438), .ZN(n318) );
  XOR2_X1 U365 ( .A(G183GAT), .B(KEYINPUT17), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n399) );
  XOR2_X1 U368 ( .A(G15GAT), .B(n399), .Z(n316) );
  NAND2_X1 U369 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U371 ( .A(n318), .B(n317), .Z(n326) );
  XOR2_X1 U372 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n320) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(G99GAT), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U375 ( .A(G176GAT), .B(KEYINPUT85), .Z(n322) );
  XNOR2_X1 U376 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n532) );
  XOR2_X1 U380 ( .A(KEYINPUT72), .B(KEYINPUT68), .Z(n328) );
  NAND2_X1 U381 ( .A1(G229GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U383 ( .A(n329), .B(KEYINPUT29), .Z(n335) );
  XOR2_X1 U384 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n331) );
  XNOR2_X1 U385 ( .A(G197GAT), .B(G113GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n337) );
  XNOR2_X1 U389 ( .A(G15GAT), .B(G1GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n336), .B(KEYINPUT71), .ZN(n364) );
  XOR2_X1 U391 ( .A(n337), .B(n364), .Z(n339) );
  XOR2_X1 U392 ( .A(G141GAT), .B(G22GAT), .Z(n416) );
  XOR2_X1 U393 ( .A(G169GAT), .B(G8GAT), .Z(n395) );
  XNOR2_X1 U394 ( .A(n416), .B(n395), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n576) );
  XOR2_X1 U396 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n341) );
  NAND2_X1 U397 ( .A1(G230GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n343) );
  INV_X1 U399 ( .A(KEYINPUT31), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U401 ( .A(G78GAT), .B(G148GAT), .Z(n345) );
  XNOR2_X1 U402 ( .A(KEYINPUT75), .B(G204GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n425) );
  XNOR2_X1 U404 ( .A(n425), .B(n346), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U406 ( .A(G57GAT), .B(KEYINPUT13), .Z(n360) );
  XNOR2_X1 U407 ( .A(n360), .B(KEYINPUT33), .ZN(n350) );
  INV_X1 U408 ( .A(KEYINPUT76), .ZN(n349) );
  XOR2_X1 U409 ( .A(n354), .B(n353), .Z(n355) );
  XNOR2_X1 U410 ( .A(G176GAT), .B(G64GAT), .ZN(n394) );
  XNOR2_X1 U411 ( .A(n355), .B(n394), .ZN(n386) );
  XNOR2_X1 U412 ( .A(KEYINPUT41), .B(n386), .ZN(n564) );
  INV_X1 U413 ( .A(n564), .ZN(n551) );
  NOR2_X1 U414 ( .A1(n576), .A2(n551), .ZN(n357) );
  XNOR2_X1 U415 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n377) );
  XOR2_X1 U417 ( .A(G78GAT), .B(G211GAT), .Z(n359) );
  XNOR2_X1 U418 ( .A(G183GAT), .B(G71GAT), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n361) );
  XOR2_X1 U420 ( .A(n361), .B(n360), .Z(n363) );
  XNOR2_X1 U421 ( .A(G22GAT), .B(G155GAT), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U423 ( .A(n364), .B(KEYINPUT12), .Z(n366) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U426 ( .A(n368), .B(n367), .Z(n376) );
  XOR2_X1 U427 ( .A(KEYINPUT81), .B(G64GAT), .Z(n370) );
  XNOR2_X1 U428 ( .A(G8GAT), .B(G127GAT), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U430 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n372) );
  XNOR2_X1 U431 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n581) );
  NAND2_X1 U435 ( .A1(n377), .A2(n581), .ZN(n379) );
  INV_X1 U436 ( .A(KEYINPUT116), .ZN(n378) );
  NAND2_X1 U437 ( .A1(n380), .A2(n557), .ZN(n382) );
  XOR2_X1 U438 ( .A(KEYINPUT117), .B(KEYINPUT47), .Z(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n390) );
  XNOR2_X1 U440 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n542), .B(KEYINPUT101), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n383), .B(KEYINPUT36), .ZN(n584) );
  NOR2_X1 U443 ( .A1(n581), .A2(n584), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n388) );
  XOR2_X1 U445 ( .A(n576), .B(KEYINPUT73), .Z(n534) );
  NAND2_X1 U446 ( .A1(n386), .A2(n534), .ZN(n387) );
  NOR2_X1 U447 ( .A1(n388), .A2(n387), .ZN(n389) );
  NOR2_X1 U448 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n391), .B(KEYINPUT48), .ZN(n530) );
  XOR2_X1 U450 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n393) );
  XNOR2_X1 U451 ( .A(G204GAT), .B(KEYINPUT92), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n406) );
  XNOR2_X1 U453 ( .A(n394), .B(G218GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n395), .B(G190GAT), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U456 ( .A(G92GAT), .B(n398), .Z(n404) );
  XOR2_X1 U457 ( .A(n399), .B(KEYINPUT90), .Z(n402) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n411) );
  XOR2_X1 U461 ( .A(KEYINPUT21), .B(KEYINPUT88), .Z(n408) );
  XNOR2_X1 U462 ( .A(KEYINPUT87), .B(G211GAT), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U464 ( .A(G197GAT), .B(n409), .Z(n426) );
  INV_X1 U465 ( .A(n426), .ZN(n410) );
  INV_X1 U466 ( .A(n506), .ZN(n521) );
  NOR2_X1 U467 ( .A1(n530), .A2(n521), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n412), .B(KEYINPUT54), .ZN(n573) );
  XOR2_X1 U469 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n414) );
  XNOR2_X1 U470 ( .A(KEYINPUT86), .B(KEYINPUT23), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n420) );
  XOR2_X1 U472 ( .A(G106GAT), .B(n415), .Z(n418) );
  XNOR2_X1 U473 ( .A(G50GAT), .B(n416), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U475 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U476 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U478 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n423), .B(KEYINPUT3), .ZN(n437) );
  XOR2_X1 U480 ( .A(n424), .B(n437), .Z(n428) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n462) );
  XOR2_X1 U483 ( .A(KEYINPUT1), .B(G57GAT), .Z(n430) );
  XNOR2_X1 U484 ( .A(G1GAT), .B(G120GAT), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n446) );
  XOR2_X1 U486 ( .A(G85GAT), .B(G162GAT), .Z(n432) );
  XNOR2_X1 U487 ( .A(G141GAT), .B(G148GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U489 ( .A(G29GAT), .B(G134GAT), .Z(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n442) );
  XNOR2_X1 U491 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n435), .B(KEYINPUT4), .ZN(n436) );
  XOR2_X1 U493 ( .A(n436), .B(KEYINPUT89), .Z(n440) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n444) );
  NAND2_X1 U497 ( .A1(G225GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n503) );
  INV_X1 U500 ( .A(n503), .ZN(n572) );
  AND2_X1 U501 ( .A1(n462), .A2(n572), .ZN(n447) );
  NAND2_X1 U502 ( .A1(n573), .A2(n447), .ZN(n449) );
  INV_X1 U503 ( .A(KEYINPUT55), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n450) );
  NOR2_X1 U505 ( .A1(n532), .A2(n450), .ZN(n451) );
  XNOR2_X1 U506 ( .A(KEYINPUT122), .B(n451), .ZN(n568) );
  NAND2_X1 U507 ( .A1(n542), .A2(n568), .ZN(n454) );
  XOR2_X1 U508 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n452) );
  XOR2_X1 U509 ( .A(KEYINPUT27), .B(n521), .Z(n464) );
  INV_X1 U510 ( .A(n532), .ZN(n508) );
  NOR2_X1 U511 ( .A1(n508), .A2(n462), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n455), .B(KEYINPUT26), .ZN(n574) );
  NAND2_X1 U513 ( .A1(n464), .A2(n574), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n506), .A2(n508), .ZN(n456) );
  NAND2_X1 U515 ( .A1(n462), .A2(n456), .ZN(n457) );
  XOR2_X1 U516 ( .A(KEYINPUT25), .B(n457), .Z(n458) );
  NAND2_X1 U517 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n460), .A2(n572), .ZN(n461) );
  XNOR2_X1 U519 ( .A(KEYINPUT95), .B(n461), .ZN(n468) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT67), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT28), .ZN(n531) );
  NAND2_X1 U522 ( .A1(n503), .A2(n464), .ZN(n529) );
  NOR2_X1 U523 ( .A1(n531), .A2(n529), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n532), .A2(n465), .ZN(n466) );
  XOR2_X1 U525 ( .A(KEYINPUT94), .B(n466), .Z(n467) );
  NOR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n483) );
  NOR2_X1 U527 ( .A1(n584), .A2(n483), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n581), .A2(n469), .ZN(n471) );
  INV_X1 U529 ( .A(n534), .ZN(n559) );
  AND2_X1 U530 ( .A1(n559), .A2(n386), .ZN(n484) );
  NAND2_X1 U531 ( .A1(n517), .A2(n484), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT103), .ZN(n473) );
  XNOR2_X1 U533 ( .A(KEYINPUT38), .B(n473), .ZN(n498) );
  NAND2_X1 U534 ( .A1(n498), .A2(n503), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n474) );
  XNOR2_X1 U536 ( .A(n474), .B(G29GAT), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(G1328GAT) );
  NAND2_X1 U538 ( .A1(n498), .A2(n508), .ZN(n480) );
  XOR2_X1 U539 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n478) );
  XNOR2_X1 U540 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n477) );
  XOR2_X1 U541 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n487) );
  NOR2_X1 U542 ( .A1(n581), .A2(n542), .ZN(n481) );
  XOR2_X1 U543 ( .A(KEYINPUT16), .B(n481), .Z(n482) );
  NOR2_X1 U544 ( .A1(n483), .A2(n482), .ZN(n501) );
  NAND2_X1 U545 ( .A1(n484), .A2(n501), .ZN(n485) );
  XOR2_X1 U546 ( .A(KEYINPUT96), .B(n485), .Z(n495) );
  NAND2_X1 U547 ( .A1(n495), .A2(n503), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n495), .A2(n506), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n489), .B(KEYINPUT98), .ZN(n490) );
  XNOR2_X1 U552 ( .A(G8GAT), .B(n490), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n492) );
  NAND2_X1 U554 ( .A1(n495), .A2(n508), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n494) );
  XOR2_X1 U556 ( .A(G15GAT), .B(KEYINPUT99), .Z(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U558 ( .A1(n495), .A2(n531), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n506), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT107), .Z(n500) );
  NAND2_X1 U563 ( .A1(n531), .A2(n498), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n505) );
  AND2_X1 U566 ( .A1(n564), .A2(n576), .ZN(n516) );
  NAND2_X1 U567 ( .A1(n501), .A2(n516), .ZN(n502) );
  XOR2_X1 U568 ( .A(KEYINPUT108), .B(n502), .Z(n511) );
  NAND2_X1 U569 ( .A1(n503), .A2(n511), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n511), .A2(n506), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT109), .Z(n510) );
  NAND2_X1 U574 ( .A1(n511), .A2(n508), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U577 ( .A1(n531), .A2(n511), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n515) );
  XOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT111), .Z(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT112), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n572), .A2(n526), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(KEYINPUT113), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U586 ( .A1(n526), .A2(n521), .ZN(n522) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U588 ( .A1(n532), .A2(n526), .ZN(n523) );
  XOR2_X1 U589 ( .A(KEYINPUT114), .B(n523), .Z(n524) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  INV_X1 U591 ( .A(n531), .ZN(n525) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U593 ( .A(G106GAT), .B(n527), .Z(n528) );
  XNOR2_X1 U594 ( .A(KEYINPUT44), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n546) );
  NOR2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n546), .A2(n533), .ZN(n541) );
  NOR2_X1 U598 ( .A1(n534), .A2(n541), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT118), .B(n535), .Z(n536) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n536), .ZN(G1340GAT) );
  NOR2_X1 U601 ( .A1(n551), .A2(n541), .ZN(n538) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NOR2_X1 U604 ( .A1(n581), .A2(n541), .ZN(n539) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(n539), .Z(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  INV_X1 U608 ( .A(n541), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n546), .A2(n574), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n576), .A2(n556), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n551), .A2(n556), .ZN(n552) );
  XOR2_X1 U619 ( .A(n553), .B(n552), .Z(G1345GAT) );
  NOR2_X1 U620 ( .A1(n581), .A2(n556), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NAND2_X1 U625 ( .A1(n568), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(n563), .Z(n566) );
  NAND2_X1 U631 ( .A1(n568), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  INV_X1 U633 ( .A(n581), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n571) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n578) );
  AND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n583) );
  NOR2_X1 U641 ( .A1(n576), .A2(n583), .ZN(n577) );
  XOR2_X1 U642 ( .A(n578), .B(n577), .Z(G1352GAT) );
  NOR2_X1 U643 ( .A1(n386), .A2(n583), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

