//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT92), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n202), .A2(new_n203), .A3(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n202), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G8gat), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n206), .A2(new_n212), .A3(new_n207), .A4(new_n209), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G57gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G64gat), .ZN(new_n216));
  INV_X1    g015(.A(G64gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(G57gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT96), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G71gat), .A2(G78gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(KEYINPUT97), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT97), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n217), .A2(G57gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n215), .A2(G64gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT96), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n219), .A2(new_n222), .A3(new_n225), .A4(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G71gat), .B(G78gat), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT98), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT100), .ZN(new_n234));
  OR2_X1    g033(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n234), .B(new_n226), .C1(new_n237), .C2(new_n217), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n217), .B1(new_n235), .B2(new_n236), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT100), .B1(new_n239), .B2(new_n216), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n225), .A2(new_n222), .ZN(new_n241));
  INV_X1    g040(.A(new_n231), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n238), .A2(new_n240), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT98), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n230), .A2(new_n244), .A3(new_n231), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n233), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT21), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n214), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT102), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n247), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G155gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n249), .B(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G231gat), .A2(G233gat), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n253), .A2(new_n254), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G183gat), .B(G211gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT20), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n261), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT39), .ZN(new_n266));
  XOR2_X1   g065(.A(G141gat), .B(G148gat), .Z(new_n267));
  INV_X1    g066(.A(KEYINPUT76), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT2), .ZN(new_n269));
  INV_X1    g068(.A(G155gat), .ZN(new_n270));
  INV_X1    g069(.A(G162gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n267), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(new_n268), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT79), .B(G155gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G162gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT2), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n271), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n273), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT78), .B(G148gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G141gat), .ZN(new_n283));
  INV_X1    g082(.A(G148gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G141gat), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n285), .A2(KEYINPUT77), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(KEYINPUT77), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n283), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n275), .B1(new_n281), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G120gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(G113gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT68), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n290), .B2(G113gat), .ZN(new_n294));
  INV_X1    g093(.A(G113gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n292), .B(new_n294), .C1(new_n295), .C2(G120gat), .ZN(new_n296));
  XOR2_X1   g095(.A(G127gat), .B(G134gat), .Z(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT1), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n295), .A2(G120gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(new_n291), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n296), .A2(new_n298), .B1(new_n301), .B2(new_n297), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n289), .A2(new_n303), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n277), .A2(KEYINPUT2), .B1(new_n273), .B2(new_n279), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n283), .A2(new_n286), .A3(new_n287), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n305), .A2(new_n306), .B1(new_n272), .B2(new_n274), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n302), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT80), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n266), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n313), .A2(KEYINPUT88), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(KEYINPUT4), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n307), .A2(new_n316), .A3(new_n302), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n302), .B1(new_n289), .B2(KEYINPUT3), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n275), .B(new_n319), .C1(new_n281), .C2(new_n288), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n315), .A2(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n321), .A2(new_n312), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n313), .A2(KEYINPUT88), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n314), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G1gat), .B(G29gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(KEYINPUT0), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(G57gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(G85gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n324), .B(new_n329), .C1(KEYINPUT39), .C2(new_n322), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT40), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT5), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n321), .A2(new_n312), .ZN(new_n333));
  OR2_X1    g132(.A1(new_n309), .A2(new_n312), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT5), .B1(new_n321), .B2(new_n312), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n330), .A2(new_n331), .B1(new_n328), .B2(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n330), .A2(new_n331), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT87), .ZN(new_n340));
  INV_X1    g139(.A(G211gat), .ZN(new_n341));
  INV_X1    g140(.A(G218gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G211gat), .A2(G218gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G197gat), .B(G204gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT22), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n345), .B1(new_n348), .B2(new_n346), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G226gat), .ZN(new_n353));
  INV_X1    g152(.A(G233gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G190gat), .ZN(new_n357));
  AND2_X1   g156(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT27), .B(G183gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(KEYINPUT28), .A3(new_n357), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n364), .A3(KEYINPUT66), .ZN(new_n365));
  NAND2_X1  g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT26), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT67), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n368), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT67), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n372), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n375), .A3(new_n361), .ZN(new_n376));
  NAND2_X1  g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n365), .A2(new_n374), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT24), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(new_n377), .ZN(new_n381));
  NAND3_X1  g180(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n366), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT25), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(KEYINPUT65), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT64), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n382), .A2(new_n390), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n381), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n394), .B(new_n366), .C1(new_n385), .C2(new_n386), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n389), .A2(new_n393), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n388), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT72), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT72), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n378), .A2(new_n400), .A3(new_n388), .A4(new_n397), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n356), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n355), .A2(KEYINPUT29), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n352), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n399), .A2(new_n401), .A3(new_n403), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n397), .A2(new_n388), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n378), .A3(new_n355), .ZN(new_n408));
  INV_X1    g207(.A(new_n352), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G8gat), .B(G36gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(new_n217), .ZN(new_n412));
  INV_X1    g211(.A(G92gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n405), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT73), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n405), .A2(new_n410), .ZN(new_n418));
  INV_X1    g217(.A(new_n414), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(KEYINPUT30), .A3(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n405), .A2(KEYINPUT73), .A3(new_n410), .A4(new_n414), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(KEYINPUT75), .B(KEYINPUT30), .Z(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n418), .B2(new_n419), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n340), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n427), .A2(KEYINPUT87), .A3(new_n424), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n338), .B(new_n339), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT31), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(G50gat), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n433), .B(new_n434), .C1(new_n350), .C2(new_n351), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n319), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n346), .A2(new_n348), .ZN(new_n437));
  INV_X1    g236(.A(new_n345), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT29), .B1(new_n439), .B2(new_n349), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(new_n433), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n289), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n320), .A2(new_n434), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n352), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT83), .B(new_n289), .C1(new_n436), .C2(new_n441), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G228gat), .A2(G233gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI211_X1 g249(.A(KEYINPUT85), .B(KEYINPUT29), .C1(new_n307), .C2(new_n319), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n320), .B2(new_n434), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n352), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n449), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n440), .A2(KEYINPUT3), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(new_n307), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n289), .B(KEYINPUT84), .C1(KEYINPUT3), .C2(new_n440), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(new_n455), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G22gat), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n450), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(new_n450), .B2(new_n460), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n432), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n450), .A2(new_n460), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G22gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n432), .A2(KEYINPUT86), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n460), .A3(new_n461), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(KEYINPUT86), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n464), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n329), .B1(new_n335), .B2(new_n336), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n333), .A2(new_n332), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n309), .A2(new_n312), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n312), .B2(new_n321), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n328), .B(new_n474), .C1(new_n476), .C2(new_n332), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n478), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n337), .A2(new_n328), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n418), .A2(new_n419), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT89), .B(KEYINPUT38), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n419), .B1(new_n418), .B2(new_n485), .ZN(new_n486));
  OR3_X1    g285(.A1(new_n402), .A2(new_n352), .A3(new_n404), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n406), .A2(new_n408), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n487), .B(KEYINPUT37), .C1(new_n409), .C2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n484), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n405), .A2(KEYINPUT37), .A3(new_n410), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n486), .A2(new_n484), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n482), .B(new_n483), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n429), .A2(new_n472), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n427), .A2(KEYINPUT74), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT74), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n417), .A2(new_n420), .A3(new_n496), .A4(new_n421), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n481), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n425), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n407), .A2(new_n501), .A3(new_n302), .A4(new_n378), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n378), .A2(new_n302), .A3(new_n388), .A4(new_n397), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT69), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n398), .A2(new_n303), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT32), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT34), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n507), .B2(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n512), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(KEYINPUT32), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n506), .A2(new_n508), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n514), .B1(new_n509), .B2(KEYINPUT32), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n520));
  AOI211_X1 g319(.A(new_n520), .B(new_n512), .C1(new_n506), .C2(new_n508), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n516), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT33), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G43gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT70), .ZN(new_n527));
  XNOR2_X1  g326(.A(G71gat), .B(G99gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n530), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n518), .A2(new_n522), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(KEYINPUT36), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n518), .A2(new_n522), .A3(new_n532), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n532), .B1(new_n518), .B2(new_n522), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n500), .A2(new_n471), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n494), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n464), .A2(new_n469), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n541), .A2(new_n533), .A3(new_n531), .A4(new_n470), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT35), .B1(new_n500), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n426), .A2(new_n428), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n471), .A2(new_n536), .A3(new_n537), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n499), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G162gat), .B(G218gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G29gat), .ZN(new_n552));
  INV_X1    g351(.A(G36gat), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT14), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(new_n552), .B2(new_n553), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G43gat), .ZN(new_n559));
  INV_X1    g358(.A(G50gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT15), .ZN(new_n562));
  NAND2_X1  g361(.A1(G43gat), .A2(G50gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n563), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT15), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n564), .A2(new_n565), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n558), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n557), .B1(KEYINPUT15), .B2(new_n567), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT17), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT104), .ZN(new_n574));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT7), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(G85gat), .A3(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(G85gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n581), .B2(new_n413), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G99gat), .B(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n574), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n579), .A2(new_n582), .A3(new_n584), .A4(KEYINPUT104), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n570), .A2(new_n568), .A3(new_n566), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n557), .ZN(new_n592));
  INV_X1    g391(.A(new_n572), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT17), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n590), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n571), .A2(new_n572), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n588), .A3(new_n589), .ZN(new_n598));
  NAND3_X1  g397(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n600), .A2(G134gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(G134gat), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n603), .B(KEYINPUT103), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G190gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n601), .B2(new_n602), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n551), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(new_n550), .A3(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT105), .B1(new_n579), .B2(new_n582), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n579), .A2(new_n582), .A3(KEYINPUT105), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n585), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n588), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT106), .B1(new_n246), .B2(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n230), .A2(new_n244), .A3(new_n231), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n244), .B1(new_n230), .B2(new_n231), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT106), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n579), .A2(KEYINPUT105), .A3(new_n582), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n614), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n625), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n622), .A2(new_n623), .A3(new_n243), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT107), .B(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n246), .A2(new_n590), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n619), .A2(new_n627), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n246), .A2(new_n590), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n629), .A3(new_n627), .ZN(new_n636));
  INV_X1    g435(.A(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT108), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  INV_X1    g440(.A(G176gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(G204gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n636), .A2(KEYINPUT108), .A3(new_n637), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n635), .A2(new_n640), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n638), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n637), .B1(new_n630), .B2(new_n632), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n648), .A2(KEYINPUT109), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT109), .B1(new_n648), .B2(new_n651), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n573), .A2(new_n214), .A3(new_n595), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n211), .A2(new_n213), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n597), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G229gat), .A2(G233gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT93), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT18), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT94), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n656), .A2(KEYINPUT18), .A3(new_n658), .A4(new_n661), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n660), .B(KEYINPUT13), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n597), .A2(new_n657), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n597), .A2(new_n657), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT94), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n662), .A2(new_n672), .A3(new_n663), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n665), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT95), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT90), .B(KEYINPUT12), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G113gat), .B(G141gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G197gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT11), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G169gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(G169gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n677), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n680), .A2(G169gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n681), .A3(new_n676), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n674), .A2(new_n675), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n674), .A2(new_n688), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n664), .A2(new_n687), .A3(new_n670), .A4(new_n666), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT95), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n689), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n655), .A2(new_n693), .ZN(new_n694));
  AND4_X1   g493(.A1(new_n265), .A2(new_n549), .A3(new_n613), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n482), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G1gat), .ZN(G1324gat));
  INV_X1    g496(.A(new_n544), .ZN(new_n698));
  NAND2_X1  g497(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n208), .B2(new_n212), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n212), .B1(new_n695), .B2(new_n698), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT42), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(KEYINPUT42), .B2(new_n701), .ZN(G1325gat));
  NOR2_X1   g503(.A1(new_n536), .A2(new_n537), .ZN(new_n705));
  AOI21_X1  g504(.A(G15gat), .B1(new_n695), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n538), .A2(new_n534), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G15gat), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT110), .Z(new_n710));
  AOI21_X1  g509(.A(new_n706), .B1(new_n695), .B2(new_n710), .ZN(G1326gat));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n471), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  AOI21_X1  g513(.A(new_n613), .B1(new_n540), .B2(new_n548), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n264), .A2(new_n694), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n552), .A3(new_n482), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n613), .A2(KEYINPUT44), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n549), .A2(KEYINPUT111), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n540), .A2(new_n548), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n721), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n715), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n716), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT112), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n730), .B(new_n716), .C1(new_n725), .C2(new_n727), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n499), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n719), .B1(new_n732), .B2(new_n552), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT113), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n735), .B(new_n719), .C1(new_n732), .C2(new_n552), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1328gat));
  NAND3_X1  g536(.A1(new_n717), .A2(new_n553), .A3(new_n698), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT46), .Z(new_n739));
  AOI21_X1  g538(.A(new_n544), .B1(new_n729), .B2(new_n731), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n553), .ZN(G1329gat));
  OAI21_X1  g540(.A(G43gat), .B1(new_n728), .B2(new_n707), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n717), .A2(new_n559), .A3(new_n705), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(KEYINPUT47), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n743), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n731), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n708), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n744), .B1(new_n748), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g548(.A(G50gat), .B1(new_n728), .B2(new_n472), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n717), .A2(new_n560), .A3(new_n471), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(KEYINPUT48), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n751), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n746), .A2(new_n471), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(G50gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(new_n755), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g555(.A1(new_n722), .A2(new_n724), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n262), .A2(new_n263), .A3(new_n613), .A4(new_n693), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n655), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n482), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n237), .ZN(G1332gat));
  NOR2_X1   g562(.A1(new_n760), .A2(new_n544), .ZN(new_n764));
  NAND2_X1  g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OR2_X1    g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n764), .B2(new_n766), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT114), .B(KEYINPUT115), .Z(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1333gat));
  NAND3_X1  g569(.A1(new_n761), .A2(G71gat), .A3(new_n708), .ZN(new_n771));
  INV_X1    g570(.A(new_n705), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n760), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(G71gat), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n761), .A2(new_n471), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g576(.A1(new_n725), .A2(new_n727), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n692), .B1(new_n688), .B2(new_n674), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n674), .A2(new_n675), .A3(new_n688), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n778), .A2(new_n265), .A3(new_n654), .A4(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n581), .B1(new_n782), .B2(new_n482), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n265), .A2(new_n781), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n786), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n715), .A2(new_n784), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n655), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n715), .A2(new_n784), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n787), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n794), .A2(G85gat), .A3(new_n499), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT117), .B1(new_n783), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n795), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n725), .A2(new_n727), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n655), .A3(new_n784), .ZN(new_n799));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799), .B2(new_n499), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n797), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n796), .A2(new_n802), .ZN(G1336gat));
  OAI21_X1  g602(.A(new_n413), .B1(new_n794), .B2(new_n544), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT118), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n544), .A2(new_n413), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n798), .A2(new_n655), .A3(new_n784), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n805), .A2(KEYINPUT118), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n809), .B(new_n810), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n799), .B2(new_n707), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n794), .A2(G99gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n772), .B2(new_n813), .ZN(G1338gat));
  INV_X1    g613(.A(G106gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n782), .B2(new_n471), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n794), .A2(G106gat), .A3(new_n472), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT53), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n817), .ZN(new_n819));
  OAI21_X1  g618(.A(G106gat), .B1(new_n799), .B2(new_n472), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n822), .ZN(G1339gat));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n630), .A2(new_n637), .A3(new_n632), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n650), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n633), .A2(new_n828), .A3(new_n634), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n645), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n824), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n646), .B1(new_n650), .B2(new_n828), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n832), .B(KEYINPUT55), .C1(new_n650), .C2(new_n826), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n648), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n613), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n668), .A2(new_n669), .A3(new_n667), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n661), .B1(new_n656), .B2(new_n658), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n681), .B(new_n685), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n691), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n652), .B2(new_n653), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n841), .B(new_n842), .C1(new_n693), .C2(new_n834), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n613), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n833), .A2(new_n648), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n781), .A2(new_n845), .A3(new_n831), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n842), .B1(new_n846), .B2(new_n841), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n840), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n264), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n758), .A2(new_n655), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n542), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n698), .A2(new_n499), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n693), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(new_n295), .ZN(G1340gat));
  OAI21_X1  g655(.A(G120gat), .B1(new_n854), .B2(new_n654), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n654), .A2(G120gat), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT120), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n854), .B2(new_n859), .ZN(G1341gat));
  NOR2_X1   g659(.A1(new_n854), .A2(new_n264), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g661(.A1(new_n854), .A2(new_n613), .ZN(new_n863));
  INV_X1    g662(.A(G134gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT121), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(KEYINPUT56), .A3(new_n868), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n871), .B(new_n872), .C1(new_n864), .C2(new_n863), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n831), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n831), .A2(new_n874), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n845), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n841), .B1(new_n877), .B2(new_n693), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n613), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n265), .B1(new_n879), .B2(new_n840), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n471), .B1(new_n880), .B2(new_n850), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n472), .B1(new_n849), .B2(new_n851), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n853), .A2(new_n707), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G141gat), .B1(new_n888), .B2(new_n693), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n887), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n693), .A2(G141gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT58), .ZN(G1344gat));
  OAI21_X1  g692(.A(KEYINPUT59), .B1(new_n890), .B2(new_n654), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n282), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n472), .A2(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n835), .A2(KEYINPUT123), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n834), .B2(new_n613), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n839), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n265), .B1(new_n879), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n897), .B1(new_n902), .B2(new_n850), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(new_n883), .B2(new_n884), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n904), .A2(new_n654), .A3(new_n886), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n896), .B1(new_n905), .B2(G148gat), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n654), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(KEYINPUT59), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n895), .B1(new_n906), .B2(new_n908), .ZN(G1345gat));
  INV_X1    g708(.A(new_n276), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n888), .A2(new_n910), .A3(new_n264), .ZN(new_n911));
  INV_X1    g710(.A(new_n890), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n276), .B1(new_n912), .B2(new_n265), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n911), .A2(new_n913), .ZN(G1346gat));
  OAI21_X1  g713(.A(G162gat), .B1(new_n888), .B2(new_n613), .ZN(new_n915));
  INV_X1    g714(.A(new_n613), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n271), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n544), .A2(new_n482), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n852), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n693), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(G169gat), .Z(G1348gat));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n654), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n642), .A2(KEYINPUT124), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g724(.A(KEYINPUT124), .B(G176gat), .Z(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n923), .B2(new_n926), .ZN(G1349gat));
  NOR2_X1   g726(.A1(new_n920), .A2(new_n264), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n363), .ZN(new_n929));
  INV_X1    g728(.A(G183gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(new_n928), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT60), .ZN(G1350gat));
  XNOR2_X1  g731(.A(KEYINPUT61), .B(G190gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n920), .A2(new_n613), .ZN(new_n935));
  MUX2_X1   g734(.A(new_n933), .B(new_n934), .S(new_n935), .Z(G1351gat));
  NAND2_X1  g735(.A1(new_n904), .A2(KEYINPUT126), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n707), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n903), .B(new_n940), .C1(new_n883), .C2(new_n884), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n937), .A2(new_n781), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(KEYINPUT125), .B(G197gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n883), .A2(new_n939), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n945), .A2(new_n693), .A3(new_n943), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n944), .A2(KEYINPUT127), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1352gat));
  NOR3_X1   g750(.A1(new_n945), .A2(G204gat), .A3(new_n654), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n937), .A2(new_n939), .A3(new_n941), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(new_n655), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n953), .B1(new_n955), .B2(new_n644), .ZN(G1353gat));
  INV_X1    g755(.A(new_n945), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(new_n341), .A3(new_n265), .ZN(new_n958));
  OR3_X1    g757(.A1(new_n904), .A2(new_n264), .A3(new_n938), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1354gat));
  AOI21_X1  g761(.A(G218gat), .B1(new_n957), .B2(new_n916), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n613), .A2(new_n342), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n954), .B2(new_n964), .ZN(G1355gat));
endmodule


