//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT30), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n209), .B(new_n204), .C1(KEYINPUT22), .C2(new_n207), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT73), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n214), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT74), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(new_n218), .A3(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G226gat), .A2(G233gat), .ZN(new_n222));
  XOR2_X1   g021(.A(new_n222), .B(KEYINPUT75), .Z(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT27), .B(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT28), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(KEYINPUT28), .A3(new_n225), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G169gat), .ZN(new_n231));
  INV_X1    g030(.A(G176gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n233), .A2(KEYINPUT26), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(KEYINPUT26), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(new_n225), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n243));
  MUX2_X1   g042(.A(G183gat), .B(new_n243), .S(G190gat), .Z(new_n244));
  INV_X1    g043(.A(KEYINPUT24), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n237), .B2(new_n225), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n234), .B2(KEYINPUT23), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT23), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n250), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n233), .B1(KEYINPUT23), .B2(new_n234), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n246), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(KEYINPUT65), .B(new_n245), .C1(new_n237), .C2(new_n225), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n244), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n260), .A2(KEYINPUT25), .A3(new_n252), .A4(new_n253), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n230), .A2(KEYINPUT66), .A3(new_n239), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n242), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT29), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n223), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n262), .A2(new_n240), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(new_n222), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n221), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n222), .B1(new_n267), .B2(KEYINPUT29), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n223), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n220), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT76), .ZN(new_n275));
  XOR2_X1   g074(.A(G64gat), .B(G92gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n203), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n273), .B2(new_n277), .ZN(new_n279));
  OR3_X1    g078(.A1(new_n273), .A2(KEYINPUT30), .A3(new_n277), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n282));
  XNOR2_X1  g081(.A(G113gat), .B(G120gat), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n285));
  NOR2_X1   g084(.A1(G127gat), .A2(G134gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G127gat), .A2(G134gat), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT67), .B(G127gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n286), .B1(new_n291), .B2(G134gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT68), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n283), .A2(KEYINPUT1), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n292), .A2(KEYINPUT68), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n290), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G141gat), .ZN(new_n300));
  INV_X1    g099(.A(G141gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G148gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  INV_X1    g103(.A(G155gat), .ZN(new_n305));
  INV_X1    g104(.A(G162gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT77), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n303), .A2(new_n304), .A3(new_n307), .A4(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT78), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(new_n299), .B2(G141gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n301), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n313), .B(new_n314), .C1(new_n301), .C2(G148gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT79), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n304), .B1(new_n308), .B2(KEYINPUT2), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(new_n315), .B2(new_n317), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n311), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n282), .B1(new_n297), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n311), .ZN(new_n323));
  INV_X1    g122(.A(new_n320), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n318), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n283), .A2(KEYINPUT1), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n292), .B2(KEYINPUT68), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(KEYINPUT68), .B2(new_n292), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n325), .A2(new_n328), .A3(KEYINPUT4), .A4(new_n290), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n321), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(KEYINPUT80), .B(new_n311), .C1(new_n319), .C2(new_n320), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(KEYINPUT3), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n335), .B(new_n311), .C1(new_n319), .C2(new_n320), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n297), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n330), .A2(new_n338), .A3(KEYINPUT5), .A4(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n330), .A2(new_n338), .A3(new_n339), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT5), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n332), .A2(new_n333), .A3(new_n297), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n321), .B2(new_n297), .ZN(new_n344));
  INV_X1    g143(.A(new_n339), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n340), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G1gat), .B(G29gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT0), .ZN(new_n351));
  XNOR2_X1  g150(.A(G57gat), .B(G85gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(KEYINPUT85), .B(new_n340), .C1(new_n341), .C2(new_n346), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n349), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n347), .B2(new_n353), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n354), .B(new_n340), .C1(new_n341), .C2(new_n346), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(new_n357), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n202), .B(new_n281), .C1(new_n360), .C2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n356), .B2(new_n359), .ZN(new_n364));
  INV_X1    g163(.A(new_n281), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT87), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n297), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n264), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n297), .A2(new_n242), .A3(new_n262), .A4(new_n263), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n368), .A2(G227gat), .A3(G233gat), .A4(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G15gat), .B(G43gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT33), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(KEYINPUT32), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT70), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n370), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n373), .B1(new_n370), .B2(KEYINPUT32), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n370), .A2(new_n374), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n385));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OR3_X1    g186(.A1(new_n387), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(KEYINPUT34), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT71), .B1(new_n387), .B2(KEYINPUT34), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n390), .A2(new_n389), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n393), .A2(new_n388), .A3(new_n380), .A4(new_n383), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT72), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n384), .A2(KEYINPUT72), .A3(new_n391), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n336), .A2(new_n265), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n217), .A3(new_n219), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n213), .A2(new_n265), .A3(new_n215), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n335), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n332), .A3(new_n333), .ZN(new_n403));
  AND2_X1   g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n211), .A2(new_n212), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT3), .B1(new_n407), .B2(new_n265), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n325), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n404), .B1(new_n400), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(G22gat), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G22gat), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n400), .A2(new_n410), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n413), .B(new_n405), .C1(new_n414), .C2(new_n404), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(G78gat), .B(G106gat), .Z(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT31), .B(G50gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT82), .B(G22gat), .C1(new_n406), .C2(new_n411), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n411), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n412), .A2(KEYINPUT83), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n426), .B(G22gat), .C1(new_n406), .C2(new_n411), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(KEYINPUT35), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n363), .A2(new_n366), .A3(new_n398), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n347), .A2(new_n353), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n361), .A3(new_n357), .ZN(new_n434));
  INV_X1    g233(.A(new_n362), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n281), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n429), .A2(new_n392), .A3(new_n394), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT35), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT88), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n441), .B(KEYINPUT35), .C1(new_n437), .C2(new_n438), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT39), .B1(new_n344), .B2(new_n345), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n339), .B1(new_n330), .B2(new_n338), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n448), .A2(KEYINPUT84), .A3(new_n353), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT84), .B1(new_n448), .B2(new_n353), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT40), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n446), .B(KEYINPUT40), .C1(new_n449), .C2(new_n450), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n365), .A2(new_n453), .A3(new_n356), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n429), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n273), .A2(new_n277), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n273), .A2(KEYINPUT37), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n458), .A2(new_n277), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n220), .B1(new_n266), .B2(new_n268), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n460), .A2(KEYINPUT37), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n270), .A2(new_n221), .A3(new_n271), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT38), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n457), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n364), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n273), .A2(KEYINPUT37), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n465), .A2(KEYINPUT86), .B1(KEYINPUT38), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n464), .A2(new_n364), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n456), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT36), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n396), .A2(new_n472), .A3(new_n397), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT36), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n437), .A2(new_n430), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n443), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G22gat), .ZN(new_n479));
  INV_X1    g278(.A(G1gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT16), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT93), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n479), .B2(G1gat), .ZN(new_n485));
  OAI21_X1  g284(.A(G8gat), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n479), .A2(G1gat), .ZN(new_n487));
  INV_X1    g286(.A(G8gat), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(new_n482), .A3(new_n484), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492));
  OR2_X1    g291(.A1(G43gat), .A2(G50gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(G43gat), .A2(G50gat), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT14), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT14), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(KEYINPUT91), .A2(G36gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(KEYINPUT91), .A2(G36gat), .ZN(new_n504));
  OAI21_X1  g303(.A(G29gat), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n498), .B2(new_n500), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n495), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n492), .A3(new_n494), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n509), .A2(new_n505), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n498), .A2(new_n500), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT17), .B1(new_n514), .B2(KEYINPUT92), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517));
  AOI211_X1 g316(.A(new_n516), .B(new_n517), .C1(new_n508), .C2(new_n513), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n491), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n490), .A2(new_n514), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT18), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n519), .A2(KEYINPUT18), .A3(new_n520), .A4(new_n521), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n511), .A2(KEYINPUT90), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(new_n502), .A3(new_n505), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n527), .A2(new_n495), .B1(new_n510), .B2(new_n512), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n491), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n521), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n520), .B(KEYINPUT13), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n524), .A2(new_n525), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G113gat), .B(G141gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G169gat), .B(G197gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT12), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n532), .A4(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n478), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G57gat), .B(G64gat), .Z(new_n545));
  OR2_X1    g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G57gat), .B(G64gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n547), .B(new_n546), .C1(new_n552), .C2(new_n549), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G99gat), .B(G106gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT7), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G85gat), .ZN(new_n560));
  INV_X1    g359(.A(G92gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT8), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n559), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n556), .A2(new_n557), .ZN(new_n566));
  NAND3_X1  g365(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(KEYINPUT7), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n555), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n563), .B1(new_n560), .B2(new_n561), .ZN(new_n570));
  AND4_X1   g369(.A1(new_n555), .A2(new_n568), .A3(new_n559), .A4(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n554), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT10), .ZN(new_n573));
  INV_X1    g372(.A(new_n555), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n566), .A2(KEYINPUT7), .A3(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n562), .A3(new_n564), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n568), .A2(new_n555), .A3(new_n559), .A4(new_n570), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n577), .A2(new_n553), .A3(new_n551), .A4(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n572), .A2(new_n573), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n569), .A2(new_n571), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n551), .A2(new_n553), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT97), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n579), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(G230gat), .A3(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  NAND4_X1  g393(.A1(new_n587), .A2(new_n589), .A3(new_n591), .A4(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT98), .B1(new_n584), .B2(new_n585), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597));
  INV_X1    g396(.A(new_n585), .ZN(new_n598));
  AOI211_X1 g397(.A(new_n597), .B(new_n598), .C1(new_n580), .C2(new_n583), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n591), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT99), .ZN(new_n601));
  INV_X1    g400(.A(new_n594), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n600), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n595), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(G231gat), .ZN(new_n606));
  INV_X1    g405(.A(G233gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n582), .B2(KEYINPUT21), .ZN(new_n609));
  INV_X1    g408(.A(G127gat), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT21), .ZN(new_n611));
  INV_X1    g410(.A(new_n608), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n554), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n554), .B2(new_n611), .ZN(new_n615));
  AOI211_X1 g414(.A(KEYINPUT21), .B(new_n608), .C1(new_n551), .C2(new_n553), .ZN(new_n616));
  OAI21_X1  g415(.A(G127gat), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G183gat), .B(G211gat), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n614), .B2(new_n617), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT21), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n486), .A2(new_n489), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT94), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT94), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n486), .A2(new_n489), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(new_n305), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n625), .B2(new_n627), .ZN(new_n633));
  OAI22_X1  g432(.A1(new_n621), .A2(new_n622), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n617), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n618), .ZN(new_n636));
  INV_X1    g435(.A(new_n633), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n636), .A2(new_n620), .A3(new_n637), .A4(new_n631), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n577), .A2(new_n578), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n640), .B1(new_n528), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n581), .A2(new_n514), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(KEYINPUT96), .A3(new_n640), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n641), .B1(new_n515), .B2(new_n518), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n650), .B1(new_n647), .B2(new_n648), .ZN(new_n653));
  XNOR2_X1  g452(.A(G190gat), .B(G218gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G134gat), .B(G162gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n652), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT96), .B1(new_n645), .B2(new_n640), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n648), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n649), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n656), .B1(new_n662), .B2(new_n651), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n639), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT100), .B1(new_n605), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n634), .A2(new_n638), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n657), .B1(new_n652), .B2(new_n653), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n662), .A2(new_n651), .A3(new_n656), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n600), .A2(new_n602), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT99), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n669), .A2(new_n673), .A3(new_n674), .A4(new_n595), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n665), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n544), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n436), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(new_n480), .ZN(G1324gat));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  NAND4_X1  g479(.A1(new_n544), .A2(new_n365), .A3(new_n676), .A4(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G8gat), .B1(new_n677), .B2(new_n281), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n681), .ZN(new_n683));
  MUX2_X1   g482(.A(new_n681), .B(new_n683), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g483(.A(G15gat), .B1(new_n677), .B2(new_n475), .ZN(new_n685));
  INV_X1    g484(.A(new_n398), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n677), .B2(new_n687), .ZN(G1326gat));
  NAND3_X1  g487(.A1(new_n544), .A2(new_n430), .A3(new_n676), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT101), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NOR2_X1   g491(.A1(new_n658), .A2(new_n663), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(new_n605), .A3(new_n639), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n544), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n436), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n496), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n468), .A2(new_n470), .ZN(new_n702));
  INV_X1    g501(.A(new_n456), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n477), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n443), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n432), .A2(new_n440), .A3(KEYINPUT104), .A4(new_n442), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n701), .B1(new_n708), .B2(new_n694), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n478), .A2(KEYINPUT44), .A3(new_n693), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n605), .B(KEYINPUT103), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n543), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n639), .B(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n436), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n719), .ZN(G1328gat));
  OR2_X1    g519(.A1(new_n503), .A2(new_n504), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n696), .A2(new_n281), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n721), .B1(new_n718), .B2(new_n281), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1329gat));
  INV_X1    g525(.A(new_n475), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n709), .A2(new_n727), .A3(new_n710), .A4(new_n717), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G43gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n686), .A2(G43gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n697), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT47), .B1(new_n732), .B2(KEYINPUT106), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n728), .A2(G43gat), .B1(new_n697), .B2(new_n730), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n733), .A2(new_n737), .ZN(G1330gat));
  NAND4_X1  g537(.A1(new_n709), .A2(new_n430), .A3(new_n710), .A4(new_n717), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G50gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n429), .A2(G50gat), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n478), .A2(new_n543), .A3(new_n695), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT48), .B1(new_n742), .B2(KEYINPUT107), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT108), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n743), .B(new_n745), .ZN(G1331gat));
  NOR3_X1   g545(.A1(new_n712), .A2(new_n543), .A3(new_n664), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT109), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n708), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n698), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g550(.A1(new_n708), .A2(new_n281), .A3(new_n748), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  AND2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n752), .B2(new_n753), .ZN(G1333gat));
  INV_X1    g555(.A(G71gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n749), .A2(new_n757), .A3(new_n398), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n708), .A2(new_n475), .A3(new_n748), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n757), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g560(.A1(new_n749), .A2(new_n430), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n708), .A2(new_n694), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n543), .A2(new_n639), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT51), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  INV_X1    g566(.A(new_n765), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n708), .A2(new_n767), .A3(new_n694), .A4(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(new_n560), .A3(new_n698), .A4(new_n605), .ZN(new_n771));
  INV_X1    g570(.A(new_n605), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n711), .A2(new_n698), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n560), .B2(new_n774), .ZN(G1336gat));
  NOR2_X1   g574(.A1(new_n281), .A2(G92gat), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n713), .B(new_n776), .C1(new_n766), .C2(new_n769), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n709), .A2(new_n365), .A3(new_n710), .A4(new_n773), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G92gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1337gat));
  INV_X1    g584(.A(G99gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n770), .A2(new_n786), .A3(new_n398), .A4(new_n605), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n709), .A2(new_n727), .A3(new_n710), .A4(new_n773), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n786), .B1(new_n788), .B2(KEYINPUT111), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(KEYINPUT111), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1338gat));
  NAND4_X1  g590(.A1(new_n709), .A2(new_n430), .A3(new_n710), .A4(new_n773), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n792), .A2(G106gat), .B1(KEYINPUT112), .B2(KEYINPUT53), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n429), .A2(G106gat), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n713), .B(new_n794), .C1(new_n766), .C2(new_n769), .ZN(new_n795));
  OR2_X1    g594(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n793), .B2(new_n795), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(G1339gat));
  NOR3_X1   g598(.A1(new_n605), .A2(new_n664), .A3(new_n543), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n580), .A2(new_n598), .A3(new_n583), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n587), .A2(KEYINPUT54), .A3(new_n589), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n586), .A2(new_n597), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n584), .A2(KEYINPUT98), .A3(new_n585), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n802), .A2(new_n806), .A3(KEYINPUT55), .A4(new_n602), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(new_n595), .ZN(new_n808));
  INV_X1    g607(.A(new_n531), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n529), .A2(new_n521), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n810), .B(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n538), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n542), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n802), .A2(new_n602), .A3(new_n806), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n808), .A2(new_n693), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n541), .A2(new_n542), .B1(new_n816), .B2(new_n817), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n820), .A2(new_n808), .B1(new_n605), .B2(new_n815), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n821), .B2(new_n693), .ZN(new_n822));
  INV_X1    g621(.A(new_n716), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n800), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n436), .ZN(new_n825));
  INV_X1    g624(.A(new_n438), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n365), .ZN(new_n828));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n543), .ZN(new_n829));
  AND4_X1   g628(.A1(new_n543), .A2(new_n595), .A3(new_n818), .A4(new_n807), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n542), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n673), .B2(new_n595), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n694), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n716), .B1(new_n833), .B2(new_n819), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n429), .B1(new_n834), .B2(new_n800), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n365), .A2(new_n436), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n398), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT115), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n838), .A2(new_n842), .A3(new_n398), .A4(new_n839), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n543), .A2(G113gat), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n829), .B1(new_n844), .B2(new_n845), .ZN(G1340gat));
  INV_X1    g645(.A(G120gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n847), .A3(new_n605), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n841), .A2(new_n713), .A3(new_n843), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n849), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT116), .B1(new_n849), .B2(G120gat), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(G1341gat));
  XOR2_X1   g651(.A(KEYINPUT67), .B(G127gat), .Z(new_n853));
  NAND3_X1  g652(.A1(new_n828), .A2(new_n853), .A3(new_n639), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n844), .A2(new_n716), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n853), .ZN(G1342gat));
  NOR4_X1   g655(.A1(new_n827), .A2(G134gat), .A3(new_n365), .A4(new_n694), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT56), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n844), .A2(new_n693), .ZN(new_n859));
  INV_X1    g658(.A(G134gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(G1343gat));
  NAND2_X1  g660(.A1(new_n475), .A2(new_n839), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n824), .B2(new_n429), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n429), .A2(new_n864), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n820), .A2(new_n808), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n605), .A2(new_n815), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n693), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(KEYINPUT117), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n819), .B1(new_n870), .B2(KEYINPUT117), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n666), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n800), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n865), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI211_X1 g676(.A(KEYINPUT118), .B(new_n867), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n863), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n714), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n727), .A2(new_n429), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n825), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n365), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n301), .A3(new_n543), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT58), .ZN(G1344gat));
  OAI211_X1 g685(.A(new_n605), .B(new_n863), .C1(new_n877), .C2(new_n878), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n299), .A2(KEYINPUT59), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n822), .A2(new_n666), .B1(new_n676), .B2(new_n714), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n864), .B1(new_n890), .B2(new_n429), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT119), .B1(new_n824), .B2(new_n867), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n893), .B(new_n866), .C1(new_n834), .C2(new_n800), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n862), .A2(new_n772), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(KEYINPUT120), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G148gat), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT120), .B1(new_n895), .B2(new_n896), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT59), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g701(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n898), .C2(new_n899), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n889), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n883), .A2(new_n299), .A3(new_n605), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT122), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n888), .ZN(new_n908));
  INV_X1    g707(.A(new_n903), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n895), .A2(new_n896), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(G148gat), .A3(new_n897), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT121), .B1(new_n913), .B2(KEYINPUT59), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n908), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n905), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n907), .A2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(G155gat), .B1(new_n879), .B2(new_n823), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n883), .A2(new_n305), .A3(new_n639), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n879), .B2(new_n694), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n281), .A2(new_n306), .A3(new_n693), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n882), .B2(new_n923), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n824), .A2(new_n698), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n438), .A2(new_n281), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n543), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n698), .A2(new_n281), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n838), .A2(new_n398), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n714), .A2(new_n231), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1348gat));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n232), .A3(new_n605), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n931), .A2(new_n713), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(new_n232), .ZN(G1349gat));
  AOI21_X1  g735(.A(new_n237), .B1(new_n931), .B2(new_n716), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n928), .A2(new_n224), .A3(new_n639), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n940), .B(new_n941), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n928), .A2(new_n225), .A3(new_n693), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n931), .A2(new_n693), .ZN(new_n944));
  XNOR2_X1  g743(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n944), .A2(G190gat), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n944), .B2(G190gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1351gat));
  AND3_X1   g747(.A1(new_n881), .A2(new_n925), .A3(new_n365), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n543), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n475), .A2(new_n930), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n895), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n543), .A2(G197gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(G1352gat));
  XOR2_X1   g754(.A(KEYINPUT124), .B(G204gat), .Z(new_n956));
  NOR2_X1   g755(.A1(new_n772), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n949), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT62), .Z(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n952), .B2(new_n712), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT125), .Z(G1353gat));
  NAND3_X1  g761(.A1(new_n953), .A2(KEYINPUT126), .A3(new_n639), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n964), .B1(new_n952), .B2(new_n666), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n963), .A2(G211gat), .A3(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n967), .A3(KEYINPUT63), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n949), .A2(new_n205), .A3(new_n639), .ZN(new_n969));
  XOR2_X1   g768(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n970));
  OAI211_X1 g769(.A(new_n968), .B(new_n969), .C1(new_n966), .C2(new_n970), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n952), .B2(new_n694), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n949), .A2(new_n206), .A3(new_n693), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1355gat));
endmodule


