//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  XOR2_X1   g000(.A(KEYINPUT90), .B(G8gat), .Z(new_n202));
  INV_X1    g001(.A(G15gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G15gat), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n202), .B(new_n209), .C1(G1gat), .C2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT91), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n204), .A2(new_n206), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(new_n207), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G8gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n215), .A2(KEYINPUT91), .A3(new_n209), .A4(new_n202), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G50gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G43gat), .ZN(new_n222));
  INV_X1    g021(.A(G43gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G50gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT87), .ZN(new_n225));
  OR3_X1    g024(.A1(new_n223), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT88), .A4(new_n227), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT83), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n223), .A2(G50gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n221), .A2(G43gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT83), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(KEYINPUT15), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G29gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT86), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT86), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G29gat), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n240), .A2(new_n242), .A3(G36gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT84), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(KEYINPUT84), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(G29gat), .A2(G36gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT14), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n244), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT85), .ZN(new_n255));
  NOR4_X1   g054(.A1(new_n255), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT85), .B1(new_n250), .B2(new_n251), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n243), .B1(new_n258), .B2(new_n249), .ZN(new_n259));
  OAI22_X1  g058(.A1(new_n232), .A2(new_n254), .B1(new_n238), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT89), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT17), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n260), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n260), .B2(new_n261), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n220), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G229gat), .A2(G233gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT92), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n219), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n213), .A2(new_n217), .A3(new_n218), .A4(KEYINPUT92), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT83), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT83), .B1(new_n222), .B2(new_n224), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n243), .B1(new_n274), .B2(KEYINPUT15), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n275), .A2(new_n253), .A3(new_n230), .A4(new_n231), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n259), .A2(new_n238), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n270), .A2(new_n271), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n267), .A2(new_n268), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT93), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT18), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n276), .A2(new_n262), .A3(new_n277), .A4(new_n263), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n260), .A2(new_n261), .A3(new_n264), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n278), .B1(new_n286), .B2(new_n220), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(KEYINPUT93), .A3(new_n268), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n282), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n268), .B(KEYINPUT94), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT13), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n271), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(new_n260), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n293), .B2(new_n278), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n287), .A2(KEYINPUT18), .A3(new_n268), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n289), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G113gat), .B(G141gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(G197gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT11), .ZN(new_n299));
  INV_X1    g098(.A(G169gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n301), .B(KEYINPUT12), .Z(new_n302));
  AOI21_X1  g101(.A(KEYINPUT93), .B1(new_n287), .B2(new_n268), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n219), .B1(new_n284), .B2(new_n285), .ZN(new_n304));
  INV_X1    g103(.A(new_n268), .ZN(new_n305));
  NOR4_X1   g104(.A1(new_n304), .A2(new_n281), .A3(new_n305), .A4(new_n278), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n303), .A2(new_n306), .A3(KEYINPUT18), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n302), .B1(new_n307), .B2(KEYINPUT95), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n296), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n302), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT95), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(new_n289), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n289), .A2(new_n294), .A3(new_n295), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G71gat), .ZN(new_n317));
  INV_X1    g116(.A(G78gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT96), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT96), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(G71gat), .B2(G78gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G71gat), .A2(G78gat), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT97), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT97), .ZN(new_n325));
  AND2_X1   g124(.A1(G71gat), .A2(G78gat), .ZN(new_n326));
  AOI211_X1 g125(.A(new_n325), .B(new_n326), .C1(new_n319), .C2(new_n321), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(KEYINPUT9), .ZN(new_n328));
  XNOR2_X1  g127(.A(G57gat), .B(G64gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n324), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT98), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n317), .B(new_n318), .C1(new_n332), .C2(KEYINPUT9), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n323), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(KEYINPUT98), .B2(new_n328), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(new_n329), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G85gat), .A2(G92gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT100), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT100), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(G85gat), .A3(G92gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT7), .ZN(new_n342));
  NAND2_X1  g141(.A1(G99gat), .A2(G106gat), .ZN(new_n343));
  INV_X1    g142(.A(G85gat), .ZN(new_n344));
  INV_X1    g143(.A(G92gat), .ZN(new_n345));
  AOI22_X1  g144(.A1(KEYINPUT8), .A2(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT7), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n338), .A2(KEYINPUT100), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G99gat), .B(G106gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(KEYINPUT103), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n349), .A2(new_n351), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n342), .A2(new_n350), .A3(new_n346), .A4(new_n348), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT103), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n352), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n349), .A2(new_n351), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT101), .A3(new_n354), .ZN(new_n361));
  OR3_X1    g160(.A1(new_n349), .A2(KEYINPUT101), .A3(new_n351), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n361), .B(new_n362), .C1(new_n331), .C2(new_n336), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n362), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(new_n337), .A3(KEYINPUT10), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G230gat), .A2(G233gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n358), .A2(new_n363), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(G230gat), .A3(G233gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G120gat), .B(G148gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT104), .ZN(new_n373));
  INV_X1    g172(.A(G176gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G204gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n369), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n368), .B(KEYINPUT105), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n367), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n377), .B1(new_n381), .B2(new_n371), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n316), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G148gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(G141gat), .ZN(new_n388));
  INV_X1    g187(.A(G141gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(G148gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT72), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT2), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n391), .A2(new_n392), .B1(KEYINPUT73), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT72), .B1(new_n388), .B2(new_n390), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n394), .B(new_n395), .C1(KEYINPUT73), .C2(new_n393), .ZN(new_n396));
  XOR2_X1   g195(.A(G155gat), .B(G162gat), .Z(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n390), .A2(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n390), .A2(KEYINPUT74), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n399), .B(new_n400), .C1(G141gat), .C2(new_n387), .ZN(new_n401));
  INV_X1    g200(.A(G155gat), .ZN(new_n402));
  INV_X1    g201(.A(G162gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n393), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n402), .B2(new_n403), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n398), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT75), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n396), .A2(new_n397), .B1(new_n405), .B2(new_n401), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G127gat), .B(G134gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT64), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G113gat), .ZN(new_n416));
  INV_X1    g215(.A(G120gat), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT1), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n416), .B2(new_n417), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(KEYINPUT65), .B(G113gat), .Z(new_n421));
  OAI211_X1 g220(.A(new_n413), .B(new_n418), .C1(new_n421), .C2(new_n417), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n410), .A2(new_n411), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n408), .A2(new_n412), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT4), .B1(new_n407), .B2(new_n423), .ZN(new_n426));
  INV_X1    g225(.A(new_n423), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n433));
  AND2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n410), .B(new_n427), .ZN(new_n435));
  INV_X1    g234(.A(new_n431), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n433), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT0), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G57gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(new_n344), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT6), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n434), .B2(new_n438), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(KEYINPUT77), .B(new_n443), .C1(new_n434), .C2(new_n438), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT78), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT78), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n445), .A2(new_n448), .A3(new_n452), .A4(new_n449), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n444), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT27), .B(G183gat), .ZN(new_n457));
  INV_X1    g256(.A(G190gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n459), .A2(KEYINPUT28), .ZN(new_n460));
  NAND2_X1  g259(.A1(G183gat), .A2(G190gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(KEYINPUT28), .ZN(new_n462));
  NOR2_X1   g261(.A1(G169gat), .A2(G176gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT26), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n465), .B(new_n466), .C1(new_n300), .C2(new_n374), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n460), .A2(new_n461), .A3(new_n462), .A4(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT23), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n463), .B(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n461), .A2(KEYINPUT24), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n300), .A2(new_n374), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(G183gat), .A2(G190gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(KEYINPUT24), .A3(new_n461), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n470), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT25), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n476), .A2(new_n477), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n468), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n480), .A2(G226gat), .A3(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n480), .A2(new_n482), .B1(G226gat), .B2(G233gat), .ZN(new_n483));
  OR2_X1    g282(.A1(KEYINPUT69), .A2(KEYINPUT22), .ZN(new_n484));
  NAND2_X1  g283(.A1(KEYINPUT69), .A2(KEYINPUT22), .ZN(new_n485));
  INV_X1    g284(.A(G211gat), .ZN(new_n486));
  INV_X1    g285(.A(G218gat), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G197gat), .B(G204gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G211gat), .B(G218gat), .Z(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT70), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n490), .B(new_n492), .ZN(new_n493));
  OR3_X1    g292(.A1(new_n481), .A2(new_n483), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n481), .B2(new_n483), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G8gat), .B(G36gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT71), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(G64gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(G92gat), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT30), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n501), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n504), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n493), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(new_n424), .B2(new_n482), .ZN(new_n509));
  INV_X1    g308(.A(new_n491), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT29), .B1(new_n490), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n510), .B2(new_n490), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n410), .B1(new_n411), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G228gat), .ZN(new_n514));
  INV_X1    g313(.A(G233gat), .ZN(new_n515));
  OAI22_X1  g314(.A1(new_n509), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT79), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n508), .A2(new_n482), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n410), .B1(new_n518), .B2(new_n411), .ZN(new_n519));
  OR4_X1    g318(.A1(new_n514), .A2(new_n509), .A3(new_n515), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G22gat), .B(G78gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n521), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G50gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(G106gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n521), .B(new_n522), .ZN(new_n528));
  INV_X1    g327(.A(new_n526), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n480), .A2(new_n427), .ZN(new_n532));
  INV_X1    g331(.A(G227gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(new_n515), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n423), .B(new_n468), .C1(new_n478), .C2(new_n479), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G43gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G71gat), .ZN(new_n538));
  INV_X1    g337(.A(G99gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT33), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(KEYINPUT32), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT66), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n536), .A2(KEYINPUT66), .A3(KEYINPUT32), .A4(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT33), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n536), .B1(KEYINPUT32), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n540), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT34), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n535), .ZN(new_n552));
  INV_X1    g351(.A(new_n534), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI211_X1 g353(.A(KEYINPUT34), .B(new_n534), .C1(new_n532), .C2(new_n535), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n544), .A2(new_n545), .B1(new_n548), .B2(new_n540), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n556), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(KEYINPUT67), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT67), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n550), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n456), .A2(new_n507), .A3(new_n531), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT35), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n450), .A2(new_n455), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT35), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n558), .A2(new_n569), .A3(new_n560), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n559), .A2(KEYINPUT68), .A3(new_n556), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n531), .A2(new_n568), .A3(new_n507), .A4(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n566), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n527), .A2(new_n530), .A3(KEYINPUT80), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT80), .B1(new_n527), .B2(new_n530), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n456), .A2(new_n507), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(KEYINPUT81), .A2(KEYINPUT40), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n431), .B1(new_n425), .B2(new_n430), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n444), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n435), .A2(new_n436), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n585), .B2(new_n582), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n507), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n439), .A2(new_n444), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n587), .B(new_n588), .C1(new_n580), .C2(new_n586), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n496), .A2(KEYINPUT37), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n496), .A2(KEYINPUT37), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n503), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(KEYINPUT82), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(KEYINPUT38), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(KEYINPUT38), .B2(new_n593), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n504), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n567), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n589), .A2(new_n531), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n570), .A2(new_n571), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n561), .B2(new_n563), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n579), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n386), .B1(new_n574), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n486), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n337), .A2(KEYINPUT21), .ZN(new_n609));
  INV_X1    g408(.A(G127gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n292), .B1(KEYINPUT21), .B2(new_n337), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n616));
  XNOR2_X1  g415(.A(G155gat), .B(G183gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n615), .A2(new_n618), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n608), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(new_n607), .A3(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT99), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n629));
  XOR2_X1   g428(.A(G190gat), .B(G218gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n260), .A2(new_n365), .ZN(new_n633));
  INV_X1    g432(.A(new_n365), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n286), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT102), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n635), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n638), .B1(new_n635), .B2(new_n639), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n632), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n635), .A2(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n637), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(new_n631), .A3(new_n640), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n625), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n605), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n456), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n207), .ZN(G1324gat));
  INV_X1    g451(.A(new_n507), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n605), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(KEYINPUT106), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(KEYINPUT106), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(G8gat), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT16), .B(G8gat), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT42), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n661));
  OAI221_X1 g460(.A(new_n658), .B1(new_n654), .B2(new_n660), .C1(new_n661), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n570), .A2(new_n571), .A3(new_n599), .ZN(new_n664));
  INV_X1    g463(.A(new_n564), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n663), .B(new_n664), .C1(new_n665), .C2(new_n599), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT108), .B1(new_n600), .B2(new_n601), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n203), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT109), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n650), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n572), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n650), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(G15gat), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(KEYINPUT107), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(KEYINPUT107), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(G1326gat));
  INV_X1    g476(.A(new_n577), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT110), .B1(new_n650), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n605), .A2(new_n681), .A3(new_n649), .A4(new_n577), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n680), .B1(new_n679), .B2(new_n682), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n205), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(G22gat), .A3(new_n683), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n574), .A2(new_n604), .ZN(new_n690));
  INV_X1    g489(.A(new_n625), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n386), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n648), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n240), .A2(new_n242), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n693), .A2(new_n456), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n690), .A2(new_n697), .A3(new_n648), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n690), .B2(new_n648), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n692), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n694), .B1(new_n701), .B2(new_n456), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n696), .A2(new_n702), .ZN(G1328gat));
  NOR3_X1   g502(.A1(new_n693), .A2(G36gat), .A3(new_n507), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n701), .B2(new_n507), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  OAI21_X1  g506(.A(G43gat), .B1(new_n701), .B2(new_n603), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n693), .A2(G43gat), .A3(new_n672), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(KEYINPUT47), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n668), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n712), .B(new_n692), .C1(new_n699), .C2(new_n700), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n709), .B1(new_n713), .B2(G43gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n711), .B1(KEYINPUT47), .B2(new_n714), .ZN(G1330gat));
  OAI21_X1  g514(.A(G50gat), .B1(new_n701), .B2(new_n531), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n693), .A2(G50gat), .A3(new_n678), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(KEYINPUT48), .A3(new_n718), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n577), .B(new_n692), .C1(new_n699), .C2(new_n700), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n717), .B1(new_n720), .B2(G50gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(KEYINPUT48), .B2(new_n721), .ZN(G1331gat));
  AOI21_X1  g521(.A(new_n383), .B1(new_n574), .B2(new_n604), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n625), .A2(new_n315), .A3(new_n648), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n456), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT111), .B(G57gat), .Z(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1332gat));
  NOR2_X1   g527(.A1(new_n725), .A2(new_n507), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  OAI21_X1  g532(.A(G71gat), .B1(new_n725), .B2(new_n668), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n572), .A2(new_n317), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n725), .B2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g536(.A1(new_n725), .A2(new_n678), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n318), .ZN(G1335gat));
  NOR2_X1   g538(.A1(new_n691), .A2(new_n315), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n384), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT112), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n579), .A2(new_n598), .A3(new_n603), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n573), .A2(new_n567), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(KEYINPUT35), .B2(new_n565), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n648), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT44), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n743), .B1(new_n748), .B2(new_n698), .ZN(new_n749));
  INV_X1    g548(.A(new_n455), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n451), .B2(new_n453), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G85gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n690), .A2(new_n648), .A3(new_n740), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n690), .A2(KEYINPUT51), .A3(new_n648), .A4(new_n740), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT113), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n754), .B2(new_n755), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n751), .A2(new_n344), .A3(new_n384), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT114), .Z(new_n763));
  OAI21_X1  g562(.A(new_n753), .B1(new_n761), .B2(new_n763), .ZN(G1336gat));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n653), .B(new_n742), .C1(new_n699), .C2(new_n700), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(new_n345), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n507), .A2(G92gat), .A3(new_n383), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n758), .ZN(new_n771));
  INV_X1    g570(.A(new_n760), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n770), .B1(new_n756), .B2(new_n757), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(G92gat), .B2(new_n766), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n768), .A2(new_n773), .B1(new_n775), .B2(new_n765), .ZN(G1337gat));
  NAND2_X1  g575(.A1(new_n749), .A2(new_n712), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G99gat), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n539), .B(new_n572), .C1(new_n758), .C2(new_n760), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(new_n383), .ZN(G1338gat));
  INV_X1    g579(.A(G106gat), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n749), .B2(new_n577), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n531), .A2(G106gat), .A3(new_n383), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n756), .B2(new_n757), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT53), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n761), .B2(new_n784), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n527), .A2(new_n530), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n781), .B1(new_n749), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n786), .B1(new_n788), .B2(new_n790), .ZN(G1339gat));
  NOR4_X1   g590(.A1(new_n625), .A2(new_n315), .A3(new_n648), .A4(new_n384), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n369), .B(KEYINPUT54), .C1(new_n380), .C2(new_n367), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n367), .A2(new_n794), .A3(new_n380), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796));
  INV_X1    g595(.A(new_n377), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n796), .B1(new_n795), .B2(new_n797), .ZN(new_n799));
  OAI211_X1 g598(.A(KEYINPUT55), .B(new_n793), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n800), .A2(KEYINPUT116), .A3(new_n378), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT116), .B1(new_n800), .B2(new_n378), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n289), .A2(new_n310), .A3(new_n294), .A4(new_n295), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n287), .A2(new_n268), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n293), .A2(new_n278), .A3(new_n291), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n301), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n793), .B1(new_n798), .B2(new_n799), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n647), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n803), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n804), .A2(new_n384), .A3(new_n807), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n810), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n309), .B2(new_n314), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n815), .B1(new_n818), .B2(new_n803), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n813), .B1(new_n819), .B2(new_n648), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n792), .B1(new_n820), .B2(new_n625), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n751), .A2(new_n507), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n789), .A2(new_n665), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n421), .A3(new_n315), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n678), .A2(new_n572), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(new_n822), .A3(new_n821), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n315), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n830), .B2(new_n416), .ZN(G1340gat));
  NAND3_X1  g630(.A1(new_n826), .A2(new_n417), .A3(new_n384), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n829), .A2(new_n384), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n417), .ZN(G1341gat));
  AOI21_X1  g633(.A(G127gat), .B1(new_n826), .B2(new_n691), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n625), .A2(new_n610), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n829), .B2(new_n836), .ZN(G1342gat));
  NAND2_X1  g636(.A1(new_n823), .A2(new_n648), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(G134gat), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n824), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT56), .Z(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n838), .B2(new_n828), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1343gat));
  NOR2_X1   g642(.A1(new_n821), .A2(new_n531), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n751), .A3(new_n668), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n847), .A2(new_n507), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n316), .A2(G141gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n844), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n800), .A2(new_n378), .ZN(new_n855));
  AOI211_X1 g654(.A(new_n855), .B(new_n817), .C1(new_n309), .C2(new_n314), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n814), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n804), .A2(new_n384), .A3(KEYINPUT117), .A4(new_n807), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n647), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n813), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n792), .B1(new_n862), .B2(new_n625), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT57), .B1(new_n863), .B2(new_n678), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n822), .A2(new_n602), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n854), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G141gat), .B1(new_n866), .B2(new_n316), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n712), .A2(new_n531), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n823), .A2(new_n850), .A3(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n315), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n870), .B1(new_n874), .B2(G141gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n868), .B1(new_n875), .B2(new_n852), .ZN(G1344gat));
  AOI211_X1 g675(.A(KEYINPUT59), .B(new_n387), .C1(new_n873), .C2(new_n384), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT57), .B1(new_n821), .B2(new_n531), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT57), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n855), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n800), .A2(KEYINPUT116), .A3(new_n378), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n812), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT121), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n803), .A2(new_n886), .A3(new_n812), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n887), .A3(new_n809), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n691), .B1(new_n861), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n880), .B1(new_n889), .B2(new_n792), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n384), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n865), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n878), .B1(new_n893), .B2(G148gat), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n847), .A2(new_n387), .A3(new_n507), .A4(new_n848), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n383), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n895), .A2(new_n898), .A3(new_n383), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n877), .A2(new_n894), .B1(new_n897), .B2(new_n899), .ZN(G1345gat));
  NAND4_X1  g699(.A1(new_n847), .A2(new_n691), .A3(new_n507), .A4(new_n848), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n402), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n873), .A2(G155gat), .A3(new_n691), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  NAND3_X1  g705(.A1(new_n849), .A2(new_n403), .A3(new_n648), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n647), .B1(new_n871), .B2(new_n872), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n403), .ZN(G1347gat));
  INV_X1    g708(.A(new_n792), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n884), .A2(new_n808), .ZN(new_n911));
  INV_X1    g710(.A(new_n314), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n312), .A2(new_n313), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n816), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n882), .A2(new_n883), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n814), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n911), .B1(new_n916), .B2(new_n647), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n910), .B1(new_n917), .B2(new_n691), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n456), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n920), .A2(new_n653), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n824), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n300), .A3(new_n315), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n678), .A2(new_n653), .A3(new_n572), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G169gat), .B1(new_n926), .B2(new_n316), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(new_n927), .ZN(G1348gat));
  NOR3_X1   g727(.A1(new_n926), .A2(new_n374), .A3(new_n383), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n922), .A2(new_n384), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(new_n374), .ZN(G1349gat));
  OAI21_X1  g730(.A(G183gat), .B1(new_n926), .B2(new_n625), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n921), .A2(new_n457), .A3(new_n824), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n625), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT60), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n936), .B(new_n932), .C1(new_n933), .C2(new_n625), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n458), .A3(new_n648), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n458), .B1(new_n925), .B2(new_n648), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT61), .Z(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1351gat));
  AND3_X1   g741(.A1(new_n920), .A2(new_n653), .A3(new_n869), .ZN(new_n943));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(new_n315), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n668), .A2(new_n456), .A3(new_n653), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n668), .A2(new_n456), .A3(KEYINPUT124), .A4(new_n653), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n891), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n316), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n945), .A2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n943), .A2(new_n954), .A3(new_n376), .A4(new_n384), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n892), .A2(new_n950), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G204gat), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n920), .A2(new_n376), .A3(new_n653), .A4(new_n869), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT62), .B1(new_n958), .B2(new_n383), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT125), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n955), .A2(new_n957), .A3(new_n959), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1353gat));
  NAND3_X1  g763(.A1(new_n943), .A2(new_n486), .A3(new_n691), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n879), .A2(new_n691), .A3(new_n890), .A4(new_n950), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n891), .A2(new_n967), .A3(new_n691), .A4(new_n950), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n971));
  AND4_X1   g770(.A1(KEYINPUT63), .A2(new_n970), .A3(G211gat), .A4(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n965), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n975), .B(new_n965), .C1(new_n969), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(G1354gat));
  NOR3_X1   g776(.A1(new_n951), .A2(new_n487), .A3(new_n647), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n943), .A2(new_n648), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n979), .B2(new_n487), .ZN(G1355gat));
endmodule


