//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT74), .ZN(new_n194));
  XNOR2_X1  g008(.A(G110), .B(G140), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(new_n198), .B2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n199), .A2(new_n201), .A3(new_n204), .A4(new_n202), .ZN(new_n207));
  XOR2_X1   g021(.A(KEYINPUT0), .B(G128), .Z(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n200), .A2(G143), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n211));
  OAI21_X1  g025(.A(G146), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n198), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(KEYINPUT0), .A3(G128), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G104), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT3), .B1(new_n220), .B2(G107), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(G107), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G101), .ZN(new_n225));
  INV_X1    g039(.A(G101), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n226), .B(new_n219), .C1(new_n221), .C2(new_n222), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT4), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n217), .B1(new_n218), .B2(G104), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n218), .A2(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n226), .B1(new_n231), .B2(new_n219), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT75), .B(new_n225), .C1(new_n228), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n223), .A2(G101), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT75), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT4), .A4(new_n227), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n216), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n199), .A2(new_n201), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n213), .B1(new_n240), .B2(G146), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT64), .B(G143), .ZN(new_n242));
  OAI211_X1 g056(.A(G128), .B(new_n214), .C1(new_n242), .C2(new_n202), .ZN(new_n243));
  OAI22_X1  g057(.A1(new_n239), .A2(new_n241), .B1(new_n243), .B2(KEYINPUT1), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n218), .A2(G104), .ZN(new_n245));
  OAI21_X1  g059(.A(G101), .B1(new_n222), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n227), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT10), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n227), .A2(KEYINPUT10), .A3(new_n246), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g065(.A(G128), .B1(new_n213), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n206), .A2(new_n207), .A3(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n212), .A2(new_n251), .A3(G128), .A4(new_n214), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n237), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT11), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G137), .ZN(new_n259));
  INV_X1    g073(.A(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT11), .A3(G134), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G131), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(G131), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n259), .A2(new_n261), .A3(new_n266), .A4(new_n262), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n197), .B1(new_n256), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n239), .A2(new_n241), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n202), .B1(new_n199), .B2(new_n201), .ZN(new_n272));
  NOR4_X1   g086(.A1(new_n272), .A2(KEYINPUT1), .A3(new_n238), .A4(new_n213), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n248), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n255), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n233), .A2(new_n236), .ZN(new_n277));
  INV_X1    g091(.A(new_n216), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n276), .A2(new_n279), .A3(new_n197), .A4(new_n269), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n196), .B1(new_n270), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT81), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n253), .A2(new_n254), .A3(new_n247), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT78), .A4(new_n247), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT79), .A3(new_n274), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n286), .A2(new_n287), .B1(new_n248), .B2(new_n244), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n291));
  OR3_X1    g105(.A1(new_n291), .A2(KEYINPUT79), .A3(KEYINPUT12), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n288), .A2(new_n274), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n269), .A2(new_n291), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n293), .A2(new_n268), .B1(KEYINPUT12), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n196), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n276), .A2(new_n279), .A3(new_n269), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT76), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n298), .B1(new_n300), .B2(new_n280), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT81), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n283), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(new_n280), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n256), .A2(new_n269), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n298), .ZN(new_n308));
  AOI21_X1  g122(.A(G902), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n288), .A2(KEYINPUT79), .A3(new_n274), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n292), .B1(new_n288), .B2(new_n274), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n268), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n296), .A2(KEYINPUT12), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n305), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n314), .A2(new_n298), .B1(new_n306), .B2(new_n301), .ZN(new_n315));
  OAI21_X1  g129(.A(G469), .B1(new_n315), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n191), .A2(new_n309), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT80), .B(G469), .C1(new_n315), .C2(G902), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n190), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(G472), .A2(G902), .ZN(new_n321));
  INV_X1    g135(.A(new_n262), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n258), .A2(G137), .ZN(new_n323));
  OAI21_X1  g137(.A(G131), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n263), .B2(G131), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n253), .B2(new_n254), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n268), .A2(new_n215), .A3(new_n209), .ZN(new_n328));
  NAND2_X1  g142(.A1(KEYINPUT2), .A2(G113), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT67), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT67), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT2), .A3(G113), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OR2_X1    g147(.A1(KEYINPUT2), .A2(G113), .ZN(new_n334));
  XNOR2_X1  g148(.A(G116), .B(G119), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n334), .ZN(new_n337));
  INV_X1    g151(.A(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G116), .ZN(new_n339));
  INV_X1    g153(.A(G116), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G119), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n335), .A2(KEYINPUT68), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n336), .B1(new_n337), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n327), .A2(new_n328), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n347), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n268), .A2(new_n215), .A3(new_n209), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(new_n326), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT28), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT28), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G237), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(new_n192), .A3(G210), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(G101), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT69), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n353), .A2(new_n354), .A3(new_n356), .A4(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n327), .A2(KEYINPUT30), .A3(new_n328), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT30), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n350), .B2(new_n326), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n366), .A3(new_n349), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n348), .ZN(new_n368));
  INV_X1    g182(.A(new_n361), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n370), .A3(G472), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n355), .B1(new_n348), .B2(new_n351), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n348), .A2(new_n355), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n354), .B1(new_n374), .B2(new_n361), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n321), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT70), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n367), .A2(new_n361), .A3(new_n348), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT31), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT31), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n367), .A2(new_n380), .A3(new_n361), .A4(new_n348), .ZN(new_n381));
  INV_X1    g195(.A(new_n362), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n372), .B2(new_n373), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G472), .ZN(new_n385));
  INV_X1    g199(.A(G902), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT32), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n384), .A2(KEYINPUT32), .A3(new_n385), .A4(new_n386), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT70), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(new_n321), .C1(new_n371), .C2(new_n375), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n377), .A2(new_n389), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G217), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(G234), .B2(new_n386), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n338), .A2(G128), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n238), .A2(G119), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT24), .B(G110), .Z(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n397), .B1(KEYINPUT71), .B2(KEYINPUT23), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT71), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n338), .B2(G128), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G110), .ZN(new_n408));
  XNOR2_X1  g222(.A(G125), .B(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT16), .ZN(new_n410));
  INV_X1    g224(.A(G125), .ZN(new_n411));
  OR3_X1    g225(.A1(new_n411), .A2(KEYINPUT16), .A3(G140), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(G146), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n410), .A2(G146), .A3(new_n412), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n401), .B(new_n408), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n415), .ZN(new_n417));
  OAI22_X1  g231(.A1(new_n407), .A2(G110), .B1(new_n399), .B2(new_n400), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n409), .A2(new_n202), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT72), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT22), .B(G137), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n416), .A2(new_n420), .A3(new_n425), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n386), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT25), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n427), .A2(KEYINPUT25), .A3(new_n386), .A4(new_n428), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n396), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n427), .A2(new_n428), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n395), .A2(G902), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT73), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n393), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G478), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT93), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n340), .A2(G122), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n218), .B1(new_n450), .B2(KEYINPUT14), .ZN(new_n451));
  XNOR2_X1  g265(.A(G116), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n242), .A2(new_n238), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n198), .A2(G128), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT92), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT92), .ZN(new_n457));
  INV_X1    g271(.A(new_n455), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n457), .B(new_n458), .C1(new_n242), .C2(new_n238), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n258), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n258), .B1(new_n456), .B2(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n453), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT13), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n455), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n464), .B1(new_n454), .B2(new_n466), .ZN(new_n467));
  OAI221_X1 g281(.A(KEYINPUT90), .B1(new_n465), .B2(new_n455), .C1(new_n242), .C2(new_n238), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n454), .A2(KEYINPUT13), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT91), .A3(G134), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n452), .B(new_n218), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI22_X1  g287(.A1(KEYINPUT91), .A2(new_n460), .B1(new_n470), .B2(G134), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n188), .A2(new_n394), .A3(G953), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n476), .B(new_n463), .C1(new_n473), .C2(new_n474), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n449), .B1(new_n480), .B2(new_n386), .ZN(new_n481));
  AOI211_X1 g295(.A(G902), .B(new_n448), .C1(new_n478), .C2(new_n479), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G952), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n485), .A2(KEYINPUT94), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(KEYINPUT94), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n192), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(G234), .B2(G237), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT21), .B(G898), .Z(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n386), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G214), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n494), .A2(G237), .A3(G953), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G143), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n242), .B2(new_n495), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT87), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(G131), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n497), .B2(G131), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT17), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n242), .A2(new_n495), .ZN(new_n503));
  NOR4_X1   g317(.A1(new_n198), .A2(new_n494), .A3(G237), .A4(G953), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G131), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT87), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n497), .A2(G131), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n499), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n414), .A2(new_n415), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n502), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G113), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT89), .B(G104), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT86), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n409), .B(new_n202), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n517), .A2(new_n518), .B1(new_n505), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n497), .A2(KEYINPUT18), .A3(G131), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n409), .A2(new_n202), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n419), .A3(KEYINPUT86), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n508), .A4(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n512), .A2(new_n516), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n516), .B1(new_n512), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n386), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G475), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT20), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n507), .A2(new_n508), .A3(new_n499), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT88), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT19), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n409), .B(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n533), .B2(G146), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n409), .B(KEYINPUT19), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT88), .A3(new_n202), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n417), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n524), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n515), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n512), .A2(new_n516), .A3(new_n524), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(G475), .A2(G902), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n529), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n542), .ZN(new_n544));
  AOI211_X1 g358(.A(KEYINPUT20), .B(new_n544), .C1(new_n539), .C2(new_n540), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n528), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n484), .A2(new_n493), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G214), .B1(G237), .B2(G902), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT82), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n216), .A2(G125), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n253), .A2(new_n254), .A3(new_n411), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n550), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT85), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT83), .B(G224), .Z(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n192), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI22_X1  g373(.A1(new_n553), .A2(new_n555), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(KEYINPUT7), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT5), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT5), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n338), .A3(G116), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n566), .A2(G113), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(KEYINPUT84), .B(new_n247), .C1(new_n568), .C2(new_n336), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT84), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n336), .B1(new_n564), .B2(new_n567), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(new_n248), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n567), .B1(new_n565), .B2(new_n342), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n248), .B(new_n573), .C1(new_n337), .C2(new_n342), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(G110), .B(G122), .Z(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(KEYINPUT8), .Z(new_n577));
  AOI22_X1  g391(.A1(new_n277), .A2(new_n349), .B1(new_n248), .B2(new_n571), .ZN(new_n578));
  INV_X1    g392(.A(new_n576), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n575), .A2(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI221_X1 g394(.A(new_n561), .B1(new_n556), .B2(new_n559), .C1(new_n553), .C2(new_n555), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n563), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n559), .B1(new_n553), .B2(new_n555), .ZN(new_n583));
  INV_X1    g397(.A(new_n552), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n411), .B1(new_n209), .B2(new_n215), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT82), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n558), .A3(new_n554), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n277), .A2(new_n349), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n571), .A2(new_n248), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n579), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n347), .B1(new_n233), .B2(new_n236), .ZN(new_n592));
  AOI211_X1 g406(.A(new_n336), .B(new_n247), .C1(new_n564), .C2(new_n567), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n576), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n594), .A3(KEYINPUT6), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT6), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(new_n576), .C1(new_n592), .C2(new_n593), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n588), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n582), .A2(new_n598), .A3(new_n386), .ZN(new_n599));
  OAI21_X1  g413(.A(G210), .B1(G237), .B2(G902), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n582), .A2(new_n598), .A3(new_n386), .A4(new_n600), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n549), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n320), .A2(new_n442), .A3(new_n547), .A4(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT95), .B(G101), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G3));
  NAND2_X1  g421(.A1(new_n314), .A2(new_n298), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n301), .A2(new_n306), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n317), .B1(new_n610), .B2(new_n191), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n612));
  AOI211_X1 g426(.A(KEYINPUT81), .B(new_n298), .C1(new_n300), .C2(new_n280), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n308), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n191), .A3(new_n386), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n319), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n440), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n616), .A2(new_n189), .A3(new_n620), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n493), .B(new_n549), .C1(new_n602), .C2(new_n603), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n480), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n478), .A2(KEYINPUT33), .A3(new_n479), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n443), .A2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n480), .A2(new_n386), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n443), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n546), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n623), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n621), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NOR2_X1   g450(.A1(new_n483), .A2(new_n546), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n622), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n621), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NOR2_X1   g455(.A1(new_n426), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n421), .B(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n643), .A2(new_n437), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n433), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n618), .A2(new_n619), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(KEYINPUT96), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n618), .A2(new_n619), .A3(new_n645), .A4(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n320), .A2(new_n650), .A3(new_n547), .A4(new_n604), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n489), .B1(new_n654), .B2(new_n492), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n637), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n645), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n393), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n320), .A2(new_n604), .A3(new_n658), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XNOR2_X1  g477(.A(new_n655), .B(KEYINPUT39), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n320), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT40), .Z(new_n667));
  INV_X1    g481(.A(new_n378), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n352), .B2(new_n382), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n669), .B2(G902), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n389), .A2(new_n390), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT97), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n602), .A2(new_n603), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT38), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n541), .A2(new_n542), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT20), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n541), .A2(new_n529), .A3(new_n542), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n676), .A2(new_n677), .B1(G475), .B2(new_n527), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n483), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n548), .A3(new_n645), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT98), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n667), .A2(new_n672), .A3(new_n674), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n242), .ZN(G45));
  NOR2_X1   g497(.A1(new_n632), .A2(new_n655), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n320), .A2(new_n604), .A3(new_n661), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NAND2_X1  g500(.A1(new_n614), .A2(new_n386), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n688), .A2(new_n615), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n689), .A2(new_n189), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n690), .A2(new_n442), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n633), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n638), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NAND4_X1  g510(.A1(new_n688), .A2(new_n604), .A3(new_n189), .A4(new_n615), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n698), .A2(new_n393), .A3(new_n547), .A4(new_n659), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT99), .B(G119), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G21));
  XOR2_X1   g515(.A(new_n440), .B(KEYINPUT100), .Z(new_n702));
  NOR2_X1   g516(.A1(new_n618), .A2(new_n619), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n493), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n679), .A2(new_n705), .ZN(new_n706));
  OR3_X1    g520(.A1(new_n697), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT101), .B(G122), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G24));
  INV_X1    g523(.A(new_n646), .ZN(new_n710));
  INV_X1    g524(.A(new_n632), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n656), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n697), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n411), .ZN(G27));
  INV_X1    g528(.A(KEYINPUT42), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n389), .A2(new_n717), .A3(new_n390), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n717), .B1(new_n389), .B2(new_n390), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n377), .A2(new_n392), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n702), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n716), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n389), .A2(new_n390), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n389), .A2(new_n717), .A3(new_n390), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n377), .A3(new_n392), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT105), .A3(new_n702), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n615), .A2(new_n316), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n602), .A2(new_n731), .A3(new_n548), .A4(new_n603), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n602), .A2(new_n548), .A3(new_n603), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT102), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n730), .A2(new_n189), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT103), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n190), .B1(new_n615), .B2(new_n316), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT103), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n732), .A4(new_n734), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n712), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n715), .B1(new_n729), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n684), .A2(new_n715), .ZN(new_n742));
  AOI211_X1 g556(.A(new_n441), .B(new_n742), .C1(new_n736), .C2(new_n739), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  AOI211_X1 g559(.A(new_n441), .B(new_n657), .C1(new_n736), .C2(new_n739), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n258), .ZN(G36));
  AOI21_X1  g561(.A(new_n546), .B1(new_n630), .B2(new_n628), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT43), .Z(new_n749));
  OAI21_X1  g563(.A(new_n659), .B1(new_n618), .B2(new_n619), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n734), .A2(new_n732), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(new_n752), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n753), .A2(KEYINPUT107), .A3(new_n755), .A4(new_n756), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n315), .A2(KEYINPUT45), .ZN(new_n761));
  OAI21_X1  g575(.A(G469), .B1(new_n315), .B2(KEYINPUT45), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(G469), .A2(G902), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n615), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT46), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n189), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(new_n664), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n759), .A2(new_n760), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  XOR2_X1   g586(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n773));
  OR2_X1    g587(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n768), .B1(KEYINPUT108), .B2(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n754), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n778), .A2(new_n440), .A3(new_n393), .A4(new_n712), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  INV_X1    g595(.A(KEYINPUT48), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(KEYINPUT118), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n690), .A2(new_n489), .A3(new_n754), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(new_n749), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n783), .B(new_n785), .C1(new_n723), .C2(new_n728), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(KEYINPUT118), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n786), .B(new_n787), .Z(new_n788));
  NOR3_X1   g602(.A1(new_n784), .A2(new_n617), .A3(new_n672), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT116), .Z(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n711), .ZN(new_n791));
  INV_X1    g605(.A(new_n489), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n749), .A2(new_n792), .A3(new_n704), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(new_n690), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n488), .B1(new_n794), .B2(new_n604), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n788), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n631), .A2(new_n546), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n790), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n790), .A2(KEYINPUT117), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n674), .A2(new_n548), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n794), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT50), .ZN(new_n805));
  INV_X1    g619(.A(new_n785), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n805), .B1(new_n646), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n793), .A2(new_n755), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n689), .A2(new_n190), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n810), .B1(new_n776), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n796), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n712), .A2(new_n710), .ZN(new_n816));
  INV_X1    g630(.A(new_n739), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n738), .B1(new_n754), .B2(new_n737), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n678), .A2(new_n483), .A3(new_n656), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT112), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n678), .A2(new_n822), .A3(new_n483), .A4(new_n656), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n645), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n320), .A2(new_n393), .A3(new_n754), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n741), .A2(new_n826), .A3(new_n743), .A4(new_n746), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n698), .A2(new_n816), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n645), .A2(new_n656), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT113), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n679), .A2(new_n604), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n671), .A3(new_n831), .A4(new_n737), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n662), .A2(new_n685), .A3(new_n828), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n616), .A2(new_n604), .A3(new_n189), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n660), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n713), .B1(new_n836), .B2(new_n658), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n685), .A4(new_n832), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n690), .B(new_n442), .C1(new_n633), .C2(new_n638), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n699), .A3(new_n707), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT110), .B1(new_n622), .B2(new_n637), .ZN(new_n843));
  AND4_X1   g657(.A1(KEYINPUT110), .A2(new_n637), .A3(new_n604), .A4(new_n705), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n632), .A2(KEYINPUT109), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n632), .A2(KEYINPUT109), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n623), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n621), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n605), .A3(new_n651), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(new_n651), .A3(new_n605), .A4(KEYINPUT111), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n827), .A2(new_n840), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n833), .A2(new_n858), .A3(KEYINPUT52), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT52), .B1(new_n833), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n827), .A4(new_n854), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n855), .A2(new_n856), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n861), .A2(new_n854), .A3(new_n827), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(KEYINPUT53), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n867), .B2(KEYINPUT54), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n777), .A2(KEYINPUT115), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n776), .A2(new_n870), .B1(new_n190), .B2(new_n689), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n810), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n813), .B1(new_n808), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n815), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT49), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n689), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n689), .A2(new_n876), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n702), .A2(new_n548), .A3(new_n189), .A4(new_n748), .ZN(new_n879));
  OR4_X1    g693(.A1(new_n674), .A2(new_n877), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n874), .A2(new_n875), .B1(new_n672), .B2(new_n880), .ZN(G75));
  NOR2_X1   g695(.A1(new_n192), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n386), .B1(new_n857), .B2(new_n862), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT56), .B1(new_n884), .B2(G210), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n595), .A2(new_n597), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n588), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n883), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n863), .B2(G902), .ZN(new_n893));
  AOI211_X1 g707(.A(KEYINPUT119), .B(new_n386), .C1(new_n857), .C2(new_n862), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n600), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n891), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT120), .B1(new_n895), .B2(new_n600), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(G51));
  XOR2_X1   g714(.A(new_n863), .B(KEYINPUT54), .Z(new_n901));
  XNOR2_X1  g715(.A(new_n764), .B(KEYINPUT57), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n614), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n895), .A2(new_n763), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n882), .B1(new_n903), .B2(new_n904), .ZN(G54));
  AND2_X1   g719(.A1(KEYINPUT58), .A2(G475), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n893), .B2(new_n894), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n908));
  INV_X1    g722(.A(new_n541), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n883), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n541), .B(new_n906), .C1(new_n893), .C2(new_n894), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT121), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(G60));
  AND2_X1   g729(.A1(new_n625), .A2(new_n626), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT59), .Z(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n883), .B1(new_n901), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n924), .B(new_n883), .C1(new_n901), .C2(new_n921), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n917), .B1(new_n868), .B2(new_n919), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(G63));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT60), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n857), .B2(new_n862), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n643), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n931), .B(new_n883), .C1(new_n434), .C2(new_n930), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT124), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g748(.A(new_n557), .ZN(new_n935));
  OAI21_X1  g749(.A(G953), .B1(new_n491), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n854), .B2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n886), .B1(G898), .B2(new_n192), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  NAND3_X1  g753(.A1(new_n682), .A2(new_n685), .A3(new_n837), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  INV_X1    g755(.A(new_n780), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n846), .A2(new_n847), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n442), .B(new_n754), .C1(new_n944), .C2(new_n637), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(new_n666), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n771), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n192), .B1(new_n943), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n364), .A2(new_n366), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(new_n535), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n952), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n837), .A2(new_n685), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n729), .A2(new_n831), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n770), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n771), .A2(new_n780), .A3(new_n955), .A4(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  AOI21_X1  g776(.A(G953), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n192), .A2(G900), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT126), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n954), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n953), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n953), .B2(new_n966), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(G72));
  NAND3_X1  g784(.A1(new_n961), .A2(new_n854), .A3(new_n962), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n321), .B(KEYINPUT63), .Z(new_n972));
  AOI211_X1 g786(.A(new_n361), .B(new_n368), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n368), .A2(new_n361), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n947), .B(KEYINPUT125), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n941), .A2(new_n942), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(new_n976), .A3(new_n854), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n974), .B1(new_n977), .B2(new_n972), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n370), .A2(new_n378), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n867), .A2(new_n972), .A3(new_n979), .ZN(new_n980));
  NOR4_X1   g794(.A1(new_n973), .A2(new_n978), .A3(new_n980), .A4(new_n882), .ZN(G57));
endmodule


