//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT16), .A3(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT92), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n204), .B(new_n206), .C1(new_n203), .C2(new_n202), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n205), .A2(KEYINPUT92), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT14), .B(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n219), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n221), .A2(KEYINPUT90), .A3(new_n214), .A4(new_n216), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  OR3_X1    g023(.A1(new_n218), .A2(KEYINPUT91), .A3(KEYINPUT15), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT15), .B1(new_n218), .B2(KEYINPUT91), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n217), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n223), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n224), .B1(new_n223), .B2(new_n227), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n210), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(new_n227), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n209), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT18), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n232), .A4(new_n234), .ZN(new_n238));
  INV_X1    g037(.A(new_n233), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n210), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(KEYINPUT93), .A3(new_n234), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n232), .B(KEYINPUT13), .Z(new_n242));
  OR3_X1    g041(.A1(new_n233), .A2(new_n209), .A3(KEYINPUT93), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n237), .A2(new_n238), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(G169gat), .B(G197gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n245), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n244), .A4(new_n251), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G15gat), .B(G43gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G71gat), .B(G99gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G127gat), .B(G134gat), .Z(new_n260));
  INV_X1    g059(.A(G113gat), .ZN(new_n261));
  INV_X1    g060(.A(G120gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(G120gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n263), .B1(new_n261), .B2(new_n262), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n260), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n277), .A2(KEYINPUT26), .A3(new_n278), .ZN(new_n279));
  AOI211_X1 g078(.A(new_n274), .B(new_n279), .C1(KEYINPUT26), .C2(new_n278), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT27), .B(G183gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT67), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n282), .A2(new_n283), .A3(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT28), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n280), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n277), .B1(KEYINPUT23), .B2(new_n278), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n273), .A2(KEYINPUT24), .ZN(new_n291));
  XOR2_X1   g090(.A(G183gat), .B(G190gat), .Z(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(KEYINPUT24), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n278), .A2(KEYINPUT23), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT25), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(KEYINPUT65), .A3(new_n294), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n297), .A2(new_n298), .A3(new_n293), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n288), .A2(new_n294), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(KEYINPUT65), .B2(new_n300), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n287), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n272), .B1(new_n302), .B2(KEYINPUT69), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(KEYINPUT69), .B2(new_n302), .ZN(new_n304));
  NAND2_X1  g103(.A1(G227gat), .A2(G233gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT64), .ZN(new_n306));
  OR3_X1    g105(.A1(new_n302), .A2(KEYINPUT69), .A3(new_n271), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n259), .B1(new_n308), .B2(KEYINPUT32), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT33), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n308), .B2(new_n311), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT34), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n304), .A2(new_n307), .ZN(new_n316));
  INV_X1    g115(.A(new_n306), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI211_X1 g117(.A(KEYINPUT34), .B(new_n306), .C1(new_n304), .C2(new_n307), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n308), .B(KEYINPUT32), .C1(new_n311), .C2(new_n259), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n314), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n320), .B1(new_n314), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT72), .B(G218gat), .ZN(new_n326));
  INV_X1    g125(.A(G211gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n325), .B1(new_n328), .B2(KEYINPUT22), .ZN(new_n329));
  XNOR2_X1  g128(.A(G211gat), .B(G218gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G141gat), .B(G148gat), .Z(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT2), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G155gat), .B(G162gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n337), .B(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n333), .A2(new_n336), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n342), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT74), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n332), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n345), .A2(new_n348), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT3), .ZN(new_n354));
  AND2_X1   g153(.A1(G228gat), .A2(G233gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n350), .A3(new_n332), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n352), .A2(new_n354), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  OR3_X1    g156(.A1(new_n331), .A2(KEYINPUT83), .A3(KEYINPUT29), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT83), .B1(new_n331), .B2(KEYINPUT29), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n346), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n351), .B1(new_n360), .B2(new_n353), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n355), .B(KEYINPUT82), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n363), .A2(G22gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(G22gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT84), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n363), .B2(G22gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G78gat), .B(G106gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT81), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT31), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n371), .B(G50gat), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n366), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n364), .A2(new_n367), .A3(new_n365), .A4(new_n372), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT78), .ZN(new_n378));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G57gat), .B(G85gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n353), .A2(new_n271), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n343), .A2(new_n344), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(new_n272), .A3(new_n348), .A4(new_n338), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT75), .Z(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n392));
  INV_X1    g191(.A(new_n389), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n393), .B1(new_n384), .B2(new_n386), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT5), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n349), .A2(new_n271), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n389), .B1(new_n400), .B2(new_n354), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n391), .A2(new_n396), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n397), .A2(KEYINPUT79), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n354), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n397), .A2(KEYINPUT79), .A3(new_n398), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n389), .A2(KEYINPUT5), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n383), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n401), .A2(new_n399), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT76), .B1(new_n390), .B2(KEYINPUT5), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n394), .A2(new_n392), .A3(new_n395), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(new_n382), .A3(new_n407), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n409), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(KEYINPUT6), .B(new_n383), .C1(new_n402), .C2(new_n408), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n287), .A2(new_n301), .A3(new_n296), .ZN(new_n419));
  AND2_X1   g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n419), .B2(new_n350), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n332), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n331), .B1(new_n421), .B2(new_n422), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n424), .A2(new_n429), .A3(new_n425), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n433));
  OR3_X1    g232(.A1(new_n426), .A2(KEYINPUT30), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n418), .A2(KEYINPUT80), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT80), .B1(new_n418), .B2(new_n435), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n324), .B(new_n376), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT35), .ZN(new_n439));
  INV_X1    g238(.A(new_n376), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n435), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT88), .B(KEYINPUT35), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n322), .B2(new_n323), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n314), .A2(new_n321), .ZN(new_n446));
  INV_X1    g245(.A(new_n320), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n314), .A2(new_n320), .A3(new_n321), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT87), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n439), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n441), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n418), .A2(KEYINPUT80), .A3(new_n435), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n440), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT36), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n324), .B2(KEYINPUT71), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n389), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n382), .B1(new_n461), .B2(KEYINPUT39), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT39), .B1(new_n387), .B2(new_n389), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n460), .B2(new_n389), .ZN(new_n465));
  OR3_X1    g264(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n435), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n463), .B1(new_n462), .B2(new_n465), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n409), .A4(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n429), .B1(new_n424), .B2(new_n425), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n430), .A2(KEYINPUT37), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n426), .A2(KEYINPUT37), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n472), .B2(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n473), .A2(KEYINPUT85), .A3(new_n474), .A4(new_n476), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n432), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n469), .B(new_n376), .C1(new_n480), .C2(new_n418), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT71), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n482), .B(KEYINPUT36), .C1(new_n322), .C2(new_n323), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n457), .A2(new_n459), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n256), .B1(new_n453), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G71gat), .ZN(new_n486));
  INV_X1    g285(.A(G78gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G71gat), .A2(G78gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(KEYINPUT94), .A2(KEYINPUT9), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G57gat), .B(G64gat), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n488), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n495));
  INV_X1    g294(.A(new_n493), .ZN(new_n496));
  INV_X1    g295(.A(G57gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G64gat), .ZN(new_n498));
  INV_X1    g297(.A(G64gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G57gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT95), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n494), .A2(new_n502), .A3(KEYINPUT95), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(KEYINPUT21), .ZN(new_n508));
  NAND2_X1  g307(.A1(G231gat), .A2(G233gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(G127gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n209), .B1(new_n507), .B2(KEYINPUT21), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n511), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(new_n334), .ZN(new_n516));
  XNOR2_X1  g315(.A(G183gat), .B(G211gat), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n516), .B(new_n517), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n514), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(KEYINPUT96), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT96), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n523), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT8), .ZN(new_n526));
  OR2_X1    g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n522), .A2(new_n524), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n525), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT97), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n532), .A3(new_n525), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n528), .B2(new_n531), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n233), .A2(new_n538), .B1(KEYINPUT41), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n542));
  INV_X1    g341(.A(new_n230), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n228), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n542), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  AOI211_X1 g344(.A(KEYINPUT98), .B(new_n538), .C1(new_n543), .C2(new_n228), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n541), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT99), .Z(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n547), .A2(new_n550), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT100), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n547), .B2(new_n550), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT41), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G134gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n335), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI22_X1  g358(.A1(new_n552), .A2(new_n553), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n547), .A2(new_n550), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n561), .A2(new_n554), .A3(new_n551), .A4(new_n558), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n494), .A2(new_n502), .A3(KEYINPUT95), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT95), .B1(new_n494), .B2(new_n502), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n567), .A2(new_n537), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT102), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT101), .ZN(new_n572));
  INV_X1    g371(.A(new_n530), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n528), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n528), .B2(new_n572), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n503), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n567), .A2(new_n537), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n571), .B1(new_n577), .B2(new_n568), .ZN(new_n578));
  INV_X1    g377(.A(new_n536), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n505), .A2(new_n579), .A3(new_n534), .A4(new_n506), .ZN(new_n580));
  INV_X1    g379(.A(new_n575), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n581), .A2(new_n502), .A3(new_n494), .A4(new_n574), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n580), .A2(new_n571), .A3(new_n582), .A4(new_n568), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n570), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n577), .ZN(new_n588));
  INV_X1    g387(.A(new_n586), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n587), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n585), .A2(KEYINPUT103), .A3(new_n586), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n580), .A2(new_n568), .A3(new_n582), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT102), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n569), .B1(new_n601), .B2(new_n583), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n599), .B1(new_n602), .B2(new_n589), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n591), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n597), .B1(new_n604), .B2(new_n594), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n519), .A2(new_n564), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n485), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(new_n418), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(new_n203), .ZN(G1324gat));
  INV_X1    g408(.A(KEYINPUT104), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n485), .A2(new_n467), .A3(new_n606), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT16), .B(G8gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n613), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(KEYINPUT42), .B2(new_n613), .ZN(G1325gat));
  NAND2_X1  g414(.A1(new_n459), .A2(new_n483), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(G15gat), .B1(new_n607), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n451), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n619), .A2(G15gat), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n607), .B2(new_n620), .ZN(G1326gat));
  NOR2_X1   g420(.A1(new_n607), .A2(new_n376), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT43), .B(G22gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(G1327gat));
  AOI21_X1  g423(.A(new_n563), .B1(new_n453), .B2(new_n484), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n587), .A2(new_n596), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT103), .B1(new_n585), .B2(new_n586), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n602), .A2(new_n599), .A3(new_n589), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n590), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n629), .B2(new_n595), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n519), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n256), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n633), .A2(G29gat), .A3(new_n418), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  AND4_X1   g435(.A1(new_n457), .A2(new_n459), .A3(new_n481), .A4(new_n483), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n438), .A2(KEYINPUT35), .B1(new_n443), .B2(new_n451), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n564), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n453), .A2(new_n484), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(KEYINPUT44), .A3(new_n564), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n418), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n644), .A2(new_n645), .A3(new_n632), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n636), .B1(new_n215), .B2(new_n646), .ZN(G1328gat));
  NAND4_X1  g446(.A1(new_n641), .A2(new_n643), .A3(new_n467), .A4(new_n632), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n213), .B1(new_n648), .B2(KEYINPUT106), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(KEYINPUT106), .B2(new_n648), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n633), .A2(G36gat), .A3(new_n435), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT46), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(G1329gat));
  NAND3_X1  g452(.A1(new_n625), .A2(new_n451), .A3(new_n632), .ZN(new_n654));
  INV_X1    g453(.A(G43gat), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT107), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n654), .A2(new_n655), .B1(new_n656), .B2(KEYINPUT47), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n617), .A2(new_n655), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n641), .A2(new_n643), .A3(new_n632), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n656), .A2(KEYINPUT47), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT108), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(G1330gat));
  NAND4_X1  g462(.A1(new_n641), .A2(new_n643), .A3(new_n440), .A4(new_n632), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(G50gat), .ZN(new_n665));
  NOR4_X1   g464(.A1(new_n631), .A2(new_n376), .A3(G50gat), .A4(new_n563), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n485), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT48), .B1(new_n667), .B2(KEYINPUT109), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n665), .B(new_n667), .C1(KEYINPUT109), .C2(KEYINPUT48), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(G1331gat));
  NOR4_X1   g471(.A1(new_n519), .A2(new_n255), .A3(new_n564), .A4(new_n630), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n642), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n418), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT110), .B(G57gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1332gat));
  NOR2_X1   g476(.A1(new_n674), .A2(new_n435), .ZN(new_n678));
  NOR2_X1   g477(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n679));
  AND2_X1   g478(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n678), .B2(new_n679), .ZN(G1333gat));
  NAND4_X1  g481(.A1(new_n642), .A2(G71gat), .A3(new_n616), .A4(new_n673), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT111), .B1(new_n674), .B2(new_n619), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n486), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n674), .A2(KEYINPUT111), .A3(new_n619), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT50), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT50), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n689), .B(new_n683), .C1(new_n685), .C2(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1334gat));
  NOR2_X1   g490(.A1(new_n674), .A2(new_n376), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT112), .B(G78gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1335gat));
  INV_X1    g493(.A(new_n519), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n255), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n605), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n644), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G85gat), .B1(new_n699), .B2(new_n418), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n564), .B(new_n696), .C1(new_n637), .C2(new_n638), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT51), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n642), .A2(KEYINPUT51), .A3(new_n564), .A4(new_n696), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n630), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n418), .A2(G85gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n700), .B1(new_n706), .B2(new_n707), .ZN(G1336gat));
  NOR2_X1   g507(.A1(new_n435), .A2(G92gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n641), .A2(new_n643), .A3(new_n467), .A4(new_n698), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G92gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT52), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n710), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1337gat));
  OAI21_X1  g516(.A(G99gat), .B1(new_n699), .B2(new_n617), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n619), .A2(G99gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n706), .B2(new_n719), .ZN(G1338gat));
  INV_X1    g519(.A(KEYINPUT53), .ZN(new_n721));
  AOI21_X1  g520(.A(G106gat), .B1(new_n705), .B2(new_n440), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n440), .A2(G106gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  AND4_X1   g523(.A1(new_n641), .A2(new_n643), .A3(new_n698), .A4(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n721), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n725), .ZN(new_n727));
  AOI211_X1 g526(.A(new_n376), .B(new_n630), .C1(new_n703), .C2(new_n704), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n727), .B(KEYINPUT53), .C1(new_n728), .C2(G106gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(G1339gat));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT54), .B1(new_n602), .B2(new_n589), .ZN(new_n733));
  AOI211_X1 g532(.A(new_n586), .B(new_n569), .C1(new_n601), .C2(new_n583), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n602), .A2(new_n589), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n587), .A2(KEYINPUT113), .A3(KEYINPUT54), .A4(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n598), .A2(new_n603), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n595), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n731), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n735), .A2(new_n737), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n743), .A2(KEYINPUT55), .A3(new_n595), .A4(new_n740), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n742), .A2(new_n255), .A3(new_n597), .A4(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n242), .B1(new_n241), .B2(new_n243), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n232), .B1(new_n231), .B2(new_n234), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n250), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n254), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n605), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n564), .B1(new_n745), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n254), .A2(new_n748), .A3(KEYINPUT115), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n560), .A2(new_n562), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n744), .A2(new_n597), .ZN(new_n757));
  INV_X1    g556(.A(new_n741), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT55), .B1(new_n758), .B2(new_n743), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n519), .B1(new_n752), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n695), .A2(new_n256), .A3(new_n563), .A4(new_n630), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT116), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n761), .A2(new_n765), .A3(new_n762), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(new_n645), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n324), .A2(new_n376), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n467), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(G113gat), .B1(new_n772), .B2(new_n255), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n418), .A2(new_n467), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n767), .A2(new_n376), .A3(new_n451), .A4(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n256), .A2(new_n261), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n773), .B1(new_n779), .B2(new_n780), .ZN(G1340gat));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n605), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G120gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n772), .A2(new_n267), .A3(new_n605), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1341gat));
  NAND3_X1  g584(.A1(new_n777), .A2(new_n695), .A3(new_n778), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G127gat), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n519), .A2(G127gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n771), .B2(new_n788), .ZN(G1342gat));
  NAND3_X1  g588(.A1(new_n777), .A2(new_n564), .A3(new_n778), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G134gat), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792));
  AOI21_X1  g591(.A(G134gat), .B1(new_n792), .B2(KEYINPUT56), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n564), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n771), .A2(new_n795), .B1(new_n792), .B2(KEYINPUT56), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n792), .A2(KEYINPUT56), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n772), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n791), .A2(new_n796), .A3(new_n798), .ZN(G1343gat));
  NOR3_X1   g598(.A1(new_n616), .A2(new_n376), .A3(new_n467), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n767), .A2(new_n645), .A3(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n801), .A2(G141gat), .A3(new_n256), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(KEYINPUT58), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n459), .A2(new_n483), .A3(new_n774), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n630), .A2(new_n805), .A3(new_n749), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT119), .B1(new_n605), .B2(new_n750), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n564), .B1(new_n808), .B2(new_n745), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n519), .B1(new_n809), .B2(new_n760), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n762), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n440), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n804), .B1(new_n812), .B2(KEYINPUT57), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n764), .A2(new_n814), .A3(new_n440), .A4(new_n766), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G141gat), .B1(new_n816), .B2(new_n256), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n803), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(KEYINPUT120), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n813), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n255), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n802), .B1(new_n822), .B2(G141gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(G1344gat));
  NAND4_X1  g624(.A1(new_n764), .A2(KEYINPUT57), .A3(new_n440), .A4(new_n766), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827));
  NOR4_X1   g626(.A1(new_n519), .A2(new_n255), .A3(new_n564), .A4(new_n605), .ZN(new_n828));
  INV_X1    g627(.A(new_n760), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n805), .B1(new_n630), .B2(new_n749), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n605), .A2(new_n750), .A3(KEYINPUT119), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n757), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n759), .A2(new_n256), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n829), .B1(new_n835), .B2(new_n564), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n828), .B1(new_n836), .B2(new_n519), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n827), .B(new_n814), .C1(new_n837), .C2(new_n376), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n376), .B1(new_n810), .B2(new_n762), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT122), .B1(new_n839), .B2(KEYINPUT57), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n826), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n804), .A2(new_n630), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(G148gat), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n842), .B1(new_n841), .B2(new_n843), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT59), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(G148gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(KEYINPUT59), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n819), .A2(new_n821), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n630), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n801), .A2(G148gat), .A3(new_n630), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT121), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1345gat));
  OAI21_X1  g654(.A(G155gat), .B1(new_n850), .B2(new_n519), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n695), .A2(new_n334), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n801), .B2(new_n857), .ZN(G1346gat));
  OAI21_X1  g657(.A(G162gat), .B1(new_n850), .B2(new_n563), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n564), .A2(new_n335), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n801), .B2(new_n860), .ZN(G1347gat));
  NAND3_X1  g660(.A1(new_n451), .A2(new_n418), .A3(new_n467), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT125), .Z(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n376), .A3(new_n767), .ZN(new_n864));
  OAI21_X1  g663(.A(G169gat), .B1(new_n864), .B2(new_n256), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT126), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(KEYINPUT126), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n767), .A2(new_n418), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n769), .A2(new_n435), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n255), .A2(new_n275), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n870), .A2(KEYINPUT124), .A3(new_n871), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n866), .B(new_n867), .C1(new_n874), .C2(new_n875), .ZN(G1348gat));
  OAI21_X1  g675(.A(G176gat), .B1(new_n864), .B2(new_n630), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n605), .A2(new_n276), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n870), .B2(new_n878), .ZN(G1349gat));
  OAI21_X1  g678(.A(G183gat), .B1(new_n864), .B2(new_n519), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n519), .A2(new_n282), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n868), .A2(new_n869), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(KEYINPUT127), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT60), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n880), .A2(KEYINPUT127), .A3(new_n885), .A4(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n864), .B2(new_n563), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(KEYINPUT61), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n890), .B(G190gat), .C1(new_n864), .C2(new_n563), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n564), .A2(new_n285), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n889), .A2(new_n892), .B1(new_n870), .B2(new_n893), .ZN(G1351gat));
  NOR3_X1   g693(.A1(new_n616), .A2(new_n376), .A3(new_n435), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n868), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(G197gat), .B1(new_n896), .B2(new_n255), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n616), .A2(new_n645), .A3(new_n435), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n841), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n255), .A2(G197gat), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(G1352gat));
  NOR2_X1   g700(.A1(new_n630), .A2(G204gat), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT62), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n605), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G204gat), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n896), .A2(new_n907), .A3(new_n902), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n904), .A2(new_n906), .A3(new_n908), .ZN(G1353gat));
  NAND3_X1  g708(.A1(new_n896), .A2(new_n327), .A3(new_n695), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n841), .A2(new_n695), .A3(new_n898), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n911), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT63), .B1(new_n911), .B2(G211gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1354gat));
  AOI21_X1  g713(.A(G218gat), .B1(new_n896), .B2(new_n564), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n563), .A2(new_n326), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n899), .B2(new_n916), .ZN(G1355gat));
endmodule


