//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874;
  XNOR2_X1  g000(.A(G134gat), .B(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XOR2_X1   g002(.A(G43gat), .B(G50gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  AOI22_X1  g004(.A1(new_n204), .A2(new_n205), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT14), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n210), .C1(new_n205), .C2(new_n204), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT88), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n204), .A2(new_n205), .ZN(new_n214));
  OAI22_X1  g013(.A1(new_n210), .A2(KEYINPUT87), .B1(new_n207), .B2(new_n208), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n210), .A2(KEYINPUT87), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT17), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT98), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT7), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT99), .B(G85gat), .ZN(new_n223));
  INV_X1    g022(.A(G92gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n223), .A2(new_n224), .B1(KEYINPUT8), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(G99gat), .B(G106gat), .Z(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT100), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n227), .A2(new_n228), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n227), .A2(KEYINPUT100), .A3(new_n228), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n230), .B(new_n231), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n218), .ZN(new_n237));
  NAND3_X1  g036(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G190gat), .ZN(new_n240));
  INV_X1    g039(.A(G190gat), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n235), .A2(new_n237), .A3(new_n241), .A4(new_n238), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G218gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT96), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(G218gat), .A3(new_n242), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT94), .B(KEYINPUT95), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n249), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n245), .A2(new_n246), .A3(new_n253), .A4(new_n247), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n250), .B2(new_n254), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n203), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n250), .A2(new_n254), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n251), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n202), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G15gat), .B(G22gat), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n263), .A2(G1gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT16), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n265), .B2(G1gat), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G8gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT90), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n267), .B2(KEYINPUT89), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(KEYINPUT89), .B2(new_n264), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G57gat), .B(G64gat), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G71gat), .B(G78gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n273), .B1(KEYINPUT21), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G183gat), .ZN(new_n280));
  XOR2_X1   g079(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n278), .A2(KEYINPUT21), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT93), .B(G211gat), .Z(new_n285));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G127gat), .B(G155gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT92), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n287), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n284), .B(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n262), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G120gat), .B(G148gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(G176gat), .B(G204gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G230gat), .ZN(new_n296));
  INV_X1    g095(.A(G233gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n278), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n236), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n231), .A2(KEYINPUT101), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n229), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n227), .A2(KEYINPUT101), .A3(new_n228), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n278), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n234), .A2(new_n306), .A3(new_n299), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n298), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n305), .A2(new_n296), .A3(new_n297), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n295), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT10), .B1(new_n300), .B2(new_n304), .ZN(new_n314));
  OAI22_X1  g113(.A1(new_n314), .A2(new_n308), .B1(new_n296), .B2(new_n297), .ZN(new_n315));
  INV_X1    g114(.A(new_n295), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT102), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n312), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(KEYINPUT102), .B(new_n295), .C1(new_n310), .C2(new_n311), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n273), .A2(new_n218), .ZN(new_n322));
  INV_X1    g121(.A(new_n273), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n219), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G229gat), .A2(G233gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT18), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n273), .A2(new_n218), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n325), .B(KEYINPUT13), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n324), .A2(KEYINPUT18), .A3(new_n325), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G113gat), .B(G141gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(G197gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT11), .B(G169gat), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  XOR2_X1   g137(.A(new_n338), .B(KEYINPUT12), .Z(new_n339));
  NAND2_X1  g138(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n339), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n328), .A2(new_n332), .A3(new_n333), .A4(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n342), .A2(KEYINPUT91), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(KEYINPUT91), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n292), .A2(new_n321), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G197gat), .B(G204gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT22), .ZN(new_n348));
  NAND2_X1  g147(.A1(G211gat), .A2(G218gat), .ZN(new_n349));
  INV_X1    g148(.A(G211gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n244), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n350), .A2(new_n244), .A3(KEYINPUT22), .ZN(new_n355));
  INV_X1    g154(.A(new_n349), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n347), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G155gat), .B(G162gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G141gat), .B(G148gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(KEYINPUT2), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  INV_X1    g163(.A(G155gat), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT2), .B1(new_n365), .B2(KEYINPUT79), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n360), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n359), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n352), .B2(new_n357), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n368), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n370), .B1(new_n359), .B2(KEYINPUT29), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n379), .A2(new_n368), .B1(new_n359), .B2(new_n373), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n380), .B2(new_n375), .ZN(new_n381));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G22gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n381), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT31), .B(G50gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT65), .B(G169gat), .ZN(new_n389));
  INV_X1    g188(.A(G176gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT23), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n392), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  OAI22_X1  g193(.A1(new_n389), .A2(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT24), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n399));
  INV_X1    g198(.A(G183gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n241), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n388), .B1(new_n395), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT66), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n392), .A2(G176gat), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT65), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(G169gat), .ZN(new_n409));
  INV_X1    g208(.A(G169gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(KEYINPUT65), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n407), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT23), .B1(new_n410), .B2(new_n390), .ZN(new_n413));
  INV_X1    g212(.A(new_n394), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(new_n415), .A3(new_n402), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT66), .A3(new_n388), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n388), .B1(new_n407), .B2(new_n410), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n418), .A3(new_n402), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n406), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT26), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n394), .A2(KEYINPUT68), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n394), .B2(KEYINPUT68), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(new_n410), .B2(new_n390), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT67), .B1(new_n400), .B2(KEYINPUT27), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT27), .B(G183gat), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n241), .B(new_n426), .C1(new_n427), .C2(KEYINPUT67), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT28), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n427), .A2(KEYINPUT28), .A3(new_n241), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n396), .B(new_n425), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n420), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G127gat), .ZN(new_n434));
  INV_X1    g233(.A(G134gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G127gat), .A2(G134gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n436), .A2(KEYINPUT69), .A3(new_n437), .ZN(new_n441));
  XNOR2_X1  g240(.A(G113gat), .B(G120gat), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n440), .B(new_n441), .C1(KEYINPUT1), .C2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT71), .B(KEYINPUT1), .ZN(new_n444));
  INV_X1    g243(.A(new_n442), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n436), .A2(KEYINPUT70), .A3(new_n437), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT70), .B1(new_n436), .B2(new_n437), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n444), .B(new_n445), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n443), .A2(new_n448), .A3(KEYINPUT72), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT72), .B1(new_n443), .B2(new_n448), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n433), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G227gat), .A2(G233gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT34), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n454), .B(KEYINPUT64), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OR3_X1    g257(.A1(new_n452), .A2(KEYINPUT34), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G43gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n452), .A2(new_n458), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n461), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n387), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n416), .A2(KEYINPUT66), .A3(new_n388), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT66), .B1(new_n416), .B2(new_n388), .ZN(new_n478));
  INV_X1    g277(.A(new_n419), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n431), .B1(new_n429), .B2(new_n428), .ZN(new_n481));
  AOI211_X1 g280(.A(new_n423), .B(new_n422), .C1(G169gat), .C2(G176gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n396), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n372), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G226gat), .A2(G233gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT74), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n476), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT29), .B1(new_n420), .B2(new_n432), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n490), .A2(KEYINPUT75), .A3(new_n487), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT76), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n433), .A2(new_n487), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n358), .ZN(new_n495));
  INV_X1    g294(.A(new_n433), .ZN(new_n496));
  MUX2_X1   g295(.A(new_n490), .B(new_n496), .S(new_n487), .Z(new_n497));
  OR2_X1    g296(.A1(new_n497), .A2(new_n358), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n485), .A2(new_n476), .A3(new_n488), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT75), .B1(new_n490), .B2(new_n487), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n494), .A4(new_n358), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT76), .ZN(new_n502));
  XNOR2_X1  g301(.A(G8gat), .B(G36gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT77), .ZN(new_n504));
  XNOR2_X1  g303(.A(G64gat), .B(G92gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n504), .B(new_n505), .Z(new_n506));
  NAND4_X1  g305(.A1(new_n495), .A2(new_n498), .A3(new_n502), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT78), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT30), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n495), .A2(new_n498), .A3(new_n502), .ZN(new_n510));
  INV_X1    g309(.A(new_n506), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(KEYINPUT78), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n475), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G1gat), .B(G29gat), .Z(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(G85gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT0), .B(G57gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT4), .B(new_n369), .C1(new_n449), .C2(new_n450), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n443), .A2(new_n448), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n368), .A2(KEYINPUT3), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n371), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G225gat), .A2(G233gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT4), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n522), .B2(new_n368), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n521), .A2(new_n524), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n522), .B(new_n368), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n528), .B(KEYINPUT5), .C1(new_n525), .C2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n526), .B1(new_n451), .B2(new_n368), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n369), .A2(KEYINPUT4), .A3(new_n448), .A4(new_n443), .ZN(new_n533));
  INV_X1    g332(.A(new_n525), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT5), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n532), .A2(new_n524), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n520), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT6), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n537), .B(KEYINPUT81), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n531), .A2(new_n520), .A3(new_n536), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT35), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n516), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n537), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n539), .B1(new_n547), .B2(new_n543), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n515), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n387), .A3(new_n474), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n473), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(KEYINPUT36), .A3(new_n471), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n472), .B2(new_n473), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n549), .B2(new_n387), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT39), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n532), .A2(new_n524), .A3(new_n533), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT80), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n534), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n561), .B2(new_n534), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n566), .A2(new_n520), .ZN(new_n567));
  INV_X1    g366(.A(new_n565), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n560), .B1(new_n530), .B2(new_n525), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT40), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n566), .A2(new_n570), .A3(KEYINPUT40), .A4(new_n520), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n540), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n386), .B1(new_n574), .B2(new_n515), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n510), .A2(KEYINPUT37), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT85), .B1(new_n578), .B2(new_n511), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT85), .ZN(new_n580));
  AOI211_X1 g379(.A(new_n580), .B(new_n506), .C1(new_n510), .C2(KEYINPUT37), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT83), .B(KEYINPUT37), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n495), .A2(new_n498), .A3(new_n502), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n577), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT84), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n499), .A2(new_n500), .A3(new_n494), .A4(new_n359), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n588), .B(KEYINPUT37), .C1(new_n497), .C2(new_n359), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n585), .A2(new_n511), .A3(new_n577), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n537), .A2(KEYINPUT81), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT81), .ZN(new_n593));
  AOI211_X1 g392(.A(new_n593), .B(new_n520), .C1(new_n531), .C2(new_n536), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n543), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n538), .A3(new_n507), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n587), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n544), .A2(KEYINPUT84), .A3(new_n590), .A4(new_n507), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n575), .B1(new_n586), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT86), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n575), .B(KEYINPUT86), .C1(new_n586), .C2(new_n599), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n559), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n553), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n346), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n548), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n515), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT42), .B1(new_n610), .B2(new_n268), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G8gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  MUX2_X1   g413(.A(KEYINPUT42), .B(new_n611), .S(new_n614), .Z(G1325gat));
  AOI21_X1  g414(.A(G15gat), .B1(new_n606), .B2(new_n474), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT104), .ZN(new_n617));
  INV_X1    g416(.A(new_n558), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n618), .A2(G15gat), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n606), .B2(new_n619), .ZN(G1326gat));
  NAND2_X1  g419(.A1(new_n606), .A2(new_n386), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT105), .B(KEYINPUT106), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT43), .B(G22gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(G1327gat));
  OAI21_X1  g424(.A(new_n262), .B1(new_n553), .B2(new_n604), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n291), .ZN(new_n628));
  INV_X1    g427(.A(new_n321), .ZN(new_n629));
  INV_X1    g428(.A(new_n345), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n632), .A2(new_n207), .A3(new_n548), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT45), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n602), .A2(new_n603), .ZN(new_n635));
  INV_X1    g434(.A(new_n559), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT107), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n638));
  AOI211_X1 g437(.A(new_n638), .B(new_n559), .C1(new_n602), .C2(new_n603), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n552), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n262), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT108), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(new_n626), .B2(KEYINPUT44), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n640), .A2(new_n643), .A3(new_n641), .A4(new_n262), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n647), .A2(new_n548), .A3(new_n631), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n634), .B1(new_n648), .B2(new_n207), .ZN(G1328gat));
  NAND4_X1  g448(.A1(new_n645), .A2(new_n515), .A3(new_n646), .A4(new_n631), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT110), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(G36gat), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n632), .A2(new_n208), .A3(new_n515), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT109), .B(KEYINPUT46), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT111), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(KEYINPUT111), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(G1329gat));
  NAND4_X1  g461(.A1(new_n647), .A2(G43gat), .A3(new_n618), .A4(new_n631), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n632), .A2(new_n474), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n663), .B1(G43gat), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g465(.A1(new_n645), .A2(new_n386), .A3(new_n646), .A4(new_n631), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G50gat), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n387), .A2(G50gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT113), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n632), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(KEYINPUT48), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT48), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT112), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n667), .A2(new_n674), .A3(G50gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n674), .B1(new_n667), .B2(G50gat), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT114), .B(new_n673), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n668), .A2(KEYINPUT112), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n671), .A3(new_n675), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT114), .B1(new_n681), .B2(new_n673), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n672), .B1(new_n679), .B2(new_n682), .ZN(G1331gat));
  NOR2_X1   g482(.A1(new_n345), .A2(new_n321), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n640), .A2(new_n292), .A3(new_n684), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n685), .A2(KEYINPUT115), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(KEYINPUT115), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n548), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G57gat), .ZN(G1332gat));
  INV_X1    g490(.A(new_n515), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n694));
  AND2_X1   g493(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n693), .B2(new_n694), .ZN(G1333gat));
  INV_X1    g496(.A(new_n474), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n688), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n618), .A2(G71gat), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n699), .A2(G71gat), .B1(new_n688), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g501(.A1(new_n689), .A2(new_n386), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g503(.A1(new_n647), .A2(new_n291), .A3(new_n684), .ZN(new_n705));
  INV_X1    g504(.A(new_n548), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n705), .A2(new_n706), .A3(new_n223), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n640), .A2(new_n291), .A3(new_n262), .A4(new_n630), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT51), .Z(new_n709));
  AND2_X1   g508(.A1(new_n709), .A2(new_n629), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n548), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n707), .B1(new_n711), .B2(new_n223), .ZN(G1336gat));
  OAI21_X1  g511(.A(G92gat), .B1(new_n705), .B2(new_n692), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n709), .A2(new_n224), .A3(new_n515), .A4(new_n629), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g515(.A(G99gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n710), .A2(new_n717), .A3(new_n474), .ZN(new_n718));
  OAI21_X1  g517(.A(G99gat), .B1(new_n705), .B2(new_n558), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(G1338gat));
  OAI21_X1  g519(.A(G106gat), .B1(new_n705), .B2(new_n387), .ZN(new_n721));
  INV_X1    g520(.A(G106gat), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n709), .A2(new_n722), .A3(new_n386), .A4(new_n629), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g524(.A1(new_n292), .A2(new_n321), .A3(new_n630), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n307), .A2(new_n298), .A3(new_n309), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n315), .A3(KEYINPUT54), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT54), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n310), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n730), .A3(new_n295), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n728), .A2(new_n730), .A3(KEYINPUT55), .A4(new_n295), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n345), .A2(new_n317), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n338), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n330), .A2(new_n331), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT116), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n324), .A2(new_n325), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n343), .B2(new_n344), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n735), .B1(new_n321), .B2(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n743), .A2(new_n257), .A3(new_n261), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n733), .A2(new_n734), .A3(new_n317), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n742), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n257), .B2(new_n261), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n291), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n706), .B1(new_n726), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n516), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n630), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g552(.A1(new_n751), .A2(new_n321), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g554(.A1(new_n751), .A2(new_n291), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(new_n434), .ZN(G1342gat));
  INV_X1    g556(.A(new_n262), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n435), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT117), .Z(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n435), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT56), .Z(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1343gat));
  NAND2_X1  g563(.A1(new_n262), .A2(new_n746), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n342), .A2(KEYINPUT91), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n342), .A2(KEYINPUT91), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n740), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n629), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT118), .B1(new_n742), .B2(new_n321), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n735), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n257), .A3(new_n261), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n628), .B1(new_n765), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(KEYINPUT119), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n772), .A2(new_n261), .A3(new_n257), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT119), .B(new_n291), .C1(new_n776), .C2(new_n748), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n726), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n386), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT57), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n387), .B1(new_n726), .B2(new_n749), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n618), .A2(new_n706), .A3(new_n515), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n780), .A2(new_n345), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(KEYINPUT121), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(KEYINPUT121), .ZN(new_n787));
  INV_X1    g586(.A(G141gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n750), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n515), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n387), .B(new_n618), .C1(new_n750), .C2(new_n790), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n788), .A4(new_n345), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n785), .A2(G141gat), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n794), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n789), .A2(new_n796), .B1(new_n795), .B2(new_n798), .ZN(G1344gat));
  NAND3_X1  g598(.A1(new_n792), .A2(new_n793), .A3(new_n629), .ZN(new_n800));
  INV_X1    g599(.A(G148gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(KEYINPUT59), .A3(new_n801), .ZN(new_n802));
  NOR4_X1   g601(.A1(new_n262), .A2(new_n291), .A3(new_n629), .A4(new_n345), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n782), .B(new_n386), .C1(new_n774), .C2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n804), .B(new_n629), .C1(new_n781), .C2(new_n782), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n784), .A2(KEYINPUT59), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n780), .A2(new_n629), .A3(new_n783), .A4(new_n784), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n802), .B1(new_n810), .B2(new_n801), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT122), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n802), .B(new_n813), .C1(new_n810), .C2(new_n801), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1345gat));
  NAND4_X1  g614(.A1(new_n780), .A2(new_n628), .A3(new_n783), .A4(new_n784), .ZN(new_n816));
  XOR2_X1   g615(.A(KEYINPUT79), .B(G155gat), .Z(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n792), .A2(new_n793), .A3(new_n628), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n820), .B(new_n821), .ZN(G1346gat));
  AND3_X1   g621(.A1(new_n792), .A2(new_n793), .A3(new_n262), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n780), .A2(new_n784), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n262), .A3(new_n783), .ZN(new_n825));
  MUX2_X1   g624(.A(new_n823), .B(new_n825), .S(G162gat), .Z(G1347gat));
  NAND2_X1  g625(.A1(new_n515), .A2(new_n706), .ZN(new_n827));
  AOI211_X1 g626(.A(new_n475), .B(new_n827), .C1(new_n726), .C2(new_n749), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n345), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n389), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT124), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(G169gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1348gat));
  NAND2_X1  g632(.A1(new_n828), .A2(new_n629), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n390), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT126), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(KEYINPUT126), .ZN(new_n837));
  AOI21_X1  g636(.A(G176gat), .B1(new_n828), .B2(new_n629), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT125), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n838), .A2(KEYINPUT125), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n836), .A2(new_n837), .B1(new_n839), .B2(new_n840), .ZN(G1349gat));
  AND3_X1   g640(.A1(new_n828), .A2(new_n427), .A3(new_n628), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT127), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n628), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT127), .B1(new_n845), .B2(G183gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n846), .B2(new_n842), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g647(.A1(new_n828), .A2(new_n262), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n849), .A2(new_n850), .A3(new_n241), .ZN(new_n851));
  XOR2_X1   g650(.A(KEYINPUT61), .B(G190gat), .Z(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n849), .B2(new_n852), .ZN(G1351gat));
  NOR2_X1   g652(.A1(new_n618), .A2(new_n827), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n804), .B(new_n854), .C1(new_n781), .C2(new_n782), .ZN(new_n855));
  OAI21_X1  g654(.A(G197gat), .B1(new_n855), .B2(new_n630), .ZN(new_n856));
  INV_X1    g655(.A(new_n781), .ZN(new_n857));
  INV_X1    g656(.A(new_n854), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(G197gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n345), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n856), .A2(new_n861), .ZN(G1352gat));
  NOR4_X1   g661(.A1(new_n857), .A2(G204gat), .A3(new_n321), .A4(new_n858), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT62), .ZN(new_n864));
  OAI21_X1  g663(.A(G204gat), .B1(new_n805), .B2(new_n858), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1353gat));
  NAND3_X1  g665(.A1(new_n859), .A2(new_n350), .A3(new_n628), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n855), .A2(new_n291), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT63), .B1(new_n868), .B2(G211gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(G1354gat));
  OAI21_X1  g671(.A(G218gat), .B1(new_n855), .B2(new_n758), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n859), .A2(new_n244), .A3(new_n262), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1355gat));
endmodule


