//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n531, new_n532, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157, new_n1158;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT66), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT68), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  NAND2_X1  g031(.A1(G113), .A2(G2104), .ZN(new_n457));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(new_n460), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  AND2_X1   g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n460), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n460), .A2(new_n466), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  OAI21_X1  g055(.A(G2104), .B1(new_n466), .B2(G114), .ZN(new_n481));
  INV_X1    g056(.A(G102), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(new_n466), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(G126), .B2(new_n475), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n473), .A2(G138), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G164));
  INV_X1    g064(.A(G651), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT6), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G651), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n491), .A2(new_n493), .A3(G543), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G50), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n491), .A2(new_n493), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g077(.A(KEYINPUT71), .B(G88), .Z(new_n503));
  OAI21_X1  g078(.A(new_n495), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(new_n490), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n504), .A2(new_n506), .ZN(G166));
  NAND3_X1  g082(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n494), .A2(G51), .ZN(new_n509));
  NAND3_X1  g084(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT7), .ZN(new_n511));
  INV_X1    g086(.A(G89), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n502), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n508), .B(new_n509), .C1(new_n513), .C2(KEYINPUT72), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n513), .A2(KEYINPUT72), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(G168));
  NAND2_X1  g091(.A1(new_n494), .A2(G52), .ZN(new_n517));
  INV_X1    g092(.A(G90), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n502), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n490), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(G171));
  NAND2_X1  g097(.A1(new_n494), .A2(G43), .ZN(new_n523));
  INV_X1    g098(.A(G81), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n502), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n490), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G860), .ZN(G153));
  NAND4_X1  g104(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g105(.A1(G1), .A2(G3), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT8), .ZN(new_n532));
  NAND4_X1  g107(.A1(G319), .A2(G483), .A3(G661), .A4(new_n532), .ZN(G188));
  AND2_X1   g108(.A1(KEYINPUT5), .A2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(KEYINPUT73), .B1(new_n499), .B2(new_n500), .ZN(new_n538));
  OAI21_X1  g113(.A(G65), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(G78), .A2(G543), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(KEYINPUT74), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  INV_X1    g117(.A(G65), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n536), .B1(new_n534), .B2(new_n535), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n500), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n540), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n541), .A2(new_n548), .A3(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n494), .A2(G53), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n494), .A2(new_n552), .A3(G53), .ZN(new_n553));
  INV_X1    g128(.A(new_n502), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n551), .A2(new_n553), .B1(new_n554), .B2(G91), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT75), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n549), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  INV_X1    g136(.A(G168), .ZN(G286));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND3_X1  g138(.A1(new_n496), .A2(G49), .A3(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT76), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n501), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n554), .A2(G87), .B1(new_n566), .B2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n554), .A2(G86), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(KEYINPUT77), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n501), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(new_n494), .B2(G48), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n569), .A2(KEYINPUT77), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n570), .A2(new_n575), .A3(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(G72), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G60), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n572), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n490), .B1(new_n580), .B2(KEYINPUT78), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n581), .B1(KEYINPUT78), .B2(new_n580), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n494), .A2(G47), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n502), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n502), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n496), .A2(KEYINPUT10), .A3(G92), .A4(new_n501), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n591), .A2(new_n592), .B1(G54), .B2(new_n494), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n544), .B2(new_n545), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT79), .Z(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT80), .Z(new_n604));
  AND3_X1   g179(.A1(new_n549), .A2(new_n558), .A3(new_n555), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n558), .B1(new_n549), .B2(new_n555), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n604), .B1(G868), .B2(new_n607), .ZN(G297));
  OAI21_X1  g183(.A(new_n604), .B1(G868), .B2(new_n607), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n600), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n600), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n528), .ZN(G323));
  XOR2_X1   g189(.A(G323), .B(KEYINPUT81), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n473), .A2(G2104), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT82), .B(G2100), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT83), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n473), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n475), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  OAI211_X1 g203(.A(new_n622), .B(new_n628), .C1(new_n619), .C2(new_n620), .ZN(G156));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT14), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n635), .A2(new_n642), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n643), .A2(new_n644), .A3(G14), .ZN(G401));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT17), .Z(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  INV_X1    g226(.A(new_n648), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(new_n646), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n650), .B(new_n651), .C1(new_n649), .C2(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n646), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT84), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  OR2_X1    g245(.A1(new_n663), .A2(new_n665), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n666), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n672), .A2(KEYINPUT86), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(KEYINPUT86), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(new_n668), .ZN(new_n675));
  OAI221_X1 g250(.A(new_n670), .B1(new_n671), .B2(new_n668), .C1(new_n673), .C2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G23), .ZN(new_n686));
  INV_X1    g261(.A(G288), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n685), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT33), .Z(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(G1976), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(G1976), .ZN(new_n691));
  MUX2_X1   g266(.A(G6), .B(G305), .S(G16), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT88), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n685), .A2(G22), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT89), .Z(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n685), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT90), .B(G1971), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n690), .A2(new_n691), .A3(new_n695), .A4(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n703));
  AND3_X1   g278(.A1(new_n685), .A2(KEYINPUT87), .A3(G24), .ZN(new_n704));
  AOI21_X1  g279(.A(KEYINPUT87), .B1(new_n685), .B2(G24), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n704), .B(new_n705), .C1(G290), .C2(G16), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(new_n677), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n677), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G25), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n473), .A2(G131), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n475), .A2(G119), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n710), .B1(new_n716), .B2(new_n709), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  XOR2_X1   g293(.A(new_n717), .B(new_n718), .Z(new_n719));
  NOR3_X1   g294(.A1(new_n707), .A2(new_n708), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n702), .A2(new_n703), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT36), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n685), .A2(G20), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT23), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n607), .B2(new_n685), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1956), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT92), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT25), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n473), .A2(G139), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n729), .B(new_n730), .C1(new_n466), .C2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G33), .B(new_n732), .S(G29), .Z(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G2072), .Z(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  NOR2_X1   g310(.A1(G164), .A2(new_n709), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G27), .B2(new_n709), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n735), .ZN(new_n739));
  INV_X1    g314(.A(G28), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n740), .B2(KEYINPUT30), .ZN(new_n742));
  OR2_X1    g317(.A1(KEYINPUT31), .A2(G11), .ZN(new_n743));
  NAND2_X1  g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n627), .B2(new_n709), .ZN(new_n746));
  NOR2_X1   g321(.A1(G171), .A2(new_n685), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G5), .B2(new_n685), .ZN(new_n748));
  INV_X1    g323(.A(G1961), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n709), .A2(G32), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n475), .A2(G129), .ZN(new_n752));
  NAND2_X1  g327(.A1(G105), .A2(G2104), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT94), .B1(new_n753), .B2(G2105), .ZN(new_n754));
  OR3_X1    g329(.A1(new_n753), .A2(KEYINPUT94), .A3(G2105), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n473), .A2(G141), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT26), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n751), .B1(new_n761), .B2(new_n709), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT27), .B(G1996), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n473), .A2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n475), .A2(G128), .ZN(new_n766));
  NOR2_X1   g341(.A1(G104), .A2(G2105), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G29), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n709), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT91), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT28), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G2067), .Z(new_n775));
  NAND4_X1  g350(.A1(new_n739), .A2(new_n750), .A3(new_n764), .A4(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT24), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n709), .B1(new_n777), .B2(G34), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(KEYINPUT93), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(KEYINPUT93), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n777), .B2(G34), .ZN(new_n781));
  AOI22_X1  g356(.A1(G160), .A2(G29), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2084), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n738), .A2(new_n776), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n600), .A2(new_n685), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G4), .B2(new_n685), .ZN(new_n786));
  INV_X1    g361(.A(G1348), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n709), .A2(G35), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G162), .B2(new_n709), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT29), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n791), .A2(G2090), .B1(new_n786), .B2(new_n787), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n685), .A2(G19), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n528), .B2(new_n685), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1341), .Z(new_n795));
  OAI221_X1 g370(.A(new_n795), .B1(new_n749), .B2(new_n748), .C1(new_n791), .C2(G2090), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n685), .A2(G21), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G168), .B2(new_n685), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1966), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n784), .A2(new_n788), .A3(new_n792), .A4(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n722), .A2(new_n726), .A3(new_n801), .ZN(G311));
  INV_X1    g377(.A(G311), .ZN(G150));
  NAND2_X1  g378(.A1(new_n494), .A2(G55), .ZN(new_n804));
  INV_X1    g379(.A(G93), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n502), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n490), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n528), .A2(new_n809), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n527), .A2(new_n525), .B1(new_n806), .B2(new_n808), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT38), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n600), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  INV_X1    g391(.A(G860), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n809), .A2(new_n817), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT96), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n819), .A2(new_n823), .ZN(G145));
  XNOR2_X1  g399(.A(new_n715), .B(KEYINPUT97), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n618), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n473), .A2(G142), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n475), .A2(G130), .ZN(new_n828));
  NOR2_X1   g403(.A1(G106), .A2(G2105), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n826), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n488), .B(new_n769), .ZN(new_n833));
  INV_X1    g408(.A(new_n761), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(new_n732), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n732), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n835), .A2(new_n732), .ZN(new_n839));
  INV_X1    g414(.A(new_n832), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n835), .A2(new_n732), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n471), .B(G162), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(new_n627), .Z(new_n845));
  AOI21_X1  g420(.A(G37), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n838), .A2(KEYINPUT98), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(new_n832), .C1(new_n836), .C2(new_n837), .ZN(new_n849));
  INV_X1    g424(.A(new_n845), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n847), .A2(new_n849), .A3(new_n842), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n846), .A2(new_n851), .A3(KEYINPUT99), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g432(.A(G305), .B(G303), .ZN(new_n858));
  XNOR2_X1  g433(.A(G290), .B(G288), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n859), .A2(new_n860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n858), .B2(new_n862), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n557), .A2(new_n559), .A3(new_n599), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G299), .B2(new_n600), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n868), .B(new_n600), .C1(new_n605), .C2(new_n606), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n867), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n612), .B(new_n812), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT100), .B1(new_n607), .B2(new_n599), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n870), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n607), .A2(KEYINPUT101), .A3(new_n599), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n873), .A2(new_n875), .A3(new_n883), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n876), .A2(new_n870), .B1(new_n607), .B2(new_n599), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(new_n875), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n866), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n892), .A2(new_n888), .A3(new_n865), .ZN(new_n893));
  OAI21_X1  g468(.A(G868), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(G868), .B2(new_n809), .ZN(G331));
  XNOR2_X1  g470(.A(G331), .B(KEYINPUT103), .ZN(G295));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT104), .B1(new_n519), .B2(new_n521), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g474(.A1(G171), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n812), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n898), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n811), .A3(new_n810), .ZN(new_n903));
  AOI21_X1  g478(.A(G168), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n903), .A3(G168), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n897), .B1(new_n907), .B2(new_n885), .ZN(new_n908));
  INV_X1    g483(.A(new_n906), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(new_n904), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n872), .A3(KEYINPUT106), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n873), .A2(new_n883), .A3(new_n907), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n873), .A2(new_n883), .A3(KEYINPUT105), .A4(new_n907), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n865), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n877), .A2(new_n881), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n910), .A2(new_n882), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n865), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n885), .B1(new_n910), .B2(new_n882), .ZN(new_n924));
  AOI21_X1  g499(.A(G37), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(new_n917), .B2(new_n865), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(KEYINPUT107), .B(new_n927), .C1(new_n917), .C2(new_n865), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n919), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n926), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n918), .B2(new_n925), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n931), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n936), .B2(new_n920), .ZN(new_n937));
  MUX2_X1   g512(.A(new_n934), .B(new_n937), .S(KEYINPUT44), .Z(G397));
  XNOR2_X1  g513(.A(KEYINPUT108), .B(G1384), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n488), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT45), .B1(new_n941), .B2(KEYINPUT109), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(KEYINPUT109), .B2(new_n941), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n465), .A2(G40), .A3(new_n470), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n834), .ZN(new_n946));
  INV_X1    g521(.A(G1996), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT111), .Z(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n947), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT110), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n761), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n769), .B(G2067), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n949), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n715), .B(new_n718), .Z(new_n957));
  NAND2_X1  g532(.A1(new_n945), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(G290), .B(G1986), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n945), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n944), .ZN(new_n962));
  AOI21_X1  g537(.A(G1384), .B1(new_n485), .B2(new_n487), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(G8), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT113), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n687), .A2(G1976), .ZN(new_n967));
  INV_X1    g542(.A(G1976), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT52), .B1(G288), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT114), .ZN(new_n971));
  OR2_X1    g546(.A1(G305), .A2(G1981), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n575), .A2(new_n569), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(G1981), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT115), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n975), .A2(KEYINPUT116), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n978), .A2(new_n966), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n974), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT116), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT49), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n966), .A2(new_n967), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n979), .A2(new_n983), .B1(new_n984), .B2(KEYINPUT52), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n971), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G8), .ZN(new_n987));
  NOR2_X1   g562(.A1(G166), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT55), .ZN(new_n989));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n488), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n488), .A2(KEYINPUT45), .A3(new_n940), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n962), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1971), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n944), .B1(new_n963), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G2090), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n989), .B1(new_n1003), .B2(G8), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(KEYINPUT117), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1000), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(KEYINPUT112), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n991), .A2(new_n1008), .A3(KEYINPUT50), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n1001), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n987), .B1(new_n1011), .B2(new_n997), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n989), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1004), .A2(KEYINPUT117), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1005), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n986), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n993), .A2(new_n962), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n991), .A2(new_n992), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(G2078), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n995), .B2(G2078), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1024), .B(new_n1025), .C1(G1961), .C2(new_n1010), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1018), .B1(new_n1026), .B2(G301), .ZN(new_n1027));
  AND4_X1   g602(.A1(G40), .A2(new_n470), .A3(new_n463), .A4(new_n1023), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n994), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n943), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n1025), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1008), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n963), .A2(KEYINPUT112), .A3(new_n999), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1000), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT123), .B1(new_n1034), .B2(new_n749), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(KEYINPUT123), .A3(new_n749), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1031), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT124), .ZN(new_n1039));
  OAI21_X1  g614(.A(G171), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1030), .A2(new_n1025), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1037), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1041), .B(new_n1039), .C1(new_n1042), .C2(new_n1035), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1027), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1038), .A2(G301), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1026), .A2(G171), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1018), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1966), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(G2084), .B2(new_n1034), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G8), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT122), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G168), .A2(new_n987), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n1051), .B2(G8), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1053), .B(new_n1055), .C1(KEYINPUT122), .C2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1056), .B(G8), .C1(new_n1051), .C2(G286), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1051), .A2(KEYINPUT121), .A3(new_n1054), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT121), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1045), .A2(new_n1048), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(new_n556), .B(KEYINPUT57), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n998), .A2(new_n1000), .ZN(new_n1066));
  INV_X1    g641(.A(G1956), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT56), .B(G2072), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n993), .A2(new_n962), .A3(new_n994), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI22_X1  g647(.A1(new_n1010), .A2(G1348), .B1(G2067), .B2(new_n964), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n964), .A2(G2067), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1034), .B2(new_n787), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n599), .B1(new_n1077), .B2(KEYINPUT60), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n993), .A2(new_n947), .A3(new_n962), .A4(new_n994), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n964), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1082), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n528), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1075), .A2(new_n1078), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1077), .A2(KEYINPUT60), .ZN(new_n1089));
  INV_X1    g664(.A(new_n528), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT119), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1092), .B2(new_n1083), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n599), .A2(new_n1089), .B1(new_n1093), .B2(KEYINPUT59), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1068), .A2(new_n1065), .A3(new_n1070), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1071), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1071), .B2(new_n1096), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1088), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1072), .B1(new_n1101), .B2(new_n1098), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1095), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1073), .A2(new_n600), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1064), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1057), .A2(KEYINPUT122), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OR3_X1    g684(.A1(new_n1109), .A2(KEYINPUT62), .A3(new_n1062), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT62), .B1(new_n1109), .B2(new_n1062), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1047), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1017), .B1(new_n1106), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n986), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1013), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n979), .A2(new_n983), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(new_n968), .A3(new_n687), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n972), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1115), .A2(new_n1116), .B1(new_n1119), .B2(new_n966), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1052), .A2(G286), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1121), .B(KEYINPUT118), .Z(new_n1122));
  NOR2_X1   g697(.A1(new_n1012), .A2(new_n989), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1116), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1122), .A2(new_n1115), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT63), .B1(new_n1016), .B2(new_n1122), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n961), .B1(new_n1114), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n716), .A2(new_n718), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n955), .A2(new_n1130), .B1(G2067), .B2(new_n769), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n945), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n946), .A2(new_n954), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT125), .Z(new_n1134));
  INV_X1    g709(.A(KEYINPUT46), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n951), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n951), .A2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT47), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n945), .A2(new_n677), .A3(new_n582), .A4(new_n586), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT48), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n956), .A2(new_n958), .A3(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1132), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1129), .A2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n1146));
  INV_X1    g720(.A(G319), .ZN(new_n1147));
  NOR2_X1   g721(.A1(G227), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g722(.A(new_n1148), .B(KEYINPUT126), .ZN(new_n1149));
  NOR2_X1   g723(.A1(new_n1149), .A2(G401), .ZN(new_n1150));
  NAND2_X1  g724(.A1(new_n683), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g725(.A(new_n1151), .B1(new_n854), .B2(new_n855), .ZN(new_n1152));
  AND3_X1   g726(.A1(new_n934), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g727(.A(new_n1146), .B1(new_n934), .B2(new_n1152), .ZN(new_n1154));
  NOR2_X1   g728(.A1(new_n1153), .A2(new_n1154), .ZN(G308));
  NAND2_X1  g729(.A1(new_n934), .A2(new_n1152), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n1156), .A2(KEYINPUT127), .ZN(new_n1157));
  NAND3_X1  g731(.A1(new_n934), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1158));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1158), .ZN(G225));
endmodule


