//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n187));
  INV_X1    g001(.A(G107), .ZN(new_n188));
  NAND4_X1  g002(.A1(new_n188), .A2(KEYINPUT78), .A3(KEYINPUT3), .A4(G104), .ZN(new_n189));
  AND3_X1   g003(.A1(new_n188), .A2(KEYINPUT78), .A3(G104), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n191), .B1(new_n188), .B2(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n189), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G107), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n188), .A2(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n191), .B(new_n197), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(G101), .A3(new_n189), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n195), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT0), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n204), .A2(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n204), .A2(new_n206), .A3(new_n210), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT67), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n204), .A2(new_n206), .A3(new_n210), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n214), .B(new_n215), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n200), .A2(new_n221), .A3(G101), .A4(new_n189), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n213), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n187), .B1(new_n202), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n220), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n205), .A2(G143), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n203), .A2(G146), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n226), .A2(new_n227), .B1(new_n216), .B2(new_n217), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n215), .B1(new_n228), .B2(new_n214), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n195), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n230), .A2(KEYINPUT79), .A3(new_n231), .A4(new_n222), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G134), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G137), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT11), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT64), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n235), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n234), .A2(G137), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n242), .A2(new_n243), .B1(KEYINPUT64), .B2(new_n238), .ZN(new_n244));
  OAI21_X1  g058(.A(G131), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n237), .A2(new_n239), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n242), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n241), .A2(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n239), .B1(new_n235), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n251), .A3(KEYINPUT65), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(G131), .C1(new_n240), .C2(new_n244), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n203), .B(G146), .C1(new_n208), .C2(KEYINPUT1), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n208), .A2(new_n205), .A3(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(KEYINPUT66), .A3(new_n257), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n219), .A2(new_n262), .A3(G128), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT80), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n198), .A2(new_n197), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n188), .A2(G104), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n194), .B1(new_n267), .B2(KEYINPUT80), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n193), .A2(new_n194), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT10), .ZN(new_n271));
  INV_X1    g085(.A(new_n258), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n263), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n271), .B1(KEYINPUT10), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n233), .A2(new_n255), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n264), .A2(new_n269), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n268), .A2(new_n266), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n273), .A2(new_n195), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT12), .B1(new_n280), .B2(new_n255), .ZN(new_n281));
  INV_X1    g095(.A(new_n255), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n274), .B1(new_n264), .B2(new_n269), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT12), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n276), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(G110), .B(G140), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G227), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n287), .B(new_n289), .Z(new_n290));
  OAI21_X1  g104(.A(KEYINPUT82), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n281), .A2(new_n285), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT82), .ZN(new_n294));
  INV_X1    g108(.A(new_n290), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .A4(new_n276), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n233), .A2(new_n255), .A3(new_n275), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n255), .B1(new_n233), .B2(new_n275), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n291), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G469), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n297), .B2(new_n292), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n276), .A2(KEYINPUT81), .A3(new_n281), .A4(new_n285), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n290), .A3(new_n308), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n297), .A2(new_n298), .A3(new_n290), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n303), .B(new_n305), .C1(new_n301), .C2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(G116), .B(G119), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT2), .B(G113), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n316), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n314), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n231), .A2(new_n320), .A3(new_n222), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(KEYINPUT5), .ZN(new_n322));
  INV_X1    g136(.A(G116), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n323), .A2(KEYINPUT5), .A3(G119), .ZN(new_n324));
  INV_X1    g138(.A(G113), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n322), .A2(new_n326), .B1(new_n318), .B2(new_n314), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n269), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G122), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n321), .A2(new_n330), .A3(new_n328), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(KEYINPUT6), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n228), .B2(new_n214), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n264), .B2(new_n335), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n288), .A2(G224), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n337), .B(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n330), .B1(new_n321), .B2(new_n328), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n341), .A2(KEYINPUT83), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT83), .B1(new_n341), .B2(new_n342), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n334), .B(new_n340), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(G210), .B1(G237), .B2(G902), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT86), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT7), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(new_n339), .B2(KEYINPUT85), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(KEYINPUT85), .B2(new_n339), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n337), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n330), .B(KEYINPUT8), .ZN(new_n353));
  INV_X1    g167(.A(new_n328), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n269), .A2(new_n327), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n339), .B1(new_n357), .B2(new_n349), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n357), .B2(new_n349), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n337), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n352), .A2(new_n356), .A3(new_n333), .A4(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n361), .A2(new_n302), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n345), .A2(new_n348), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n348), .B1(new_n345), .B2(new_n362), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G952), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n368), .A2(KEYINPUT95), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(KEYINPUT95), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n288), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(G234), .B2(G237), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT21), .B(G898), .ZN(new_n373));
  AOI211_X1 g187(.A(new_n302), .B(new_n288), .C1(G234), .C2(G237), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n365), .A2(new_n367), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G221), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT9), .B(G234), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n379), .B2(new_n302), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n380), .B(KEYINPUT77), .Z(new_n381));
  XNOR2_X1  g195(.A(G128), .B(G143), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n234), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n208), .A2(G143), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT13), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G134), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(new_n385), .A3(G134), .A4(new_n384), .ZN(new_n388));
  INV_X1    g202(.A(G122), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT90), .B1(new_n389), .B2(G116), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n323), .A3(G122), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n323), .A2(G122), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n188), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n393), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n397), .A2(G107), .A3(new_n394), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n387), .B(new_n388), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G217), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n378), .A2(new_n400), .A3(G953), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n394), .B1(new_n393), .B2(KEYINPUT14), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n402), .A2(KEYINPUT91), .B1(new_n403), .B2(new_n397), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n390), .B2(new_n392), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n394), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n188), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n382), .B(G134), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n398), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n399), .B(new_n401), .C1(new_n408), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT92), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n402), .A2(KEYINPUT91), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n397), .A2(new_n403), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n407), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G107), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n410), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n399), .A4(new_n401), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n399), .B1(new_n408), .B2(new_n411), .ZN(new_n421));
  INV_X1    g235(.A(new_n401), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n413), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT94), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n302), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT93), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n427), .A3(new_n302), .ZN(new_n428));
  INV_X1    g242(.A(G478), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT15), .ZN(new_n430));
  AOI22_X1  g244(.A1(KEYINPUT93), .A2(new_n426), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n426), .A2(KEYINPUT93), .A3(new_n430), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  NOR2_X1   g248(.A1(G237), .A2(G953), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(G143), .A3(G214), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G143), .B1(new_n435), .B2(G214), .ZN(new_n438));
  OAI21_X1  g252(.A(G131), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT17), .ZN(new_n440));
  INV_X1    g254(.A(G237), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n288), .A3(G214), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n203), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n250), .A3(new_n436), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n436), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT17), .A3(G131), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT74), .A2(G125), .ZN(new_n448));
  INV_X1    g262(.A(G140), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(KEYINPUT74), .A2(G125), .A3(G140), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(KEYINPUT16), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT16), .B1(new_n449), .B2(G125), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n205), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n454), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G146), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n445), .A2(new_n447), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n451), .ZN(new_n459));
  AOI21_X1  g273(.A(G140), .B1(KEYINPUT74), .B2(G125), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G146), .ZN(new_n462));
  XNOR2_X1  g276(.A(G125), .B(G140), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT76), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n463), .A2(new_n464), .A3(new_n205), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n464), .B1(new_n463), .B2(new_n205), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(KEYINPUT18), .A2(G131), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n443), .A2(new_n436), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n446), .A2(KEYINPUT18), .A3(G131), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(G113), .B(G122), .Z(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT88), .B(G104), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n458), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n457), .A2(KEYINPUT75), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT75), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n456), .A2(new_n477), .A3(G146), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n461), .A2(KEYINPUT19), .ZN(new_n479));
  XOR2_X1   g293(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n463), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n481), .A3(new_n205), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n439), .A2(new_n444), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n476), .A2(new_n478), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n474), .B1(new_n484), .B2(new_n471), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n433), .B(new_n434), .C1(new_n475), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT89), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n475), .A2(new_n485), .ZN(new_n488));
  INV_X1    g302(.A(new_n434), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT20), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n458), .A2(new_n471), .A3(new_n474), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n483), .A2(new_n482), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n477), .B1(new_n456), .B2(G146), .ZN(new_n493));
  AOI211_X1 g307(.A(KEYINPUT75), .B(new_n205), .C1(new_n452), .C2(new_n454), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n470), .A2(new_n469), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n492), .A2(new_n495), .B1(new_n496), .B2(new_n467), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n491), .B1(new_n497), .B2(new_n474), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n433), .A4(new_n434), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n487), .A2(new_n490), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n474), .B1(new_n458), .B2(new_n471), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n302), .B1(new_n475), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G475), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n431), .A2(new_n432), .A3(new_n505), .ZN(new_n506));
  AND4_X1   g320(.A1(new_n313), .A2(new_n376), .A3(new_n381), .A4(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT23), .ZN(new_n508));
  INV_X1    g322(.A(G119), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n508), .B1(new_n509), .B2(G128), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n510), .B(new_n511), .C1(G119), .C2(new_n208), .ZN(new_n512));
  XNOR2_X1  g326(.A(G119), .B(G128), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT24), .B(G110), .Z(new_n514));
  OAI22_X1  g328(.A1(new_n512), .A2(G110), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n495), .B(new_n515), .C1(new_n465), .C2(new_n466), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n513), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n517), .B(KEYINPUT73), .Z(new_n518));
  NAND2_X1  g332(.A1(new_n457), .A2(new_n455), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n512), .A2(G110), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT22), .B(G137), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n516), .A2(new_n521), .A3(new_n525), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n302), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n400), .B1(G234), .B2(new_n302), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n527), .A2(new_n528), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n532), .A2(G902), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n531), .A2(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n230), .A2(new_n252), .A3(new_n254), .ZN(new_n538));
  OAI21_X1  g352(.A(G131), .B1(new_n235), .B2(new_n248), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n264), .A2(new_n251), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n320), .ZN(new_n542));
  INV_X1    g356(.A(new_n320), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n538), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT28), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n542), .B2(new_n544), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(new_n546), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT26), .B(G101), .Z(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT69), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n435), .A2(G210), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT29), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n550), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT29), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n538), .A2(KEYINPUT28), .A3(new_n543), .A4(new_n540), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n228), .A2(new_n214), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n252), .A2(new_n254), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n540), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n320), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n549), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n556), .B(new_n557), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n562), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n538), .A2(KEYINPUT30), .A3(new_n540), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n320), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n559), .B1(new_n574), .B2(new_n544), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n302), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G472), .B1(new_n561), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n559), .A3(new_n544), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT70), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(KEYINPUT31), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n569), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n574), .A2(new_n559), .A3(new_n544), .A4(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(G472), .A2(G902), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(KEYINPUT32), .A3(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n577), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n588), .ZN(new_n591));
  NOR2_X1   g405(.A1(KEYINPUT71), .A2(KEYINPUT32), .ZN(new_n592));
  AND2_X1   g406(.A1(KEYINPUT71), .A2(KEYINPUT32), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n537), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n507), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT96), .B(G101), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G3));
  AND2_X1   g412(.A1(new_n313), .A2(new_n381), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n345), .A2(new_n348), .A3(new_n362), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n366), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n345), .A2(new_n362), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n347), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n601), .A3(new_n600), .ZN(new_n606));
  INV_X1    g420(.A(new_n375), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(G478), .B1(new_n424), .B2(new_n302), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n421), .B2(new_n422), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n424), .A2(new_n610), .B1(new_n412), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n429), .A2(G902), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n505), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n608), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n587), .A2(new_n302), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G472), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n591), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n537), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n599), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  NOR2_X1   g439(.A1(new_n431), .A2(new_n432), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n490), .A2(new_n486), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n504), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n608), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n599), .A2(new_n629), .A3(new_n621), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n526), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n522), .B(new_n633), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n531), .A2(new_n532), .B1(new_n535), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n620), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n507), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  AOI21_X1  g453(.A(new_n602), .B1(new_n365), .B2(new_n601), .ZN(new_n640));
  INV_X1    g454(.A(new_n635), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n313), .A2(new_n381), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n426), .A2(KEYINPUT93), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n428), .A2(new_n430), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n426), .A2(KEYINPUT93), .A3(new_n430), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n372), .B1(new_n648), .B2(new_n374), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n628), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n590), .B2(new_n594), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  XNOR2_X1  g468(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n649), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n599), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n545), .A2(new_n569), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n545), .A2(new_n569), .A3(KEYINPUT99), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n664), .A2(new_n578), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n666), .B2(G902), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(new_n589), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n594), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n365), .B(KEYINPUT38), .Z(new_n670));
  NOR2_X1   g484(.A1(new_n641), .A2(new_n367), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n501), .A2(new_n504), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n645), .B2(new_n646), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n669), .B(new_n670), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n675), .B2(new_n674), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n660), .A2(new_n661), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  INV_X1    g493(.A(new_n649), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n615), .A2(new_n505), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n590), .B2(new_n594), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n642), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  NAND2_X1  g498(.A1(new_n300), .A2(new_n302), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  INV_X1    g500(.A(new_n380), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n303), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n595), .A2(new_n617), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  NAND3_X1  g506(.A1(new_n595), .A2(new_n629), .A3(new_n689), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  NAND2_X1  g508(.A1(new_n603), .A2(new_n606), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n590), .A2(new_n594), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n635), .A2(new_n375), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(new_n697), .A3(new_n506), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  NAND4_X1  g514(.A1(new_n686), .A2(new_n303), .A3(new_n687), .A4(new_n607), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n505), .B1(new_n431), .B2(new_n432), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n702), .B1(new_n695), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n640), .A2(new_n673), .A3(KEYINPUT106), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT104), .B(G472), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n618), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n588), .B(KEYINPUT103), .ZN(new_n709));
  INV_X1    g523(.A(new_n552), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n551), .A2(new_n546), .B1(new_n548), .B2(new_n544), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n559), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n582), .A2(new_n586), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n708), .A2(new_n714), .A3(new_n536), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n708), .A2(new_n714), .A3(KEYINPUT105), .A4(new_n536), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n706), .A2(new_n719), .A3(KEYINPUT107), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT107), .B1(new_n706), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n389), .ZN(G24));
  INV_X1    g537(.A(new_n714), .ZN(new_n724));
  INV_X1    g538(.A(new_n707), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n587), .B2(new_n302), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n724), .A2(new_n635), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n681), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n696), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT108), .B(G125), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G27));
  NOR2_X1   g545(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n309), .A2(KEYINPUT109), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n295), .B1(new_n286), .B2(new_n306), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n308), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n301), .B(new_n310), .C1(new_n734), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n303), .A2(new_n305), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n733), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n309), .A2(KEYINPUT109), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n736), .B1(new_n735), .B2(new_n308), .ZN(new_n742));
  OAI211_X1 g556(.A(G469), .B(new_n311), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(KEYINPUT110), .A3(new_n303), .A4(new_n305), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n740), .A2(new_n687), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n743), .A2(new_n303), .A3(new_n305), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n380), .B1(new_n748), .B2(new_n733), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT111), .A3(new_n744), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n365), .A2(new_n366), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AND4_X1   g566(.A1(KEYINPUT112), .A2(new_n747), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n751), .B1(new_n745), .B2(new_n746), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT112), .B1(new_n754), .B2(new_n750), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n595), .B(new_n732), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT32), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n591), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n537), .B1(new_n590), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n728), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n747), .A2(new_n750), .A3(new_n752), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n754), .A2(KEYINPUT112), .A3(new_n750), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n756), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n250), .ZN(G33));
  INV_X1    g582(.A(new_n651), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n595), .B(new_n769), .C1(new_n753), .C2(new_n755), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n615), .A2(new_n672), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n620), .A2(new_n641), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n752), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT45), .B(new_n311), .C1(new_n741), .C2(new_n742), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n301), .B1(new_n312), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n304), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(KEYINPUT46), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n303), .B1(new_n783), .B2(KEYINPUT46), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n687), .B(new_n656), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n776), .A2(new_n772), .A3(new_n777), .ZN(new_n787));
  OR3_X1    g601(.A1(new_n779), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  INV_X1    g603(.A(new_n697), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n728), .A3(new_n537), .A4(new_n752), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n784), .A2(new_n785), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n687), .ZN(new_n793));
  XNOR2_X1  g607(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n687), .A3(new_n794), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n791), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n449), .ZN(G42));
  NAND2_X1  g613(.A1(new_n686), .A2(new_n303), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT49), .Z(new_n801));
  INV_X1    g615(.A(new_n669), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n536), .A2(new_n381), .A3(new_n366), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n670), .A2(new_n773), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n774), .A2(new_n372), .A3(new_n775), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n688), .A2(new_n751), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT114), .Z(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(KEYINPUT48), .A3(new_n759), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT48), .B1(new_n809), .B2(new_n759), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n806), .A2(new_n719), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n696), .ZN(new_n814));
  INV_X1    g628(.A(new_n371), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n802), .A2(new_n536), .A3(new_n372), .A4(new_n807), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n814), .B(new_n815), .C1(new_n616), .C2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n810), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n796), .B(new_n797), .C1(new_n381), .C2(new_n800), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n812), .A2(new_n751), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n816), .A2(new_n505), .A3(new_n615), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n809), .B2(new_n727), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n670), .A2(new_n688), .A3(new_n366), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n813), .A2(KEYINPUT50), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT50), .B1(new_n813), .B2(new_n825), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n822), .B(new_n828), .C1(KEYINPUT115), .C2(KEYINPUT51), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n830));
  INV_X1    g644(.A(new_n821), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n819), .B2(KEYINPUT116), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(KEYINPUT116), .B2(new_n819), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n820), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n818), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n724), .A2(new_n681), .A3(new_n635), .A4(new_n726), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n753), .B2(new_n755), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n595), .B(new_n689), .C1(new_n617), .C2(new_n629), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n507), .B1(new_n595), .B2(new_n636), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n506), .B1(new_n505), .B2(new_n614), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n599), .A2(new_n621), .A3(new_n376), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n838), .A2(new_n839), .A3(new_n699), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n599), .A2(new_n641), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n752), .A2(new_n626), .A3(new_n650), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n843), .A2(new_n790), .A3(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n722), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n653), .A2(new_n683), .A3(new_n729), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n704), .A2(new_n705), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n635), .A2(new_n680), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n668), .B2(new_n594), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n749), .A2(new_n849), .A3(new_n851), .A4(new_n744), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n847), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n696), .A2(new_n836), .B1(new_n642), .B2(new_n652), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .A3(new_n683), .A4(new_n852), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n770), .A2(new_n837), .A3(new_n846), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n595), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n763), .B2(new_n764), .ZN(new_n860));
  INV_X1    g674(.A(new_n760), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(new_n753), .B2(new_n755), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n860), .A2(new_n732), .B1(new_n862), .B2(KEYINPUT42), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT53), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n770), .A2(new_n837), .A3(new_n846), .A4(new_n857), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n865), .A2(new_n767), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT54), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n858), .A2(KEYINPUT53), .A3(new_n863), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n866), .B1(new_n865), .B2(new_n767), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n835), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n805), .B1(new_n874), .B2(new_n875), .ZN(G75));
  NOR2_X1   g690(.A1(new_n288), .A2(G952), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n302), .B1(new_n869), .B2(new_n871), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(new_n347), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n334), .B1(new_n343), .B2(new_n344), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n340), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT55), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n878), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n880), .A2(new_n883), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n880), .A2(KEYINPUT117), .A3(new_n883), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(G51));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n869), .A2(new_n871), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(KEYINPUT54), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n873), .B2(new_n890), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n304), .B(KEYINPUT57), .Z(new_n894));
  OAI21_X1  g708(.A(new_n300), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n879), .A2(new_n780), .A3(new_n782), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n877), .B1(new_n895), .B2(new_n896), .ZN(G54));
  NAND2_X1  g711(.A1(KEYINPUT58), .A2(G475), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT119), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n879), .A2(new_n498), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n498), .B1(new_n879), .B2(new_n899), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n900), .A2(new_n901), .A3(new_n877), .ZN(G60));
  XNOR2_X1  g716(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n429), .A2(new_n302), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n903), .B(new_n904), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n868), .B2(new_n872), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n878), .B1(new_n907), .B2(new_n612), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n612), .A2(new_n905), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n909), .B1(new_n893), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n910), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT118), .B1(new_n868), .B2(new_n872), .ZN(new_n913));
  OAI211_X1 g727(.A(KEYINPUT121), .B(new_n912), .C1(new_n913), .C2(new_n892), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n908), .B1(new_n911), .B2(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT60), .Z(new_n917));
  AND2_X1   g731(.A1(new_n891), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n877), .B1(new_n918), .B2(new_n634), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n891), .A2(new_n917), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n533), .B(KEYINPUT122), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n919), .B2(new_n922), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(G66));
  NOR2_X1   g740(.A1(new_n722), .A2(new_n842), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(G224), .A2(G953), .ZN(new_n929));
  OAI22_X1  g743(.A1(new_n928), .A2(G953), .B1(new_n373), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n881), .B1(G898), .B2(new_n288), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n930), .B(new_n931), .Z(G69));
  INV_X1    g746(.A(new_n678), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT62), .B1(new_n933), .B2(new_n848), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n935));
  INV_X1    g749(.A(new_n848), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n678), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n788), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n595), .A2(new_n752), .A3(new_n840), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n659), .A2(new_n939), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n798), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n934), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n288), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n572), .A2(new_n573), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n479), .A2(new_n481), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT125), .Z(new_n948));
  NAND2_X1  g762(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n288), .A2(G900), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT126), .ZN(new_n951));
  INV_X1    g765(.A(new_n798), .ZN(new_n952));
  INV_X1    g766(.A(new_n786), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n849), .A3(new_n759), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n788), .A2(new_n954), .A3(new_n936), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n863), .A2(new_n770), .A3(new_n952), .A4(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n951), .B1(new_n956), .B2(new_n288), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(KEYINPUT127), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n947), .B1(new_n957), .B2(KEYINPUT127), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n949), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n288), .B1(G227), .B2(G900), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n942), .B2(new_n928), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n574), .A2(new_n544), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(new_n569), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n569), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n956), .A2(new_n928), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n964), .ZN(new_n972));
  INV_X1    g786(.A(new_n968), .ZN(new_n973));
  AND4_X1   g787(.A1(new_n891), .A2(new_n970), .A3(new_n964), .A4(new_n973), .ZN(new_n974));
  NOR4_X1   g788(.A1(new_n969), .A2(new_n972), .A3(new_n974), .A4(new_n877), .ZN(G57));
endmodule


