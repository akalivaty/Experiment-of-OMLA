

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  XNOR2_X1 U324 ( .A(n313), .B(n312), .ZN(n377) );
  XOR2_X1 U325 ( .A(G78GAT), .B(G148GAT), .Z(n313) );
  XNOR2_X1 U326 ( .A(n293), .B(n314), .ZN(n369) );
  NOR2_X4 U327 ( .A1(n537), .A2(n476), .ZN(n569) );
  XNOR2_X1 U328 ( .A(n443), .B(n365), .ZN(n368) );
  XNOR2_X1 U329 ( .A(n448), .B(KEYINPUT106), .ZN(n449) );
  XNOR2_X1 U330 ( .A(n579), .B(n457), .ZN(n553) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U332 ( .A(G64GAT), .B(G92GAT), .Z(n293) );
  INV_X1 U333 ( .A(KEYINPUT95), .ZN(n363) );
  XNOR2_X1 U334 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U335 ( .A(G99GAT), .B(G85GAT), .Z(n430) );
  XNOR2_X1 U336 ( .A(n436), .B(n292), .ZN(n437) );
  INV_X1 U337 ( .A(KEYINPUT37), .ZN(n448) );
  XNOR2_X1 U338 ( .A(n438), .B(n437), .ZN(n442) );
  XNOR2_X1 U339 ( .A(n450), .B(n449), .ZN(n519) );
  XOR2_X1 U340 ( .A(KEYINPUT36), .B(n545), .Z(n587) );
  XOR2_X1 U341 ( .A(n446), .B(n445), .Z(n545) );
  XOR2_X1 U342 ( .A(n374), .B(n373), .Z(n523) );
  XNOR2_X1 U343 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U344 ( .A(n454), .B(KEYINPUT40), .ZN(n455) );
  XNOR2_X1 U345 ( .A(n480), .B(n479), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT67), .B(KEYINPUT20), .Z(n295) );
  XNOR2_X1 U348 ( .A(G190GAT), .B(KEYINPUT86), .ZN(n294) );
  XOR2_X1 U349 ( .A(n295), .B(n294), .Z(n310) );
  XOR2_X1 U350 ( .A(G176GAT), .B(G183GAT), .Z(n297) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n299) );
  INV_X1 U353 ( .A(G71GAT), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n305) );
  XOR2_X1 U355 ( .A(G120GAT), .B(KEYINPUT0), .Z(n301) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(G134GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n404) );
  XOR2_X1 U358 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n303) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n370) );
  XNOR2_X1 U361 ( .A(n404), .B(n370), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G127GAT), .Z(n347) );
  XOR2_X1 U364 ( .A(n306), .B(n347), .Z(n308) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(G99GAT), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n494) );
  INV_X1 U368 ( .A(n494), .ZN(n537) );
  XNOR2_X1 U369 ( .A(G71GAT), .B(G57GAT), .ZN(n311) );
  XOR2_X1 U370 ( .A(n311), .B(KEYINPUT13), .Z(n346) );
  XNOR2_X1 U371 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n312) );
  XNOR2_X1 U372 ( .A(G176GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n377), .B(n369), .ZN(n319) );
  XOR2_X1 U374 ( .A(KEYINPUT32), .B(KEYINPUT79), .Z(n316) );
  NAND2_X1 U375 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U377 ( .A(n317), .B(KEYINPUT33), .Z(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U379 ( .A(n320), .B(KEYINPUT31), .Z(n322) );
  XNOR2_X1 U380 ( .A(G120GAT), .B(n430), .ZN(n321) );
  XOR2_X1 U381 ( .A(n322), .B(n321), .Z(n323) );
  XNOR2_X1 U382 ( .A(n346), .B(n323), .ZN(n579) );
  XOR2_X1 U383 ( .A(KEYINPUT73), .B(KEYINPUT30), .Z(n325) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(KEYINPUT72), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n343) );
  XOR2_X1 U386 ( .A(G141GAT), .B(G22GAT), .Z(n327) );
  XNOR2_X1 U387 ( .A(G50GAT), .B(G36GAT), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U389 ( .A(G113GAT), .B(G15GAT), .Z(n329) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(G197GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U392 ( .A(n331), .B(n330), .Z(n341) );
  XOR2_X1 U393 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n333) );
  XNOR2_X1 U394 ( .A(KEYINPUT77), .B(KEYINPUT29), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n339) );
  XOR2_X1 U396 ( .A(G29GAT), .B(G43GAT), .Z(n335) );
  XNOR2_X1 U397 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n444) );
  XOR2_X1 U399 ( .A(KEYINPUT76), .B(G1GAT), .Z(n357) );
  XOR2_X1 U400 ( .A(n444), .B(n357), .Z(n337) );
  NAND2_X1 U401 ( .A1(G229GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U405 ( .A(n343), .B(n342), .ZN(n561) );
  AND2_X1 U406 ( .A1(n579), .A2(n561), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n344), .B(KEYINPUT80), .ZN(n487) );
  XOR2_X1 U408 ( .A(G8GAT), .B(G183GAT), .Z(n345) );
  XOR2_X1 U409 ( .A(G211GAT), .B(n345), .Z(n374) );
  XOR2_X1 U410 ( .A(n374), .B(n346), .Z(n361) );
  XOR2_X1 U411 ( .A(G22GAT), .B(G155GAT), .Z(n379) );
  XOR2_X1 U412 ( .A(n379), .B(n347), .Z(n349) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U415 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n351) );
  XNOR2_X1 U416 ( .A(KEYINPUT12), .B(KEYINPUT83), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U418 ( .A(n353), .B(n352), .Z(n359) );
  XOR2_X1 U419 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n355) );
  XNOR2_X1 U420 ( .A(G78GAT), .B(G64GAT), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n361), .B(n360), .ZN(n582) );
  XNOR2_X1 U425 ( .A(G36GAT), .B(G190GAT), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n362), .B(G218GAT), .ZN(n443) );
  NAND2_X1 U427 ( .A1(G226GAT), .A2(G233GAT), .ZN(n364) );
  XOR2_X1 U428 ( .A(G197GAT), .B(KEYINPUT21), .Z(n378) );
  XNOR2_X1 U429 ( .A(n378), .B(KEYINPUT94), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n366), .B(KEYINPUT96), .ZN(n367) );
  XOR2_X1 U431 ( .A(n368), .B(n367), .Z(n372) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  INV_X1 U434 ( .A(n523), .ZN(n492) );
  NAND2_X1 U435 ( .A1(n492), .A2(n494), .ZN(n393) );
  XOR2_X1 U436 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n376) );
  XNOR2_X1 U437 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n411) );
  XNOR2_X1 U439 ( .A(n411), .B(n377), .ZN(n392) );
  XOR2_X1 U440 ( .A(n379), .B(n378), .Z(n381) );
  NAND2_X1 U441 ( .A1(G228GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U443 ( .A(G50GAT), .B(G162GAT), .Z(n431) );
  XOR2_X1 U444 ( .A(n382), .B(n431), .Z(n390) );
  XOR2_X1 U445 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n384) );
  XNOR2_X1 U446 ( .A(G218GAT), .B(KEYINPUT89), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U448 ( .A(KEYINPUT87), .B(G211GAT), .Z(n386) );
  XNOR2_X1 U449 ( .A(KEYINPUT22), .B(G204GAT), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n474) );
  NAND2_X1 U454 ( .A1(n393), .A2(n474), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n394), .B(KEYINPUT25), .ZN(n395) );
  XNOR2_X1 U456 ( .A(KEYINPUT98), .B(n395), .ZN(n416) );
  XOR2_X1 U457 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n397) );
  XNOR2_X1 U458 ( .A(KEYINPUT92), .B(KEYINPUT4), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n415) );
  XOR2_X1 U460 ( .A(G155GAT), .B(G148GAT), .Z(n399) );
  XNOR2_X1 U461 ( .A(G29GAT), .B(G127GAT), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n401) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(G57GAT), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U466 ( .A(n403), .B(n402), .Z(n409) );
  XOR2_X1 U467 ( .A(G85GAT), .B(G162GAT), .Z(n406) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n404), .B(n407), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U472 ( .A(n410), .B(KEYINPUT6), .Z(n413) );
  XNOR2_X1 U473 ( .A(n411), .B(KEYINPUT91), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n489) );
  INV_X1 U476 ( .A(n489), .ZN(n530) );
  NAND2_X1 U477 ( .A1(n416), .A2(n530), .ZN(n427) );
  INV_X1 U478 ( .A(KEYINPUT26), .ZN(n419) );
  NOR2_X1 U479 ( .A1(n494), .A2(n474), .ZN(n417) );
  XNOR2_X1 U480 ( .A(KEYINPUT97), .B(n417), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n572) );
  NOR2_X1 U482 ( .A1(n489), .A2(n572), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n492), .B(KEYINPUT27), .ZN(n533) );
  INV_X1 U484 ( .A(n533), .ZN(n420) );
  NOR2_X1 U485 ( .A1(n421), .A2(n420), .ZN(n425) );
  XOR2_X1 U486 ( .A(n474), .B(KEYINPUT71), .Z(n422) );
  XOR2_X1 U487 ( .A(n422), .B(KEYINPUT28), .Z(n498) );
  NOR2_X1 U488 ( .A1(n494), .A2(n498), .ZN(n423) );
  OR2_X1 U489 ( .A1(n530), .A2(n423), .ZN(n424) );
  NAND2_X1 U490 ( .A1(n425), .A2(n424), .ZN(n426) );
  NAND2_X1 U491 ( .A1(n427), .A2(n426), .ZN(n428) );
  XOR2_X1 U492 ( .A(KEYINPUT99), .B(n428), .Z(n486) );
  NAND2_X1 U493 ( .A1(n582), .A2(n486), .ZN(n429) );
  XOR2_X1 U494 ( .A(KEYINPUT105), .B(n429), .Z(n447) );
  XOR2_X1 U495 ( .A(KEYINPUT68), .B(n430), .Z(n433) );
  XNOR2_X1 U496 ( .A(n431), .B(G92GAT), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n438) );
  XOR2_X1 U498 ( .A(KEYINPUT9), .B(KEYINPUT70), .Z(n435) );
  XNOR2_X1 U499 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U501 ( .A(KEYINPUT81), .B(KEYINPUT11), .Z(n440) );
  XNOR2_X1 U502 ( .A(G134GAT), .B(KEYINPUT66), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U504 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U505 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X1 U506 ( .A1(n447), .A2(n587), .ZN(n450) );
  NAND2_X1 U507 ( .A1(n487), .A2(n519), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n451) );
  XNOR2_X1 U509 ( .A(KEYINPUT38), .B(n451), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n505) );
  NOR2_X1 U511 ( .A1(n537), .A2(n505), .ZN(n456) );
  INV_X1 U512 ( .A(G43GAT), .ZN(n454) );
  INV_X1 U513 ( .A(n545), .ZN(n559) );
  XNOR2_X1 U514 ( .A(n582), .B(KEYINPUT115), .ZN(n568) );
  INV_X1 U515 ( .A(n561), .ZN(n574) );
  INV_X1 U516 ( .A(KEYINPUT41), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n574), .A2(n553), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n458), .B(KEYINPUT46), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n568), .A2(n459), .ZN(n460) );
  NAND2_X1 U520 ( .A1(n559), .A2(n460), .ZN(n461) );
  XNOR2_X1 U521 ( .A(KEYINPUT47), .B(n461), .ZN(n467) );
  NOR2_X1 U522 ( .A1(n582), .A2(n587), .ZN(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT69), .B(KEYINPUT45), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n463), .B(n462), .ZN(n465) );
  NAND2_X1 U525 ( .A1(n574), .A2(n579), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT64), .B(KEYINPUT116), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT48), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n470), .B(n469), .ZN(n531) );
  NOR2_X1 U531 ( .A1(n523), .A2(n531), .ZN(n471) );
  XNOR2_X1 U532 ( .A(KEYINPUT54), .B(n471), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n472), .A2(n530), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(KEYINPUT65), .ZN(n573) );
  NAND2_X1 U535 ( .A1(n573), .A2(n474), .ZN(n475) );
  XOR2_X1 U536 ( .A(KEYINPUT55), .B(n475), .Z(n476) );
  AND2_X1 U537 ( .A1(n569), .A2(n545), .ZN(n480) );
  XNOR2_X1 U538 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n478) );
  INV_X1 U539 ( .A(G190GAT), .ZN(n477) );
  XOR2_X1 U540 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n482) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n491) );
  NOR2_X1 U543 ( .A1(n545), .A2(n582), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n483), .B(KEYINPUT16), .ZN(n484) );
  XOR2_X1 U545 ( .A(KEYINPUT85), .B(n484), .Z(n485) );
  AND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n510) );
  NAND2_X1 U547 ( .A1(n510), .A2(n487), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT100), .B(n488), .Z(n499) );
  NAND2_X1 U549 ( .A1(n489), .A2(n499), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n499), .A2(n492), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U554 ( .A1(n494), .A2(n499), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U556 ( .A(G15GAT), .B(n497), .Z(G1326GAT) );
  INV_X1 U557 ( .A(n498), .ZN(n535) );
  NAND2_X1 U558 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n500), .B(KEYINPUT104), .ZN(n501) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n501), .ZN(G1327GAT) );
  NOR2_X1 U561 ( .A1(n530), .A2(n505), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n523), .A2(n505), .ZN(n504) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  NOR2_X1 U566 ( .A1(n535), .A2(n505), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n509) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT110), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(n512) );
  NOR2_X1 U572 ( .A1(n561), .A2(n553), .ZN(n520) );
  NAND2_X1 U573 ( .A1(n520), .A2(n510), .ZN(n516) );
  NOR2_X1 U574 ( .A1(n530), .A2(n516), .ZN(n511) );
  XOR2_X1 U575 ( .A(n512), .B(n511), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n516), .ZN(n513) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n537), .A2(n516), .ZN(n514) );
  XOR2_X1 U579 ( .A(KEYINPUT112), .B(n514), .Z(n515) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n515), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n535), .A2(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U585 ( .A1(n530), .A2(n527), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n527), .ZN(n524) );
  XOR2_X1 U589 ( .A(KEYINPUT114), .B(n524), .Z(n525) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n525), .ZN(G1337GAT) );
  NOR2_X1 U591 ( .A1(n537), .A2(n527), .ZN(n526) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n535), .A2(n527), .ZN(n528) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(KEYINPUT117), .B(n534), .ZN(n549) );
  NAND2_X1 U599 ( .A1(n549), .A2(n535), .ZN(n536) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n561), .A2(n546), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n540) );
  INV_X1 U604 ( .A(n553), .ZN(n564) );
  NAND2_X1 U605 ( .A1(n546), .A2(n564), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n543) );
  NAND2_X1 U609 ( .A1(n546), .A2(n568), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n549), .A2(n572), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n574), .A2(n558), .ZN(n550) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n552) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n553), .A2(n558), .ZN(n554) );
  XOR2_X1 U622 ( .A(n555), .B(n554), .Z(G1345GAT) );
  NOR2_X1 U623 ( .A1(n582), .A2(n558), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n569), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n566) );
  NAND2_X1 U632 ( .A1(n569), .A2(n564), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G176GAT), .ZN(G1349GAT) );
  XOR2_X1 U635 ( .A(G183GAT), .B(KEYINPUT123), .Z(n571) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1350GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n586) );
  NOR2_X1 U639 ( .A1(n586), .A2(n574), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n586), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n586), .ZN(n583) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n585) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n589) );
  NOR2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U653 ( .A(n589), .B(n588), .Z(G1355GAT) );
endmodule

