//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT4), .ZN(new_n207));
  NOR2_X1   g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR3_X1   g012(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n209), .B(new_n210), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(KEYINPUT76), .A3(new_n210), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT76), .ZN(new_n217));
  INV_X1    g016(.A(new_n210), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(new_n208), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT77), .ZN(new_n222));
  XOR2_X1   g021(.A(G155gat), .B(G162gat), .Z(new_n223));
  AND3_X1   g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n222), .B1(new_n221), .B2(new_n223), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n215), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT70), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G127gat), .B(G134gat), .Z(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n228), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(KEYINPUT1), .B2(new_n227), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n230), .B(KEYINPUT69), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n207), .B1(new_n226), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n215), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n223), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT77), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n238), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n238), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n249), .B(new_n215), .C1(new_n224), .C2(new_n225), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n248), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n245), .B1(new_n226), .B2(KEYINPUT3), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT78), .A3(new_n251), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n247), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT5), .ZN(new_n257));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n260));
  INV_X1    g059(.A(new_n247), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n250), .A2(new_n248), .A3(new_n252), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT78), .B1(new_n254), .B2(new_n251), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n258), .B(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n226), .B(new_n238), .ZN(new_n265));
  INV_X1    g064(.A(new_n258), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n257), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n259), .A2(new_n260), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n260), .A3(new_n267), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n206), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G8gat), .B(G36gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n278), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT66), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(G183gat), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT64), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT66), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(KEYINPUT25), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n282), .B(new_n292), .C1(new_n281), .C2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT67), .B(G190gat), .ZN(new_n296));
  AOI211_X1 g095(.A(new_n287), .B(new_n283), .C1(new_n296), .C2(new_n284), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT25), .B1(new_n297), .B2(new_n281), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT27), .B(G183gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G169gat), .ZN(new_n304));
  INV_X1    g103(.A(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(G183gat), .B2(G190gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n296), .A2(new_n299), .A3(new_n301), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n307), .A3(new_n280), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n303), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n298), .A3(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n313), .A2(G226gat), .A3(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n313), .A2(new_n315), .B1(G226gat), .B2(G233gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G211gat), .B(G218gat), .Z(new_n318));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G211gat), .B(G218gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G197gat), .B(G204gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT22), .ZN(new_n325));
  INV_X1    g124(.A(G211gat), .ZN(new_n326));
  INV_X1    g125(.A(G218gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n320), .A2(new_n328), .A3(new_n324), .A4(new_n322), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n332), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n314), .B2(new_n316), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n275), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT30), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n274), .B(KEYINPUT75), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n333), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n336), .B2(KEYINPUT30), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT40), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n256), .A2(new_n258), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT39), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n206), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n265), .A2(new_n266), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT39), .B(new_n347), .C1(new_n256), .C2(new_n258), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n343), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n262), .A2(new_n263), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n345), .B(new_n266), .C1(new_n350), .C2(new_n247), .ZN(new_n351));
  AND4_X1   g150(.A1(new_n343), .A2(new_n348), .A3(new_n351), .A4(new_n205), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n271), .B(new_n342), .C1(new_n349), .C2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n348), .A2(new_n351), .A3(new_n205), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT40), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n346), .A2(new_n343), .A3(new_n348), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n359), .A2(KEYINPUT83), .A3(new_n271), .A4(new_n342), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n260), .B1(new_n264), .B2(KEYINPUT5), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n264), .A2(new_n267), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n205), .A3(new_n269), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n271), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT38), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n333), .A2(new_n335), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT37), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT37), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  AND4_X1   g172(.A1(new_n368), .A2(new_n371), .A3(new_n373), .A4(new_n339), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n274), .B1(new_n369), .B2(new_n372), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n368), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n374), .A2(new_n376), .A3(new_n336), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT6), .B(new_n206), .C1(new_n268), .C2(new_n270), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n378), .A2(KEYINPUT84), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(KEYINPUT84), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n367), .B(new_n377), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382));
  INV_X1    g181(.A(G50gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(G22gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n330), .A2(new_n315), .A3(new_n331), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n244), .B1(new_n249), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n334), .B1(new_n251), .B2(new_n315), .ZN(new_n389));
  AND2_X1   g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  OR3_X1    g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT3), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n330), .A2(KEYINPUT81), .A3(new_n315), .A4(new_n331), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n244), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(G228gat), .B(G233gat), .C1(new_n395), .C2(new_n389), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n391), .B2(new_n396), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n401), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n391), .A2(new_n396), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT82), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n405), .B2(new_n398), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n386), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n401), .B1(new_n399), .B2(new_n400), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n398), .A3(new_n403), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n385), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n361), .A2(new_n381), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n313), .A2(new_n245), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n238), .A2(new_n295), .A3(new_n298), .A4(new_n312), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G227gat), .ZN(new_n417));
  INV_X1    g216(.A(G233gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT71), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT71), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n414), .A2(new_n422), .A3(new_n419), .A4(new_n415), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(new_n420), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT32), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT32), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n416), .B(new_n420), .C1(new_n422), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT34), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT72), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n430), .B1(new_n420), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT73), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n424), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G15gat), .B(G43gat), .Z(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT33), .B1(new_n421), .B2(new_n423), .ZN(new_n441));
  INV_X1    g240(.A(new_n439), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n441), .A2(new_n433), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n429), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n436), .A2(new_n434), .A3(new_n439), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n433), .B1(new_n441), .B2(new_n442), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n428), .A4(new_n426), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT36), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n367), .A2(new_n378), .ZN(new_n451));
  INV_X1    g250(.A(new_n342), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n450), .B1(new_n453), .B2(new_n411), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n451), .A2(new_n412), .A3(new_n452), .A4(new_n448), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n338), .A2(new_n341), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n407), .A2(new_n410), .A3(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n444), .A2(KEYINPUT85), .A3(new_n447), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT85), .B1(new_n444), .B2(new_n447), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n367), .B1(new_n379), .B2(new_n380), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n413), .A2(new_n454), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT12), .ZN(new_n466));
  XNOR2_X1  g265(.A(G113gat), .B(G141gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(G169gat), .B(G197gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  XOR2_X1   g268(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n469), .A2(new_n470), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(KEYINPUT12), .A3(new_n471), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n478), .B(KEYINPUT13), .Z(new_n479));
  NAND2_X1  g278(.A1(new_n383), .A2(G43gat), .ZN(new_n480));
  INV_X1    g279(.A(G43gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G50gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n482), .A3(KEYINPUT15), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G29gat), .ZN(new_n485));
  INV_X1    g284(.A(G36gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT14), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(G29gat), .B2(G36gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(G29gat), .A2(G36gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT89), .B1(new_n383), .B2(G43gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(new_n481), .A3(G50gat), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n383), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT15), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n483), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n492), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G1gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT16), .ZN(new_n506));
  INV_X1    g305(.A(G15gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G22gat), .ZN(new_n508));
  INV_X1    g307(.A(G22gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G15gat), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(G1gat), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g311(.A(G8gat), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n510), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n505), .ZN(new_n515));
  INV_X1    g314(.A(G8gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  INV_X1    g320(.A(new_n499), .ZN(new_n522));
  AOI21_X1  g321(.A(G50gat), .B1(new_n522), .B2(new_n497), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n493), .A2(new_n495), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n484), .A2(new_n491), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n527), .A2(new_n492), .B1(new_n513), .B2(new_n518), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n479), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n504), .A2(new_n519), .ZN(new_n530));
  OAI211_X1 g329(.A(KEYINPUT17), .B(new_n492), .C1(new_n501), .C2(new_n503), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n513), .A2(new_n518), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT17), .B1(new_n527), .B2(new_n492), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n478), .B(new_n530), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n477), .B(new_n529), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT92), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(KEYINPUT90), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n504), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(new_n532), .A3(new_n531), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n543), .A2(new_n544), .A3(new_n478), .A4(new_n530), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n536), .A3(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n538), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n539), .B1(new_n538), .B2(new_n546), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n529), .B1(new_n535), .B2(new_n536), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(new_n546), .B2(KEYINPUT91), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n540), .A2(new_n545), .A3(new_n552), .A4(new_n536), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n477), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n465), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n451), .ZN(new_n557));
  NAND2_X1  g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  OR2_X1    g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT9), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562));
  INV_X1    g361(.A(G57gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(G64gat), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(KEYINPUT93), .A3(G57gat), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n564), .B(new_n566), .C1(G57gat), .C2(new_n565), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n563), .A2(G64gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n565), .A2(G57gat), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT9), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n559), .A2(new_n558), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n561), .A2(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n573));
  AND2_X1   g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G127gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G183gat), .B(G211gat), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n575), .B(G127gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n519), .B1(KEYINPUT21), .B2(new_n572), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT94), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(new_n211), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n585), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n583), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT95), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n593));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n502), .A2(new_n483), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n598), .B1(new_n525), .B2(new_n526), .ZN(new_n599));
  OR2_X1    g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT97), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n603));
  AND2_X1   g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(G92gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n601), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(KEYINPUT96), .A2(G99gat), .A3(G106gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(KEYINPUT8), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n607), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT7), .ZN(new_n620));
  INV_X1    g419(.A(G85gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(G92gat), .A3(new_n610), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT8), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n601), .B2(new_n614), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n623), .A2(new_n609), .B1(new_n625), .B2(new_n616), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n602), .A2(new_n606), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n619), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n597), .B1(new_n599), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(KEYINPUT98), .B(new_n597), .C1(new_n599), .C2(new_n629), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT99), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n542), .A2(new_n531), .A3(new_n629), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n634), .B2(new_n638), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n596), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(new_n595), .A3(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n607), .B2(new_n618), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n607), .A2(new_n618), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n626), .A2(new_n627), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n648), .B(new_n572), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n567), .A2(new_n561), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n570), .A2(new_n571), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n628), .B(new_n619), .C1(new_n654), .C2(new_n647), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT10), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n629), .A2(new_n657), .A3(new_n654), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n646), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n651), .A2(new_n655), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n646), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT101), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n665), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n590), .A2(new_n645), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n556), .A2(new_n557), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n413), .A2(new_n454), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n456), .A2(new_n464), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n555), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n671), .A2(new_n452), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G8gat), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  NAND3_X1  g484(.A1(new_n556), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n676), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n676), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n675), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n689), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n691), .A2(new_n687), .A3(KEYINPUT102), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n690), .A2(new_n692), .ZN(G1325gat));
  NAND2_X1  g492(.A1(new_n556), .A2(new_n672), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n448), .B(KEYINPUT36), .ZN(new_n695));
  OAI21_X1  g494(.A(G15gat), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n460), .A2(new_n461), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n507), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n694), .B2(new_n698), .ZN(G1326gat));
  NOR2_X1   g498(.A1(new_n694), .A2(new_n412), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT43), .B(G22gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NOR3_X1   g501(.A1(new_n590), .A2(new_n645), .A3(new_n669), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n679), .A2(new_n680), .A3(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(G29gat), .A3(new_n451), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(KEYINPUT45), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n465), .B2(new_n645), .ZN(new_n709));
  INV_X1    g508(.A(new_n645), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n679), .A2(KEYINPUT44), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT103), .B1(new_n549), .B2(new_n554), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n546), .A2(KEYINPUT91), .ZN(new_n714));
  INV_X1    g513(.A(new_n550), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n553), .ZN(new_n716));
  INV_X1    g515(.A(new_n477), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n546), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT92), .B1(new_n719), .B2(new_n537), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n538), .A2(new_n539), .A3(new_n546), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n713), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n725), .A2(new_n590), .A3(new_n669), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n712), .A2(new_n557), .A3(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n706), .B(new_n707), .C1(new_n727), .C2(new_n485), .ZN(G1328gat));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n342), .A3(new_n726), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G36gat), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n452), .A2(G36gat), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT104), .B1(new_n704), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n556), .A2(new_n734), .A3(new_n703), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n736), .B2(KEYINPUT46), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739));
  AOI211_X1 g538(.A(KEYINPUT105), .B(new_n739), .C1(new_n733), .C2(new_n735), .ZN(new_n740));
  OAI221_X1 g539(.A(new_n730), .B1(KEYINPUT46), .B2(new_n736), .C1(new_n738), .C2(new_n740), .ZN(G1329gat));
  NOR2_X1   g540(.A1(new_n498), .A2(new_n499), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n695), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n712), .A2(new_n726), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n556), .A2(new_n697), .A3(new_n703), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n745), .A2(new_n742), .B1(new_n746), .B2(KEYINPUT47), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n746), .A2(KEYINPUT47), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1330gat));
  NAND4_X1  g549(.A1(new_n709), .A2(new_n711), .A3(new_n411), .A4(new_n726), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G50gat), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n556), .A2(new_n383), .A3(new_n411), .A4(new_n703), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1331gat));
  INV_X1    g555(.A(new_n725), .ZN(new_n757));
  NOR4_X1   g556(.A1(new_n757), .A2(new_n589), .A3(new_n710), .A4(new_n670), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n679), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n451), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(new_n563), .ZN(G1332gat));
  XNOR2_X1  g560(.A(new_n759), .B(KEYINPUT107), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n342), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT49), .B(G64gat), .Z(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n695), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n697), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n759), .B2(new_n770), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n769), .A2(KEYINPUT50), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT50), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n762), .A2(new_n411), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g575(.A1(new_n757), .A2(new_n590), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n342), .B1(new_n367), .B2(new_n378), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n695), .B1(new_n778), .B2(new_n412), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n411), .B1(new_n355), .B2(new_n360), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n381), .B2(new_n780), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n455), .A2(KEYINPUT35), .B1(new_n462), .B2(new_n463), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n710), .B(new_n777), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n679), .A2(KEYINPUT51), .A3(new_n710), .A4(new_n777), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n787), .A2(new_n621), .A3(new_n557), .A4(new_n669), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n757), .A2(new_n590), .A3(new_n670), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n709), .A2(new_n711), .A3(new_n557), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G85gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT108), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n788), .A2(new_n794), .A3(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1336gat));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n785), .A2(new_n797), .A3(new_n786), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT110), .A3(new_n784), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n452), .A2(G92gat), .A3(new_n670), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n709), .A2(new_n711), .A3(new_n342), .A4(new_n789), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(KEYINPUT109), .A3(G92gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT109), .B1(new_n802), .B2(G92gat), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT52), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(new_n802), .B2(G92gat), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n787), .A2(KEYINPUT111), .A3(new_n800), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT111), .B1(new_n787), .B2(new_n800), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n806), .A2(new_n810), .ZN(G1337gat));
  NAND3_X1  g610(.A1(new_n712), .A2(new_n450), .A3(new_n789), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G99gat), .ZN(new_n813));
  INV_X1    g612(.A(new_n787), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n770), .A2(G99gat), .A3(new_n670), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT112), .Z(new_n816));
  OAI21_X1  g615(.A(new_n813), .B1(new_n814), .B2(new_n816), .ZN(G1338gat));
  NOR3_X1   g616(.A1(new_n412), .A2(G106gat), .A3(new_n670), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n798), .A2(new_n799), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n709), .A2(new_n711), .A3(new_n411), .A4(new_n789), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT53), .B1(new_n787), .B2(new_n818), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n821), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1339gat));
  NOR2_X1   g625(.A1(new_n671), .A2(new_n757), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT113), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n478), .B1(new_n543), .B2(new_n530), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n520), .A2(new_n528), .A3(new_n479), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n475), .B(new_n471), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n547), .B2(new_n548), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n645), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n834), .B(new_n646), .C1(new_n656), .C2(new_n658), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n665), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(KEYINPUT114), .A3(new_n665), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n660), .A2(new_n657), .ZN(new_n841));
  INV_X1    g640(.A(new_n658), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n841), .A2(G230gat), .A3(G233gat), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(KEYINPUT54), .A3(new_n659), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n841), .A2(new_n842), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n834), .B1(new_n848), .B2(new_n646), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n849), .B2(new_n843), .ZN(new_n850));
  AOI211_X1 g649(.A(KEYINPUT115), .B(new_n666), .C1(new_n840), .C2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n835), .A2(KEYINPUT114), .A3(new_n665), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT114), .B1(new_n835), .B2(new_n665), .ZN(new_n854));
  OAI211_X1 g653(.A(KEYINPUT55), .B(new_n844), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n852), .B1(new_n855), .B2(new_n667), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n833), .B(new_n847), .C1(new_n851), .C2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n832), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n669), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n847), .B1(new_n851), .B2(new_n856), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n725), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n858), .B1(new_n862), .B2(new_n645), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n589), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI211_X1 g664(.A(KEYINPUT116), .B(new_n858), .C1(new_n645), .C2(new_n862), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n828), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(new_n557), .ZN(new_n868));
  INV_X1    g667(.A(new_n448), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n411), .A2(new_n869), .A3(new_n342), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(G113gat), .B1(new_n871), .B2(new_n757), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n412), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n557), .A2(new_n452), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n873), .A2(new_n770), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n680), .A2(G113gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(G1340gat));
  AOI21_X1  g676(.A(G120gat), .B1(new_n871), .B2(new_n669), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n669), .A2(G120gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n875), .B2(new_n879), .ZN(G1341gat));
  AND3_X1   g679(.A1(new_n868), .A2(new_n590), .A3(new_n870), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(G127gat), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n589), .A2(new_n576), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n883), .A2(new_n884), .B1(new_n875), .B2(new_n885), .ZN(G1342gat));
  INV_X1    g685(.A(G134gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n887), .A3(new_n710), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n875), .A2(new_n710), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n889), .B(new_n890), .C1(new_n887), .C2(new_n891), .ZN(G1343gat));
  NOR2_X1   g691(.A1(new_n874), .A2(new_n450), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT118), .Z(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n867), .B2(new_n411), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  INV_X1    g695(.A(new_n860), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n847), .A2(new_n667), .A3(new_n855), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n555), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n667), .A4(new_n855), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n857), .B1(new_n902), .B2(new_n710), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n589), .ZN(new_n904));
  AOI211_X1 g703(.A(new_n896), .B(new_n412), .C1(new_n904), .C2(new_n828), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n894), .B1(new_n895), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G141gat), .B1(new_n906), .B2(new_n555), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n450), .A2(new_n412), .A3(new_n342), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n868), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(G141gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(new_n680), .ZN(new_n911));
  XNOR2_X1  g710(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n907), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(G141gat), .B1(new_n906), .B2(new_n725), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(new_n911), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(G1344gat));
  OR3_X1    g716(.A1(new_n906), .A2(KEYINPUT59), .A3(new_n670), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n909), .B2(new_n669), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n671), .A2(new_n680), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n903), .B2(new_n589), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n411), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI211_X1 g723(.A(KEYINPUT121), .B(new_n921), .C1(new_n903), .C2(new_n589), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n896), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n867), .A2(KEYINPUT57), .A3(new_n411), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(new_n669), .A3(new_n894), .ZN(new_n929));
  NAND2_X1  g728(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n930));
  OAI221_X1 g729(.A(new_n918), .B1(new_n920), .B2(G148gat), .C1(new_n929), .C2(new_n930), .ZN(G1345gat));
  OAI21_X1  g730(.A(G155gat), .B1(new_n906), .B2(new_n589), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n909), .A2(new_n211), .A3(new_n590), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1346gat));
  OAI21_X1  g733(.A(G162gat), .B1(new_n906), .B2(new_n645), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n909), .A2(new_n212), .A3(new_n710), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1347gat));
  NOR3_X1   g736(.A1(new_n770), .A2(new_n557), .A3(new_n452), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n867), .A2(new_n412), .A3(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(new_n304), .A3(new_n555), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n867), .A2(new_n451), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n411), .A2(new_n869), .A3(new_n452), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n757), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n940), .B1(new_n945), .B2(new_n304), .ZN(G1348gat));
  OAI21_X1  g745(.A(G176gat), .B1(new_n939), .B2(new_n670), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n669), .A2(new_n305), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n943), .B2(new_n948), .ZN(G1349gat));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n867), .A2(new_n412), .A3(new_n590), .A4(new_n938), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G183gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n590), .A2(new_n299), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n867), .A2(new_n451), .A3(new_n942), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n952), .A2(KEYINPUT122), .A3(new_n955), .ZN(new_n959));
  AND4_X1   g758(.A1(new_n950), .A2(new_n958), .A3(KEYINPUT60), .A4(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT60), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n952), .A2(new_n961), .A3(new_n955), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT123), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n956), .B2(new_n957), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(new_n959), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n960), .A2(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n944), .A2(new_n296), .A3(new_n710), .ZN(new_n967));
  OAI21_X1  g766(.A(G190gat), .B1(new_n939), .B2(new_n645), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  NOR3_X1   g770(.A1(new_n450), .A2(new_n412), .A3(new_n452), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n941), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n757), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n557), .A2(new_n452), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n695), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n976), .B1(new_n926), .B2(new_n927), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n680), .A2(G197gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  INV_X1    g778(.A(new_n976), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n928), .A2(new_n669), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n977), .A2(new_n983), .A3(new_n669), .ZN(new_n984));
  XNOR2_X1  g783(.A(KEYINPUT124), .B(G204gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n987));
  AOI211_X1 g786(.A(new_n985), .B(new_n670), .C1(new_n987), .C2(KEYINPUT62), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n989), .B(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n986), .A2(new_n991), .ZN(G1353gat));
  INV_X1    g791(.A(KEYINPUT63), .ZN(new_n993));
  INV_X1    g792(.A(new_n977), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n993), .B(G211gat), .C1(new_n994), .C2(new_n589), .ZN(new_n995));
  AND4_X1   g794(.A1(new_n326), .A2(new_n941), .A3(new_n590), .A4(new_n972), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n996), .B(new_n997), .ZN(new_n998));
  AOI211_X1 g797(.A(new_n589), .B(new_n976), .C1(new_n926), .C2(new_n927), .ZN(new_n999));
  OAI21_X1  g798(.A(KEYINPUT63), .B1(new_n999), .B2(new_n326), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n995), .A2(new_n998), .A3(new_n1000), .ZN(G1354gat));
  OAI21_X1  g800(.A(G218gat), .B1(new_n994), .B2(new_n645), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n973), .A2(new_n327), .A3(new_n710), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1355gat));
endmodule


