

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801;

  INV_X1 U370 ( .A(KEYINPUT56), .ZN(n349) );
  INV_X1 U371 ( .A(KEYINPUT60), .ZN(n351) );
  XNOR2_X1 U372 ( .A(n702), .B(n701), .ZN(n703) );
  INV_X1 U373 ( .A(n384), .ZN(n353) );
  NOR2_X1 U374 ( .A1(n799), .A2(n604), .ZN(n605) );
  NAND2_X1 U375 ( .A1(n409), .A2(n429), .ZN(n801) );
  AND2_X1 U376 ( .A1(n433), .A2(n432), .ZN(n409) );
  AND2_X1 U377 ( .A1(n428), .A2(n451), .ZN(n435) );
  INV_X1 U378 ( .A(n572), .ZN(n355) );
  OR2_X1 U379 ( .A1(n730), .A2(n731), .ZN(n614) );
  XOR2_X1 U380 ( .A(KEYINPUT76), .B(KEYINPUT16), .Z(n529) );
  XNOR2_X1 U381 ( .A(n449), .B(n470), .ZN(n472) );
  XNOR2_X1 U382 ( .A(n438), .B(G131), .ZN(n437) );
  XNOR2_X1 U383 ( .A(G143), .B(G128), .ZN(n526) );
  XNOR2_X1 U384 ( .A(G104), .B(G107), .ZN(n509) );
  BUF_X4 U385 ( .A(n575), .Z(n583) );
  NOR2_X1 U386 ( .A1(n698), .A2(n679), .ZN(n680) );
  XNOR2_X1 U387 ( .A(n535), .B(n534), .ZN(n418) );
  XOR2_X2 U388 ( .A(KEYINPUT62), .B(n416), .Z(n675) );
  NOR2_X4 U389 ( .A1(n765), .A2(n763), .ZN(n732) );
  XNOR2_X2 U390 ( .A(KEYINPUT99), .B(n587), .ZN(n753) );
  XOR2_X2 U391 ( .A(n684), .B(KEYINPUT123), .Z(n685) );
  XNOR2_X1 U392 ( .A(n350), .B(n349), .ZN(G51) );
  NAND2_X1 U393 ( .A1(n671), .A2(n705), .ZN(n350) );
  XNOR2_X1 U394 ( .A(n352), .B(n351), .ZN(G60) );
  NAND2_X1 U395 ( .A1(n695), .A2(n705), .ZN(n352) );
  NAND2_X1 U396 ( .A1(n728), .A2(n727), .ZN(n612) );
  AND2_X2 U397 ( .A1(n354), .A2(n353), .ZN(n383) );
  NAND2_X1 U398 ( .A1(n400), .A2(n445), .ZN(n354) );
  NOR2_X2 U399 ( .A1(n753), .A2(n766), .ZN(n588) );
  AND2_X2 U400 ( .A1(n712), .A2(n713), .ZN(n592) );
  XNOR2_X2 U401 ( .A(n581), .B(n580), .ZN(n393) );
  XNOR2_X2 U402 ( .A(n356), .B(n355), .ZN(n602) );
  NOR2_X2 U403 ( .A1(n579), .A2(n448), .ZN(n356) );
  XNOR2_X1 U404 ( .A(G107), .B(G116), .ZN(n539) );
  BUF_X1 U405 ( .A(G113), .Z(n404) );
  XOR2_X1 U406 ( .A(n556), .B(n555), .Z(n357) );
  XOR2_X1 U407 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n358) );
  OR2_X1 U408 ( .A1(G953), .A2(G237), .ZN(n359) );
  NAND2_X1 U409 ( .A1(n662), .A2(n709), .ZN(n689) );
  BUF_X1 U410 ( .A(n660), .Z(n778) );
  NOR2_X1 U411 ( .A1(n602), .A2(n413), .ZN(n406) );
  NOR2_X1 U412 ( .A1(n616), .A2(n716), .ZN(n713) );
  XNOR2_X1 U413 ( .A(n634), .B(n563), .ZN(n624) );
  NAND2_X1 U414 ( .A1(n375), .A2(n373), .ZN(n616) );
  NAND2_X1 U415 ( .A1(n381), .A2(n727), .ZN(n634) );
  INV_X2 U416 ( .A(G953), .ZN(n791) );
  OR2_X2 U417 ( .A1(n689), .A2(n673), .ZN(n676) );
  NOR2_X1 U418 ( .A1(n624), .A2(n566), .ZN(n569) );
  NAND2_X1 U419 ( .A1(n387), .A2(n398), .ZN(n384) );
  OR2_X1 U420 ( .A1(n626), .A2(n372), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n569), .B(n568), .ZN(n579) );
  NAND2_X1 U422 ( .A1(n360), .A2(n616), .ZN(n403) );
  XNOR2_X1 U423 ( .A(n419), .B(n412), .ZN(n455) );
  XNOR2_X1 U424 ( .A(n511), .B(n510), .ZN(n771) );
  INV_X1 U425 ( .A(KEYINPUT44), .ZN(n402) );
  INV_X1 U426 ( .A(KEYINPUT10), .ZN(n379) );
  INV_X1 U427 ( .A(G125), .ZN(n380) );
  INV_X1 U428 ( .A(KEYINPUT105), .ZN(n405) );
  BUF_X2 U429 ( .A(n689), .Z(n698) );
  AND2_X2 U430 ( .A1(n383), .A2(n382), .ZN(n789) );
  NAND2_X1 U431 ( .A1(n386), .A2(n385), .ZN(n382) );
  AND2_X1 U432 ( .A1(n778), .A2(KEYINPUT2), .ZN(n661) );
  NAND2_X1 U433 ( .A1(n399), .A2(n445), .ZN(n387) );
  XNOR2_X1 U434 ( .A(n610), .B(KEYINPUT45), .ZN(n660) );
  AND2_X1 U435 ( .A1(n748), .A2(n743), .ZN(n388) );
  INV_X1 U436 ( .A(n444), .ZN(n396) );
  NOR2_X1 U437 ( .A1(n391), .A2(n390), .ZN(n389) );
  NAND2_X1 U438 ( .A1(n436), .A2(n450), .ZN(n434) );
  NOR2_X1 U439 ( .A1(n796), .A2(n423), .ZN(n589) );
  AND2_X1 U440 ( .A1(n637), .A2(n371), .ZN(n370) );
  XNOR2_X1 U441 ( .A(n406), .B(n405), .ZN(n796) );
  INV_X1 U442 ( .A(n392), .ZN(n723) );
  INV_X1 U443 ( .A(n743), .ZN(n390) );
  NAND2_X1 U444 ( .A1(n369), .A2(n627), .ZN(n368) );
  XNOR2_X1 U445 ( .A(n594), .B(n593), .ZN(n736) );
  NAND2_X1 U446 ( .A1(n462), .A2(n586), .ZN(n587) );
  AND2_X1 U447 ( .A1(n626), .A2(n372), .ZN(n371) );
  AND2_X1 U448 ( .A1(n632), .A2(n633), .ZN(n361) );
  NAND2_X1 U449 ( .A1(n616), .A2(n615), .ZN(n629) );
  INV_X1 U450 ( .A(n417), .ZN(n360) );
  AND2_X1 U451 ( .A1(n591), .A2(n578), .ZN(n763) );
  NOR2_X1 U452 ( .A1(n591), .A2(n590), .ZN(n640) );
  AND2_X1 U453 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U454 ( .A1(n499), .A2(n550), .ZN(n374) );
  NAND2_X1 U455 ( .A1(n378), .A2(G902), .ZN(n376) );
  OR2_X1 U456 ( .A1(G902), .A2(n692), .ZN(n561) );
  NAND2_X1 U457 ( .A1(n702), .A2(n550), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n455), .B(n454), .ZN(n664) );
  XNOR2_X1 U459 ( .A(n362), .B(n557), .ZN(n559) );
  XNOR2_X1 U460 ( .A(n771), .B(KEYINPUT73), .ZN(n525) );
  XNOR2_X1 U461 ( .A(n357), .B(n558), .ZN(n362) );
  XNOR2_X1 U462 ( .A(n523), .B(n379), .ZN(n558) );
  XNOR2_X1 U463 ( .A(n482), .B(KEYINPUT30), .ZN(n483) );
  XNOR2_X1 U464 ( .A(n380), .B(G146), .ZN(n523) );
  XNOR2_X1 U465 ( .A(n567), .B(KEYINPUT0), .ZN(n568) );
  XNOR2_X1 U466 ( .A(G104), .B(n404), .ZN(n553) );
  INV_X1 U467 ( .A(n582), .ZN(n364) );
  NOR2_X1 U468 ( .A1(n466), .A2(G953), .ZN(n465) );
  OR2_X1 U469 ( .A1(n791), .A2(G952), .ZN(n705) );
  INV_X1 U470 ( .A(KEYINPUT24), .ZN(n488) );
  XNOR2_X1 U471 ( .A(G119), .B(G128), .ZN(n486) );
  NAND2_X1 U472 ( .A1(G234), .A2(G237), .ZN(n502) );
  INV_X1 U473 ( .A(G237), .ZN(n480) );
  INV_X1 U474 ( .A(KEYINPUT72), .ZN(n470) );
  XNOR2_X1 U475 ( .A(KEYINPUT74), .B(G472), .ZN(n479) );
  XOR2_X1 U476 ( .A(KEYINPUT3), .B(G119), .Z(n471) );
  XNOR2_X1 U477 ( .A(G110), .B(G137), .ZN(n489) );
  XNOR2_X1 U478 ( .A(G101), .B(G110), .ZN(n511) );
  NAND2_X1 U479 ( .A1(n393), .A2(n462), .ZN(n365) );
  NAND2_X1 U480 ( .A1(n442), .A2(n440), .ZN(n400) );
  NAND2_X1 U481 ( .A1(n446), .A2(KEYINPUT87), .ZN(n395) );
  NAND2_X1 U482 ( .A1(n631), .A2(n361), .ZN(n646) );
  NAND2_X1 U483 ( .A1(n363), .A2(n650), .ZN(n651) );
  XNOR2_X1 U484 ( .A(n649), .B(n358), .ZN(n363) );
  XNOR2_X2 U485 ( .A(n365), .B(n364), .ZN(n766) );
  XNOR2_X2 U486 ( .A(n583), .B(n576), .ZN(n632) );
  NAND2_X1 U487 ( .A1(n367), .A2(n366), .ZN(n427) );
  OR2_X1 U488 ( .A1(n637), .A2(n372), .ZN(n366) );
  NOR2_X1 U489 ( .A1(n370), .A2(n368), .ZN(n367) );
  INV_X1 U490 ( .A(KEYINPUT47), .ZN(n372) );
  OR2_X1 U491 ( .A1(n681), .A2(n374), .ZN(n373) );
  NAND2_X1 U492 ( .A1(n681), .A2(n378), .ZN(n377) );
  INV_X1 U493 ( .A(n629), .ZN(n617) );
  INV_X1 U494 ( .A(n499), .ZN(n378) );
  XNOR2_X1 U495 ( .A(n535), .B(n534), .ZN(n381) );
  INV_X1 U496 ( .A(n400), .ZN(n385) );
  NOR2_X1 U497 ( .A1(n396), .A2(n395), .ZN(n386) );
  NAND2_X1 U498 ( .A1(n464), .A2(n388), .ZN(n749) );
  NAND2_X1 U499 ( .A1(n464), .A2(n389), .ZN(n421) );
  INV_X1 U500 ( .A(n741), .ZN(n391) );
  OR2_X1 U501 ( .A1(n722), .A2(n393), .ZN(n392) );
  XNOR2_X1 U502 ( .A(n620), .B(KEYINPUT1), .ZN(n712) );
  XNOR2_X2 U503 ( .A(n394), .B(n517), .ZN(n620) );
  XNOR2_X2 U504 ( .A(n516), .B(n515), .ZN(n702) );
  NAND2_X1 U505 ( .A1(n444), .A2(n446), .ZN(n399) );
  INV_X1 U506 ( .A(n800), .ZN(n398) );
  OR2_X2 U507 ( .A1(n401), .A2(n481), .ZN(n484) );
  NOR2_X1 U508 ( .A1(n401), .A2(n618), .ZN(n619) );
  AND2_X1 U509 ( .A1(n401), .A2(n573), .ZN(n604) );
  XNOR2_X2 U510 ( .A(n575), .B(KEYINPUT107), .ZN(n401) );
  XNOR2_X1 U511 ( .A(n605), .B(n402), .ZN(n607) );
  NOR2_X1 U512 ( .A1(n602), .A2(n403), .ZN(n573) );
  BUF_X1 U513 ( .A(n530), .Z(n407) );
  XNOR2_X1 U514 ( .A(n461), .B(n595), .ZN(n460) );
  INV_X1 U515 ( .A(n579), .ZN(n462) );
  XNOR2_X1 U516 ( .A(G902), .B(KEYINPUT15), .ZN(n496) );
  INV_X1 U517 ( .A(n795), .ZN(n446) );
  XNOR2_X1 U518 ( .A(n467), .B(n465), .ZN(n527) );
  XNOR2_X1 U519 ( .A(n526), .B(KEYINPUT18), .ZN(n456) );
  XNOR2_X1 U520 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n467) );
  NOR2_X1 U521 ( .A1(n625), .A2(KEYINPUT42), .ZN(n430) );
  NAND2_X1 U522 ( .A1(n630), .A2(KEYINPUT40), .ZN(n451) );
  INV_X1 U523 ( .A(KEYINPUT100), .ZN(n580) );
  XNOR2_X1 U524 ( .A(n425), .B(n424), .ZN(n499) );
  XNOR2_X1 U525 ( .A(n498), .B(KEYINPUT80), .ZN(n424) );
  XNOR2_X1 U526 ( .A(n571), .B(KEYINPUT22), .ZN(n572) );
  INV_X1 U527 ( .A(KEYINPUT75), .ZN(n571) );
  AND2_X1 U528 ( .A1(n426), .A2(n408), .ZN(n643) );
  NAND2_X1 U529 ( .A1(n427), .A2(n410), .ZN(n426) );
  INV_X1 U530 ( .A(G224), .ZN(n466) );
  XNOR2_X1 U531 ( .A(n497), .B(KEYINPUT20), .ZN(n500) );
  XNOR2_X1 U532 ( .A(KEYINPUT5), .B(G101), .ZN(n474) );
  INV_X1 U533 ( .A(n496), .ZN(n657) );
  XNOR2_X1 U534 ( .A(n533), .B(n532), .ZN(n534) );
  INV_X1 U535 ( .A(G902), .ZN(n550) );
  NAND2_X1 U536 ( .A1(n500), .A2(G217), .ZN(n425) );
  NAND2_X1 U537 ( .A1(n570), .A2(n615), .ZN(n448) );
  INV_X1 U538 ( .A(KEYINPUT87), .ZN(n445) );
  INV_X1 U539 ( .A(G134), .ZN(n468) );
  XNOR2_X1 U540 ( .A(n525), .B(n457), .ZN(n454) );
  XNOR2_X1 U541 ( .A(n458), .B(n524), .ZN(n457) );
  NAND2_X1 U542 ( .A1(n463), .A2(n462), .ZN(n461) );
  INV_X1 U543 ( .A(n736), .ZN(n463) );
  NAND2_X1 U544 ( .A1(n431), .A2(n430), .ZN(n429) );
  NOR2_X1 U545 ( .A1(n630), .A2(KEYINPUT40), .ZN(n450) );
  XNOR2_X1 U546 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n582) );
  NOR2_X1 U547 ( .A1(n639), .A2(n759), .ZN(n408) );
  OR2_X1 U548 ( .A1(n628), .A2(n627), .ZN(n410) );
  XOR2_X1 U549 ( .A(n529), .B(G122), .Z(n411) );
  XOR2_X1 U550 ( .A(n527), .B(n456), .Z(n412) );
  NAND2_X1 U551 ( .A1(n577), .A2(n360), .ZN(n413) );
  AND2_X1 U552 ( .A1(n420), .A2(n742), .ZN(n414) );
  BUF_X1 U553 ( .A(n674), .Z(n416) );
  BUF_X1 U554 ( .A(n712), .Z(n417) );
  XNOR2_X1 U555 ( .A(n419), .B(n771), .ZN(n772) );
  XNOR2_X2 U556 ( .A(n530), .B(n411), .ZN(n419) );
  NAND2_X1 U557 ( .A1(n421), .A2(n414), .ZN(n422) );
  NAND2_X1 U558 ( .A1(n741), .A2(G953), .ZN(n420) );
  NAND2_X1 U559 ( .A1(n422), .A2(n749), .ZN(n751) );
  NOR2_X1 U560 ( .A1(n588), .A2(n732), .ZN(n423) );
  NAND2_X1 U561 ( .A1(n653), .A2(KEYINPUT40), .ZN(n428) );
  NAND2_X2 U562 ( .A1(n622), .A2(n801), .ZN(n452) );
  INV_X1 U563 ( .A(n724), .ZN(n431) );
  NAND2_X1 U564 ( .A1(n625), .A2(KEYINPUT42), .ZN(n432) );
  NAND2_X1 U565 ( .A1(n724), .A2(KEYINPUT42), .ZN(n433) );
  NAND2_X2 U566 ( .A1(n435), .A2(n434), .ZN(n622) );
  XNOR2_X2 U567 ( .A(n614), .B(n613), .ZN(n724) );
  INV_X1 U568 ( .A(n653), .ZN(n436) );
  XNOR2_X2 U569 ( .A(n528), .B(n437), .ZN(n469) );
  XNOR2_X2 U570 ( .A(KEYINPUT69), .B(G137), .ZN(n438) );
  XNOR2_X2 U571 ( .A(n439), .B(KEYINPUT4), .ZN(n528) );
  XNOR2_X2 U572 ( .A(KEYINPUT64), .B(KEYINPUT67), .ZN(n439) );
  NAND2_X1 U573 ( .A1(n644), .A2(n441), .ZN(n440) );
  AND2_X1 U574 ( .A1(n643), .A2(n447), .ZN(n441) );
  NAND2_X1 U575 ( .A1(n443), .A2(n645), .ZN(n442) );
  INV_X1 U576 ( .A(n644), .ZN(n443) );
  OR2_X1 U577 ( .A1(n643), .A2(n447), .ZN(n444) );
  INV_X1 U578 ( .A(n645), .ZN(n447) );
  XNOR2_X2 U579 ( .A(G116), .B(G113), .ZN(n449) );
  XNOR2_X2 U580 ( .A(n452), .B(n623), .ZN(n644) );
  XNOR2_X2 U581 ( .A(n453), .B(n479), .ZN(n575) );
  OR2_X2 U582 ( .A1(n674), .A2(G902), .ZN(n453) );
  XNOR2_X2 U583 ( .A(n472), .B(n471), .ZN(n530) );
  INV_X1 U584 ( .A(n528), .ZN(n458) );
  XNOR2_X2 U585 ( .A(n459), .B(KEYINPUT35), .ZN(n797) );
  NAND2_X1 U586 ( .A1(n460), .A2(n640), .ZN(n459) );
  XNOR2_X1 U587 ( .A(n711), .B(KEYINPUT86), .ZN(n464) );
  OR2_X2 U588 ( .A1(n698), .A2(n697), .ZN(n704) );
  OR2_X2 U589 ( .A1(n698), .A2(n683), .ZN(n686) );
  XNOR2_X2 U590 ( .A(n785), .B(G146), .ZN(n516) );
  XNOR2_X2 U591 ( .A(n469), .B(n547), .ZN(n785) );
  INV_X1 U592 ( .A(n523), .ZN(n524) );
  INV_X1 U593 ( .A(KEYINPUT93), .ZN(n532) );
  XNOR2_X1 U594 ( .A(n489), .B(n488), .ZN(n490) );
  INV_X1 U595 ( .A(KEYINPUT34), .ZN(n595) );
  XNOR2_X1 U596 ( .A(n491), .B(n490), .ZN(n494) );
  XNOR2_X1 U597 ( .A(n526), .B(n468), .ZN(n547) );
  XNOR2_X1 U598 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n473) );
  XNOR2_X1 U599 ( .A(n474), .B(n473), .ZN(n476) );
  XNOR2_X1 U600 ( .A(KEYINPUT77), .B(n359), .ZN(n552) );
  NAND2_X1 U601 ( .A1(n552), .A2(G210), .ZN(n475) );
  XNOR2_X1 U602 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U603 ( .A(n407), .B(n477), .ZN(n478) );
  XNOR2_X1 U604 ( .A(n516), .B(n478), .ZN(n674) );
  NAND2_X1 U605 ( .A1(n550), .A2(n480), .ZN(n531) );
  NAND2_X1 U606 ( .A1(n531), .A2(G214), .ZN(n727) );
  INV_X1 U607 ( .A(n727), .ZN(n481) );
  INV_X1 U608 ( .A(KEYINPUT110), .ZN(n482) );
  XNOR2_X1 U609 ( .A(n484), .B(n483), .ZN(n520) );
  XOR2_X1 U610 ( .A(G140), .B(KEYINPUT68), .Z(n513) );
  INV_X1 U611 ( .A(n513), .ZN(n485) );
  XNOR2_X1 U612 ( .A(n558), .B(n485), .ZN(n783) );
  XOR2_X1 U613 ( .A(KEYINPUT84), .B(KEYINPUT23), .Z(n487) );
  XNOR2_X1 U614 ( .A(n487), .B(n486), .ZN(n491) );
  NAND2_X1 U615 ( .A1(G234), .A2(n791), .ZN(n492) );
  XOR2_X1 U616 ( .A(KEYINPUT8), .B(n492), .Z(n545) );
  NAND2_X1 U617 ( .A1(n545), .A2(G221), .ZN(n493) );
  XNOR2_X1 U618 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U619 ( .A(n783), .B(n495), .ZN(n681) );
  XOR2_X1 U620 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n498) );
  NAND2_X1 U621 ( .A1(n496), .A2(G234), .ZN(n497) );
  NAND2_X1 U622 ( .A1(G221), .A2(n500), .ZN(n501) );
  XOR2_X1 U623 ( .A(KEYINPUT21), .B(n501), .Z(n615) );
  INV_X1 U624 ( .A(n615), .ZN(n716) );
  XNOR2_X1 U625 ( .A(n502), .B(KEYINPUT94), .ZN(n503) );
  XNOR2_X1 U626 ( .A(KEYINPUT14), .B(n503), .ZN(n505) );
  NAND2_X1 U627 ( .A1(n505), .A2(G902), .ZN(n564) );
  OR2_X1 U628 ( .A1(n791), .A2(n564), .ZN(n504) );
  NOR2_X1 U629 ( .A1(G900), .A2(n504), .ZN(n506) );
  AND2_X1 U630 ( .A1(n505), .A2(G952), .ZN(n744) );
  AND2_X1 U631 ( .A1(n744), .A2(n791), .ZN(n740) );
  NOR2_X1 U632 ( .A1(n506), .A2(n740), .ZN(n508) );
  INV_X1 U633 ( .A(KEYINPUT82), .ZN(n507) );
  XNOR2_X1 U634 ( .A(n508), .B(n507), .ZN(n633) );
  NAND2_X1 U635 ( .A1(n713), .A2(n633), .ZN(n518) );
  INV_X1 U636 ( .A(n509), .ZN(n510) );
  NAND2_X1 U637 ( .A1(G227), .A2(n791), .ZN(n512) );
  XNOR2_X1 U638 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U639 ( .A(n525), .B(n514), .ZN(n515) );
  XOR2_X1 U640 ( .A(KEYINPUT71), .B(G469), .Z(n517) );
  INV_X1 U641 ( .A(n620), .ZN(n584) );
  NOR2_X1 U642 ( .A1(n518), .A2(n584), .ZN(n519) );
  NAND2_X1 U643 ( .A1(n520), .A2(n519), .ZN(n522) );
  INV_X1 U644 ( .A(KEYINPUT78), .ZN(n521) );
  XNOR2_X1 U645 ( .A(n522), .B(n521), .ZN(n642) );
  NOR2_X2 U646 ( .A1(n664), .A2(n657), .ZN(n535) );
  NAND2_X1 U647 ( .A1(G210), .A2(n531), .ZN(n533) );
  INV_X1 U648 ( .A(KEYINPUT38), .ZN(n536) );
  XNOR2_X1 U649 ( .A(n418), .B(n536), .ZN(n728) );
  NAND2_X1 U650 ( .A1(n642), .A2(n728), .ZN(n538) );
  INV_X1 U651 ( .A(KEYINPUT39), .ZN(n537) );
  XNOR2_X2 U652 ( .A(n538), .B(n537), .ZN(n653) );
  XOR2_X1 U653 ( .A(KEYINPUT102), .B(G122), .Z(n540) );
  XNOR2_X1 U654 ( .A(n540), .B(n539), .ZN(n544) );
  XOR2_X1 U655 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n542) );
  XNOR2_X1 U656 ( .A(KEYINPUT9), .B(KEYINPUT104), .ZN(n541) );
  XNOR2_X1 U657 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U658 ( .A(n544), .B(n543), .Z(n549) );
  NAND2_X1 U659 ( .A1(G217), .A2(n545), .ZN(n546) );
  XNOR2_X1 U660 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U661 ( .A(n549), .B(n548), .ZN(n684) );
  NAND2_X1 U662 ( .A1(n684), .A2(n550), .ZN(n551) );
  INV_X1 U663 ( .A(G478), .ZN(n683) );
  XNOR2_X1 U664 ( .A(n551), .B(n683), .ZN(n591) );
  XNOR2_X1 U665 ( .A(KEYINPUT13), .B(G475), .ZN(n562) );
  NAND2_X1 U666 ( .A1(n552), .A2(G214), .ZN(n560) );
  XOR2_X1 U667 ( .A(G143), .B(G122), .Z(n554) );
  XNOR2_X1 U668 ( .A(n554), .B(n553), .ZN(n557) );
  XOR2_X1 U669 ( .A(G131), .B(KEYINPUT11), .Z(n556) );
  XNOR2_X1 U670 ( .A(G140), .B(KEYINPUT12), .ZN(n555) );
  XNOR2_X1 U671 ( .A(n560), .B(n559), .ZN(n692) );
  XNOR2_X1 U672 ( .A(n562), .B(n561), .ZN(n590) );
  INV_X1 U673 ( .A(n590), .ZN(n578) );
  INV_X1 U674 ( .A(n763), .ZN(n630) );
  XNOR2_X1 U675 ( .A(n622), .B(G131), .ZN(G33) );
  XNOR2_X1 U676 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n563) );
  XNOR2_X1 U677 ( .A(G898), .B(KEYINPUT95), .ZN(n777) );
  NAND2_X1 U678 ( .A1(G953), .A2(n777), .ZN(n773) );
  NOR2_X1 U679 ( .A1(n564), .A2(n773), .ZN(n565) );
  NOR2_X1 U680 ( .A1(n740), .A2(n565), .ZN(n566) );
  INV_X1 U681 ( .A(KEYINPUT66), .ZN(n567) );
  NAND2_X1 U682 ( .A1(n590), .A2(n591), .ZN(n730) );
  INV_X1 U683 ( .A(n730), .ZN(n570) );
  INV_X1 U684 ( .A(n604), .ZN(n574) );
  XNOR2_X1 U685 ( .A(n574), .B(G110), .ZN(G12) );
  INV_X1 U686 ( .A(KEYINPUT6), .ZN(n576) );
  NOR2_X1 U687 ( .A1(n632), .A2(n616), .ZN(n577) );
  OR2_X1 U688 ( .A1(n591), .A2(n578), .ZN(n652) );
  INV_X1 U689 ( .A(n652), .ZN(n765) );
  NAND2_X1 U690 ( .A1(n592), .A2(n583), .ZN(n581) );
  INV_X1 U691 ( .A(n583), .ZN(n718) );
  NAND2_X1 U692 ( .A1(n713), .A2(n718), .ZN(n585) );
  NOR2_X1 U693 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U694 ( .A(n589), .B(KEYINPUT106), .ZN(n597) );
  NAND2_X1 U695 ( .A1(n592), .A2(n632), .ZN(n594) );
  INV_X1 U696 ( .A(KEYINPUT33), .ZN(n593) );
  NAND2_X1 U697 ( .A1(n797), .A2(KEYINPUT44), .ZN(n596) );
  NAND2_X1 U698 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U699 ( .A(n598), .B(KEYINPUT89), .ZN(n609) );
  NAND2_X1 U700 ( .A1(n616), .A2(n417), .ZN(n599) );
  NOR2_X1 U701 ( .A1(n632), .A2(n599), .ZN(n600) );
  XNOR2_X1 U702 ( .A(n600), .B(KEYINPUT81), .ZN(n601) );
  NOR2_X1 U703 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U704 ( .A(KEYINPUT32), .B(n603), .ZN(n799) );
  NAND2_X1 U705 ( .A1(n605), .A2(n797), .ZN(n606) );
  NAND2_X1 U706 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U707 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U708 ( .A1(n660), .A2(n657), .ZN(n611) );
  XNOR2_X1 U709 ( .A(n611), .B(KEYINPUT85), .ZN(n656) );
  XOR2_X1 U710 ( .A(n612), .B(KEYINPUT111), .Z(n731) );
  INV_X1 U711 ( .A(KEYINPUT41), .ZN(n613) );
  NAND2_X1 U712 ( .A1(n633), .A2(n617), .ZN(n618) );
  XNOR2_X1 U713 ( .A(KEYINPUT28), .B(n619), .ZN(n621) );
  NAND2_X1 U714 ( .A1(n621), .A2(n620), .ZN(n625) );
  XOR2_X1 U715 ( .A(KEYINPUT88), .B(KEYINPUT46), .Z(n623) );
  NOR2_X1 U716 ( .A1(n625), .A2(n624), .ZN(n637) );
  INV_X1 U717 ( .A(n732), .ZN(n626) );
  NAND2_X1 U718 ( .A1(KEYINPUT47), .A2(n626), .ZN(n628) );
  INV_X1 U719 ( .A(KEYINPUT83), .ZN(n627) );
  NOR2_X1 U720 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U721 ( .A1(n646), .A2(n634), .ZN(n635) );
  XNOR2_X1 U722 ( .A(n635), .B(KEYINPUT36), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n636), .A2(n417), .ZN(n768) );
  NAND2_X1 U724 ( .A1(n637), .A2(KEYINPUT83), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n768), .A2(n638), .ZN(n639) );
  AND2_X1 U726 ( .A1(n418), .A2(n640), .ZN(n641) );
  AND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n759) );
  XNOR2_X1 U728 ( .A(KEYINPUT70), .B(KEYINPUT48), .ZN(n645) );
  INV_X1 U729 ( .A(n646), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n647), .A2(n727), .ZN(n648) );
  NOR2_X1 U731 ( .A1(n417), .A2(n648), .ZN(n649) );
  INV_X1 U732 ( .A(n418), .ZN(n650) );
  XNOR2_X1 U733 ( .A(n651), .B(KEYINPUT109), .ZN(n795) );
  OR2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n655) );
  INV_X1 U735 ( .A(KEYINPUT112), .ZN(n654) );
  XNOR2_X1 U736 ( .A(n655), .B(n654), .ZN(n800) );
  NAND2_X1 U737 ( .A1(n656), .A2(n789), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n657), .A2(KEYINPUT2), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n661), .A2(n789), .ZN(n709) );
  INV_X1 U741 ( .A(G210), .ZN(n663) );
  NOR2_X1 U742 ( .A1(n689), .A2(n663), .ZN(n670) );
  BUF_X1 U743 ( .A(n664), .Z(n668) );
  XOR2_X1 U744 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n666) );
  XNOR2_X1 U745 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n665) );
  XOR2_X1 U746 ( .A(n666), .B(n665), .Z(n667) );
  XNOR2_X1 U747 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U748 ( .A(n670), .B(n669), .ZN(n671) );
  INV_X1 U749 ( .A(G472), .ZN(n673) );
  XNOR2_X1 U750 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U751 ( .A1(n677), .A2(n705), .ZN(n678) );
  XNOR2_X1 U752 ( .A(n678), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U753 ( .A(G217), .ZN(n679) );
  XNOR2_X1 U754 ( .A(n681), .B(n680), .ZN(n682) );
  AND2_X1 U755 ( .A1(n682), .A2(n705), .ZN(G66) );
  XNOR2_X1 U756 ( .A(n686), .B(n685), .ZN(n687) );
  AND2_X1 U757 ( .A1(n687), .A2(n705), .ZN(G63) );
  INV_X1 U758 ( .A(G475), .ZN(n688) );
  NOR2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n694) );
  XNOR2_X1 U760 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n690) );
  XOR2_X1 U761 ( .A(n690), .B(KEYINPUT65), .Z(n691) );
  XOR2_X1 U762 ( .A(n692), .B(n691), .Z(n693) );
  XNOR2_X1 U763 ( .A(n694), .B(n693), .ZN(n695) );
  INV_X1 U764 ( .A(G469), .ZN(n697) );
  XOR2_X1 U765 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n700) );
  XNOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n699) );
  XOR2_X1 U767 ( .A(n700), .B(n699), .Z(n701) );
  XNOR2_X1 U768 ( .A(n704), .B(n703), .ZN(n706) );
  AND2_X1 U769 ( .A1(n706), .A2(n705), .ZN(G54) );
  NAND2_X1 U770 ( .A1(n778), .A2(n789), .ZN(n708) );
  INV_X1 U771 ( .A(KEYINPUT2), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  OR2_X1 U774 ( .A1(n724), .A2(n736), .ZN(n743) );
  NOR2_X1 U775 ( .A1(n713), .A2(n417), .ZN(n715) );
  XNOR2_X1 U776 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n714) );
  XNOR2_X1 U777 ( .A(n715), .B(n714), .ZN(n721) );
  NAND2_X1 U778 ( .A1(n616), .A2(n716), .ZN(n717) );
  XOR2_X1 U779 ( .A(KEYINPUT49), .B(n717), .Z(n719) );
  NAND2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U781 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U782 ( .A(KEYINPUT51), .B(n723), .ZN(n725) );
  NAND2_X1 U783 ( .A1(n725), .A2(n431), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n726), .B(KEYINPUT117), .ZN(n738) );
  NOR2_X1 U785 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U786 ( .A1(n730), .A2(n729), .ZN(n734) );
  NOR2_X1 U787 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U788 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U790 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U791 ( .A(KEYINPUT52), .B(n739), .Z(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(n740), .ZN(n741) );
  INV_X1 U793 ( .A(KEYINPUT118), .ZN(n742) );
  AND2_X1 U794 ( .A1(n745), .A2(n744), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n791), .A2(KEYINPUT118), .ZN(n746) );
  NOR2_X1 U796 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U797 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n750) );
  XNOR2_X1 U798 ( .A(n751), .B(n750), .ZN(G75) );
  NAND2_X1 U799 ( .A1(n753), .A2(n763), .ZN(n752) );
  XNOR2_X1 U800 ( .A(n752), .B(G104), .ZN(G6) );
  XOR2_X1 U801 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n755) );
  NAND2_X1 U802 ( .A1(n753), .A2(n765), .ZN(n754) );
  XNOR2_X1 U803 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U804 ( .A(G107), .B(n756), .ZN(G9) );
  XOR2_X1 U805 ( .A(G128), .B(KEYINPUT29), .Z(n758) );
  NAND2_X1 U806 ( .A1(n637), .A2(n765), .ZN(n757) );
  XNOR2_X1 U807 ( .A(n758), .B(n757), .ZN(G30) );
  XNOR2_X1 U808 ( .A(G143), .B(n759), .ZN(n760) );
  XNOR2_X1 U809 ( .A(n760), .B(KEYINPUT113), .ZN(G45) );
  NAND2_X1 U810 ( .A1(n637), .A2(n763), .ZN(n761) );
  XNOR2_X1 U811 ( .A(n761), .B(KEYINPUT114), .ZN(n762) );
  XNOR2_X1 U812 ( .A(G146), .B(n762), .ZN(G48) );
  NAND2_X1 U813 ( .A1(n766), .A2(n763), .ZN(n764) );
  XNOR2_X1 U814 ( .A(n404), .B(n764), .ZN(G15) );
  NAND2_X1 U815 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U816 ( .A(n767), .B(G116), .ZN(G18) );
  XNOR2_X1 U817 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n769) );
  XNOR2_X1 U818 ( .A(n769), .B(n768), .ZN(n770) );
  XNOR2_X1 U819 ( .A(G125), .B(n770), .ZN(G27) );
  XNOR2_X1 U820 ( .A(KEYINPUT124), .B(n772), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n774), .A2(n773), .ZN(n782) );
  NAND2_X1 U822 ( .A1(G953), .A2(G224), .ZN(n775) );
  XOR2_X1 U823 ( .A(KEYINPUT61), .B(n775), .Z(n776) );
  NOR2_X1 U824 ( .A1(n777), .A2(n776), .ZN(n780) );
  AND2_X1 U825 ( .A1(n778), .A2(n791), .ZN(n779) );
  NOR2_X1 U826 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U827 ( .A(n782), .B(n781), .ZN(G69) );
  XNOR2_X1 U828 ( .A(n783), .B(KEYINPUT125), .ZN(n784) );
  XNOR2_X1 U829 ( .A(n785), .B(n784), .ZN(n790) );
  XOR2_X1 U830 ( .A(G227), .B(n790), .Z(n786) );
  NAND2_X1 U831 ( .A1(n786), .A2(G900), .ZN(n787) );
  NAND2_X1 U832 ( .A1(n787), .A2(G953), .ZN(n788) );
  XNOR2_X1 U833 ( .A(n788), .B(KEYINPUT126), .ZN(n794) );
  XNOR2_X1 U834 ( .A(n789), .B(n790), .ZN(n792) );
  NAND2_X1 U835 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U836 ( .A1(n794), .A2(n793), .ZN(G72) );
  XOR2_X1 U837 ( .A(G140), .B(n795), .Z(G42) );
  XOR2_X1 U838 ( .A(n796), .B(G101), .Z(G3) );
  XNOR2_X1 U839 ( .A(n797), .B(G122), .ZN(n798) );
  XNOR2_X1 U840 ( .A(n798), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U841 ( .A(G119), .B(n799), .Z(G21) );
  XOR2_X1 U842 ( .A(G134), .B(n800), .Z(G36) );
  XNOR2_X1 U843 ( .A(G137), .B(n801), .ZN(G39) );
endmodule

