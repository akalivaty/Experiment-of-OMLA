//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954;
  INV_X1    g000(.A(G43gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G50gat), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G43gat), .ZN(new_n205));
  AND3_X1   g004(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT15), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT14), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n209), .B(new_n211), .C1(new_n207), .C2(new_n208), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT90), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n203), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT89), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n205), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  AOI211_X1 g017(.A(new_n206), .B(new_n212), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n206), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT88), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G1gat), .B2(new_n224), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n227), .B(G8gat), .Z(new_n228));
  NOR2_X1   g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(new_n219), .B2(new_n222), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n220), .B(KEYINPUT88), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT15), .B1(new_n214), .B2(new_n216), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n212), .A2(new_n206), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n232), .B(KEYINPUT17), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT91), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n229), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n231), .A2(new_n235), .A3(KEYINPUT91), .A4(new_n228), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n238), .A2(KEYINPUT18), .A3(new_n239), .A4(new_n240), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n223), .B(new_n228), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n239), .B(KEYINPUT13), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT87), .ZN(new_n250));
  XNOR2_X1  g049(.A(G169gat), .B(G197gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT86), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n252), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT12), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n248), .B(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(G227gat), .A2(G233gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT27), .B(G183gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT28), .B1(new_n260), .B2(G190gat), .ZN(new_n261));
  INV_X1    g060(.A(G169gat), .ZN(new_n262));
  INV_X1    g061(.A(G176gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n264), .A2(KEYINPUT26), .ZN(new_n265));
  NAND2_X1  g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(KEYINPUT26), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n270));
  INV_X1    g069(.A(G190gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n259), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n261), .A2(new_n268), .A3(new_n269), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT23), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n266), .B1(new_n264), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT64), .B1(new_n276), .B2(KEYINPUT23), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n264), .A2(new_n278), .A3(new_n274), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT65), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n269), .A2(KEYINPUT24), .ZN(new_n282));
  XOR2_X1   g081(.A(G183gat), .B(G190gat), .Z(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(KEYINPUT24), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n281), .A2(KEYINPUT25), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n280), .A2(new_n286), .A3(new_n284), .A4(KEYINPUT25), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n273), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(KEYINPUT1), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G113gat), .B2(G120gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(G113gat), .B2(G120gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n292), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n273), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n277), .ZN(new_n299));
  INV_X1    g098(.A(new_n266), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n300), .B1(KEYINPUT23), .B2(new_n276), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT25), .B1(new_n302), .B2(new_n286), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n280), .A2(new_n284), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n298), .B1(new_n305), .B2(new_n287), .ZN(new_n306));
  INV_X1    g105(.A(new_n296), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n258), .B1(new_n297), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G15gat), .B(G43gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(G71gat), .B(G99gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n308), .A3(new_n258), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(KEYINPUT32), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT33), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(new_n314), .B2(new_n317), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(KEYINPUT32), .ZN(new_n322));
  INV_X1    g121(.A(new_n313), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(KEYINPUT33), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT34), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n321), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n321), .B2(new_n325), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n310), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n315), .ZN(new_n330));
  INV_X1    g129(.A(new_n320), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(new_n318), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT34), .B1(new_n332), .B2(new_n324), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n321), .A2(new_n325), .A3(new_n326), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n309), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G141gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G148gat), .ZN(new_n337));
  INV_X1    g136(.A(G148gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G141gat), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT2), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G155gat), .ZN(new_n341));
  INV_X1    g140(.A(G162gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OR3_X1    g144(.A1(new_n340), .A2(KEYINPUT73), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT73), .B1(new_n340), .B2(new_n345), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n337), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n336), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n339), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n344), .B1(new_n343), .B2(KEYINPUT2), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n346), .A2(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G197gat), .B(G204gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(G211gat), .A2(G218gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(KEYINPUT69), .A2(KEYINPUT22), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(KEYINPUT69), .A2(KEYINPUT22), .ZN(new_n358));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT70), .ZN(new_n360));
  OAI221_X1 g159(.A(new_n354), .B1(new_n357), .B2(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n353), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n353), .A2(new_n366), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n363), .B1(new_n368), .B2(new_n364), .ZN(new_n369));
  OAI211_X1 g168(.A(G228gat), .B(G233gat), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(G228gat), .B2(G233gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n366), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n346), .A2(new_n347), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n351), .A2(new_n352), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT76), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n353), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n372), .A2(new_n379), .A3(KEYINPUT80), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n371), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT80), .B1(new_n372), .B2(new_n379), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n370), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT31), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G22gat), .B(G50gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n385), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n370), .B(new_n388), .C1(new_n381), .C2(new_n382), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n387), .B1(new_n386), .B2(new_n389), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n329), .A2(new_n335), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n394));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n395), .B(KEYINPUT71), .Z(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n306), .B2(KEYINPUT29), .ZN(new_n397));
  INV_X1    g196(.A(new_n363), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n397), .B(new_n398), .C1(new_n306), .C2(new_n396), .ZN(new_n399));
  INV_X1    g198(.A(new_n396), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n289), .B2(new_n364), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n306), .A2(new_n396), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n363), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G64gat), .ZN(new_n406));
  INV_X1    g205(.A(G92gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT72), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT72), .ZN(new_n410));
  INV_X1    g209(.A(new_n408), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n399), .A2(new_n403), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n399), .B2(new_n403), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT30), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(KEYINPUT30), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT78), .ZN(new_n422));
  XOR2_X1   g221(.A(G1gat), .B(G29gat), .Z(new_n423));
  XOR2_X1   g222(.A(new_n422), .B(new_n423), .Z(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n375), .A2(new_n307), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n353), .A2(new_n296), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n427), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n429), .A2(KEYINPUT4), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n376), .A2(new_n296), .A3(new_n378), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n434), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n296), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n368), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n431), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n433), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n376), .A2(new_n296), .A3(new_n378), .A4(new_n436), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n429), .A2(KEYINPUT4), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n445), .A2(new_n427), .A3(new_n431), .A4(new_n440), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n420), .B(new_n426), .C1(new_n442), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n446), .ZN(new_n448));
  INV_X1    g247(.A(new_n426), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT6), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n442), .A2(new_n426), .A3(new_n446), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n394), .B1(new_n419), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n449), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n420), .A3(new_n451), .ZN(new_n455));
  INV_X1    g254(.A(new_n447), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n414), .B(new_n416), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(KEYINPUT79), .A3(new_n413), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT35), .B1(new_n393), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n419), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT83), .B1(new_n455), .B2(new_n456), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT83), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n447), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n462), .B(KEYINPUT84), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n456), .A2(KEYINPUT83), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n452), .B2(KEYINPUT83), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT84), .B1(new_n469), .B2(new_n462), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n329), .A2(new_n335), .A3(new_n392), .A4(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n461), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n443), .A2(new_n444), .B1(new_n368), .B2(new_n439), .ZN(new_n476));
  OAI211_X1 g275(.A(KEYINPUT39), .B(new_n475), .C1(new_n476), .C2(new_n431), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n445), .A2(new_n440), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT39), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n432), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n480), .A3(new_n426), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT40), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n454), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n458), .B2(new_n413), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT40), .B1(new_n481), .B2(KEYINPUT81), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT81), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n477), .A2(new_n480), .A3(new_n486), .A4(new_n426), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n485), .A2(KEYINPUT82), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT82), .B1(new_n485), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n484), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n404), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n399), .A2(new_n403), .A3(KEYINPUT37), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n411), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n415), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n408), .B1(new_n404), .B2(new_n491), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n493), .B1(new_n497), .B2(new_n494), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n451), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n426), .B1(new_n442), .B2(new_n446), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT6), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n464), .B1(new_n502), .B2(new_n447), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n503), .A3(new_n468), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n490), .A2(new_n504), .A3(new_n392), .ZN(new_n505));
  INV_X1    g304(.A(new_n392), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n460), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n329), .A2(new_n335), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(KEYINPUT68), .A2(KEYINPUT36), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(KEYINPUT68), .A2(KEYINPUT36), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n327), .A2(new_n328), .A3(new_n310), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n309), .B1(new_n333), .B2(new_n334), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n505), .A2(new_n507), .A3(new_n510), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n257), .B1(new_n474), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n519));
  INV_X1    g318(.A(G57gat), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n519), .B(G64gat), .C1(new_n520), .C2(KEYINPUT93), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n522));
  INV_X1    g321(.A(G64gat), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n522), .B(G57gat), .C1(new_n523), .C2(KEYINPUT92), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(G57gat), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n521), .B(new_n524), .C1(new_n519), .C2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G71gat), .ZN(new_n527));
  INV_X1    g326(.A(G78gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT9), .ZN(new_n529));
  NAND2_X1  g328(.A1(G71gat), .A2(G78gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n520), .A2(G64gat), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT9), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G71gat), .B(G78gat), .Z(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n532), .A2(KEYINPUT94), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT94), .B1(new_n532), .B2(new_n536), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n228), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(G183gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(G183gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n519), .A2(G64gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n520), .A2(KEYINPUT93), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n520), .A2(G64gat), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(KEYINPUT92), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n549), .A2(new_n521), .B1(new_n530), .B2(new_n529), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n526), .A2(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT94), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n559), .A3(new_n543), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G127gat), .B(G155gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT96), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT95), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n565), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT97), .B(G211gat), .Z(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n561), .A2(new_n562), .A3(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G85gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n576));
  OAI22_X1  g375(.A1(new_n575), .A2(new_n407), .B1(new_n576), .B2(KEYINPUT7), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n576), .A2(KEYINPUT100), .A3(KEYINPUT7), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT100), .B1(new_n576), .B2(KEYINPUT7), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n581), .A2(KEYINPUT99), .B1(G85gat), .B2(G92gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT100), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n581), .B2(KEYINPUT99), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n576), .A2(KEYINPUT100), .A3(KEYINPUT7), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT8), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n575), .A2(new_n407), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n588), .A2(KEYINPUT101), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT101), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n580), .B(new_n586), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT102), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n587), .ZN(new_n595));
  AND2_X1   g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT102), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n592), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT8), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(G99gat), .B2(G106gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n588), .A2(KEYINPUT101), .A3(new_n589), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n608), .A2(new_n599), .A3(new_n586), .A4(new_n580), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n231), .A2(new_n235), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT41), .ZN(new_n613));
  NAND2_X1  g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(KEYINPUT98), .Z(new_n615));
  OAI22_X1  g414(.A1(new_n223), .A2(new_n610), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT103), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n619), .A3(new_n611), .ZN(new_n620));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n617), .B2(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n615), .A2(new_n613), .ZN(new_n626));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n625), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n628), .B1(new_n631), .B2(new_n623), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n574), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n629), .B1(new_n624), .B2(new_n625), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n628), .A3(new_n623), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(KEYINPUT104), .A3(new_n574), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n555), .A2(new_n610), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n552), .A2(new_n554), .B1(new_n601), .B2(new_n609), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n601), .A2(new_n553), .A3(new_n609), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT105), .B1(new_n648), .B2(new_n643), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650));
  NOR4_X1   g449(.A1(new_n646), .A2(new_n647), .A3(new_n650), .A4(KEYINPUT10), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n645), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT106), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n555), .A2(new_n610), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n601), .A2(new_n553), .A3(new_n609), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n643), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n650), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n654), .A2(KEYINPUT105), .A3(new_n643), .A4(new_n655), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n644), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n642), .B1(new_n653), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G176gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(G204gat), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n663), .B1(new_n659), .B2(new_n642), .ZN(new_n670));
  INV_X1    g469(.A(new_n666), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n640), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n518), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n452), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT107), .B(G1gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1324gat));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n419), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(G8gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(G1325gat));
  NAND2_X1  g485(.A1(new_n329), .A2(new_n335), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(G15gat), .B1(new_n675), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n516), .A2(new_n510), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G15gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT108), .Z(new_n693));
  AOI21_X1  g492(.A(new_n689), .B1(new_n675), .B2(new_n693), .ZN(G1326gat));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n506), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  NOR2_X1   g496(.A1(new_n673), .A2(new_n574), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n638), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n518), .A2(new_n207), .A3(new_n452), .A4(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n699), .A2(new_n257), .ZN(new_n704));
  AOI211_X1 g503(.A(KEYINPUT44), .B(new_n638), .C1(new_n474), .C2(new_n517), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  INV_X1    g505(.A(new_n461), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n469), .A2(new_n462), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT84), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n473), .B1(new_n710), .B2(new_n466), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n517), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n638), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n706), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n704), .B1(new_n705), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT110), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n717), .B(new_n704), .C1(new_n705), .C2(new_n714), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n716), .A2(new_n452), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n703), .B1(new_n719), .B2(new_n207), .ZN(G1328gat));
  NAND4_X1  g519(.A1(new_n518), .A2(new_n208), .A3(new_n419), .A4(new_n700), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT46), .Z(new_n722));
  AND3_X1   g521(.A1(new_n716), .A2(new_n419), .A3(new_n718), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n208), .ZN(G1329gat));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n715), .B2(new_n690), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n712), .A2(new_n713), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT44), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n638), .B1(new_n474), .B2(new_n517), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n706), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n731), .A2(KEYINPUT111), .A3(new_n691), .A4(new_n704), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n726), .A2(G43gat), .A3(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n518), .A2(new_n700), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n734), .A2(new_n202), .A3(new_n688), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n716), .A2(new_n691), .A3(new_n718), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n735), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g540(.A(G50gat), .B1(new_n715), .B2(new_n392), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n506), .A2(new_n204), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT112), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(KEYINPUT48), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n745), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n716), .A2(new_n506), .A3(new_n718), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(G50gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n746), .B1(new_n749), .B2(KEYINPUT48), .ZN(G1331gat));
  XOR2_X1   g549(.A(new_n248), .B(new_n256), .Z(new_n751));
  AOI21_X1  g550(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n640), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n712), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n452), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n419), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT49), .B(G64gat), .Z(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n757), .B2(new_n759), .ZN(G1333gat));
  AOI21_X1  g559(.A(new_n527), .B1(new_n754), .B2(new_n691), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n687), .A2(G71gat), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n754), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n754), .A2(new_n506), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n574), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n727), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n729), .A2(KEYINPUT51), .A3(new_n768), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n752), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n575), .A3(new_n452), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n769), .A2(new_n752), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n728), .B2(new_n730), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n776), .A2(new_n452), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n773), .B1(new_n777), .B2(new_n575), .ZN(G1336gat));
  NAND2_X1  g577(.A1(new_n770), .A2(new_n771), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n462), .A2(G92gat), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n779), .A2(KEYINPUT113), .A3(new_n673), .A4(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n419), .B(new_n774), .C1(new_n705), .C2(new_n714), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G92gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT113), .B1(new_n772), .B2(new_n780), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT52), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(new_n772), .B2(new_n780), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n782), .A2(KEYINPUT114), .ZN(new_n788));
  OAI21_X1  g587(.A(G92gat), .B1(new_n782), .B2(KEYINPUT114), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(G1337gat));
  XNOR2_X1  g590(.A(KEYINPUT116), .B(G99gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n691), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n772), .A2(new_n688), .A3(new_n792), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1338gat));
  NAND2_X1  g597(.A1(new_n776), .A2(new_n506), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G106gat), .ZN(new_n800));
  INV_X1    g599(.A(G106gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n772), .A2(new_n801), .A3(new_n506), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT53), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n800), .A2(new_n805), .A3(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1339gat));
  NOR2_X1   g606(.A1(new_n419), .A2(new_n457), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n688), .A2(new_n392), .A3(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n635), .A2(new_n752), .A3(new_n639), .A4(new_n257), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n574), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n243), .A2(new_n256), .A3(new_n244), .A4(new_n247), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n239), .B1(new_n238), .B2(new_n240), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n245), .A2(new_n246), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n255), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n652), .A2(new_n821), .A3(new_n641), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n671), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n659), .A2(new_n660), .ZN(new_n824));
  AOI211_X1 g623(.A(KEYINPUT106), .B(new_n644), .C1(new_n657), .C2(new_n658), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n641), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n821), .B1(new_n659), .B2(new_n642), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n668), .B1(new_n828), .B2(KEYINPUT55), .ZN(new_n829));
  INV_X1    g628(.A(new_n827), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n671), .B(new_n822), .C1(new_n662), .C2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n820), .A2(new_n713), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n751), .A2(new_n829), .A3(new_n833), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n673), .A2(new_n814), .A3(new_n817), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n713), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n813), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n809), .B1(new_n812), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n751), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n673), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n574), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(G127gat), .ZN(G1342gat));
  AND2_X1   g645(.A1(new_n840), .A2(new_n713), .ZN(new_n847));
  INV_X1    g646(.A(G134gat), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT56), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n850), .B2(KEYINPUT56), .ZN(new_n853));
  OAI221_X1 g652(.A(new_n849), .B1(KEYINPUT56), .B2(new_n850), .C1(new_n852), .C2(new_n853), .ZN(G1343gat));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n837), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n638), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n574), .B1(new_n857), .B2(new_n834), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n810), .B(KEYINPUT117), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n855), .B(new_n506), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n690), .A2(new_n808), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n832), .B1(new_n828), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g663(.A(KEYINPUT120), .B(new_n823), .C1(new_n826), .C2(new_n827), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT121), .B(new_n829), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n751), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n831), .A2(KEYINPUT120), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n828), .A2(new_n863), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n832), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT121), .B1(new_n870), .B2(new_n829), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n837), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n638), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n574), .B1(new_n873), .B2(new_n834), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n506), .B1(new_n874), .B2(new_n859), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n862), .B1(new_n875), .B2(KEYINPUT57), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n336), .B1(new_n876), .B2(new_n751), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n392), .B1(new_n812), .B2(new_n839), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n861), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(G141gat), .A3(new_n257), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT58), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  INV_X1    g681(.A(new_n880), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n257), .B(new_n862), .C1(new_n875), .C2(KEYINPUT57), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n336), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n881), .A2(new_n885), .ZN(G1344gat));
  INV_X1    g685(.A(new_n879), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n338), .A3(new_n673), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT122), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT59), .B(new_n338), .C1(new_n876), .C2(new_n673), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  INV_X1    g690(.A(new_n810), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n855), .B(new_n506), .C1(new_n874), .C2(new_n892), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n878), .A2(new_n855), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n673), .A3(new_n861), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n889), .B1(new_n890), .B2(new_n896), .ZN(G1345gat));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n887), .B2(new_n574), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n879), .A2(KEYINPUT123), .A3(new_n813), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n899), .A2(new_n900), .A3(G155gat), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n813), .A2(new_n341), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n876), .B2(new_n902), .ZN(G1346gat));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n342), .A3(new_n713), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n876), .A2(new_n713), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n342), .ZN(G1347gat));
  NAND2_X1  g705(.A1(new_n812), .A2(new_n839), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n393), .A2(new_n452), .A3(new_n462), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n257), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(new_n262), .ZN(G1348gat));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n752), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(new_n263), .ZN(G1349gat));
  INV_X1    g712(.A(new_n909), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n259), .A3(new_n574), .ZN(new_n915));
  NAND2_X1  g714(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n916));
  OAI21_X1  g715(.A(G183gat), .B1(new_n909), .B2(new_n813), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n918), .B(new_n919), .Z(G1350gat));
  OAI22_X1  g719(.A1(new_n909), .A2(new_n638), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n921), .B(new_n922), .ZN(G1351gat));
  NOR2_X1   g722(.A1(new_n462), .A2(new_n452), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n690), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n878), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n751), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n893), .A2(new_n894), .A3(new_n925), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n751), .A2(G197gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  NOR3_X1   g731(.A1(new_n926), .A2(G204gat), .A3(new_n752), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT62), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n893), .A2(new_n673), .A3(new_n894), .ZN(new_n935));
  INV_X1    g734(.A(new_n925), .ZN(new_n936));
  OAI21_X1  g735(.A(G204gat), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(G1353gat));
  OAI21_X1  g737(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n940), .B1(new_n929), .B2(new_n813), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT63), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  OAI221_X1 g744(.A(new_n940), .B1(new_n942), .B2(new_n943), .C1(new_n929), .C2(new_n813), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n926), .A2(G211gat), .A3(new_n813), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G1354gat));
  AOI21_X1  g747(.A(G218gat), .B1(new_n927), .B2(new_n713), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n713), .A2(G218gat), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT127), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n930), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(G1355gat));
endmodule


