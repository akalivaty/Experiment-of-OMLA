//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G43gat), .ZN(new_n209));
  INV_X1    g008(.A(G43gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G50gat), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT15), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT15), .B1(new_n209), .B2(new_n211), .ZN(new_n213));
  NAND2_X1  g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT84), .A2(G29gat), .A3(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n212), .A2(new_n213), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220));
  INV_X1    g019(.A(new_n206), .ZN(new_n221));
  NOR3_X1   g020(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n216), .A2(new_n217), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n205), .A2(KEYINPUT83), .A3(new_n206), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n207), .A2(new_n219), .B1(new_n226), .B2(new_n212), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n212), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n218), .ZN(new_n230));
  INV_X1    g029(.A(new_n212), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(new_n207), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT7), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(KEYINPUT93), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G99gat), .ZN(new_n241));
  INV_X1    g040(.A(G106gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G99gat), .A2(G106gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT94), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT94), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n247), .A3(new_n244), .ZN(new_n248));
  INV_X1    g047(.A(G85gat), .ZN(new_n249));
  INV_X1    g048(.A(G92gat), .ZN(new_n250));
  AOI22_X1  g049(.A1(KEYINPUT8), .A2(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n240), .A2(new_n246), .A3(new_n248), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n238), .A2(new_n239), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n244), .A2(KEYINPUT8), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(G85gat), .B2(G92gat), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT94), .B(new_n245), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n228), .A2(new_n235), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT41), .ZN(new_n260));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261));
  OAI221_X1 g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .C1(new_n227), .C2(new_n258), .ZN(new_n262));
  XNOR2_X1  g061(.A(G190gat), .B(G218gat), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G134gat), .B(G162gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n260), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT95), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n263), .ZN(new_n270));
  MUX2_X1   g069(.A(new_n267), .B(new_n268), .S(new_n270), .Z(new_n271));
  AOI21_X1  g070(.A(new_n269), .B1(new_n271), .B2(new_n264), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(G71gat), .A2(G78gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(G71gat), .A2(G78gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G57gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G64gat), .ZN(new_n283));
  INV_X1    g082(.A(G64gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G57gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G78gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n280), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n281), .A2(new_n289), .A3(KEYINPUT91), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT91), .B1(new_n281), .B2(new_n289), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT21), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT92), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295));
  INV_X1    g094(.A(G1gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT16), .ZN(new_n297));
  INV_X1    g096(.A(G15gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G22gat), .ZN(new_n299));
  INV_X1    g098(.A(G22gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G15gat), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n297), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(G1gat), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n302), .A2(new_n303), .A3(G8gat), .ZN(new_n304));
  INV_X1    g103(.A(G8gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n301), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n296), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n297), .A2(new_n299), .A3(new_n301), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n295), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(G8gat), .B1(new_n302), .B2(new_n303), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n305), .A3(new_n308), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT85), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n294), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n294), .B1(new_n293), .B2(new_n314), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n275), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n317), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(new_n315), .A3(new_n274), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n292), .A2(KEYINPUT21), .ZN(new_n321));
  XOR2_X1   g120(.A(G183gat), .B(G211gat), .Z(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  NAND3_X1  g122(.A1(new_n318), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(G127gat), .B(G155gat), .Z(new_n326));
  NAND2_X1  g125(.A1(G231gat), .A2(G233gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n323), .B1(new_n318), .B2(new_n320), .ZN(new_n330));
  OR3_X1    g129(.A1(new_n325), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n325), .B2(new_n330), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n256), .B(new_n252), .C1(new_n290), .C2(new_n291), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT10), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n287), .B1(new_n288), .B2(new_n286), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n257), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n257), .A2(KEYINPUT10), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT91), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n337), .B2(new_n338), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n281), .A2(new_n289), .A3(KEYINPUT91), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT96), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT96), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n292), .A2(new_n348), .A3(KEYINPUT10), .A4(new_n257), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n341), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT97), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G230gat), .A2(G233gat), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n341), .A2(new_n347), .A3(KEYINPUT97), .A4(new_n349), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G120gat), .B(G148gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G176gat), .B(G204gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n353), .B1(new_n335), .B2(new_n340), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT98), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n360), .A2(KEYINPUT98), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n355), .A2(new_n359), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n358), .B(KEYINPUT99), .Z(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n361), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n350), .A2(new_n353), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n273), .A2(new_n334), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G1gat), .B(G29gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(new_n249), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT0), .B(G57gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT2), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377));
  INV_X1    g176(.A(G141gat), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n378), .A2(G148gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(G148gat), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n376), .B(new_n377), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G155gat), .B(G162gat), .Z(new_n384));
  OR2_X1    g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n376), .B1(new_n379), .B2(new_n380), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n383), .B(new_n384), .C1(new_n382), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT66), .ZN(new_n391));
  INV_X1    g190(.A(G127gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(G134gat), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT66), .B1(new_n392), .B2(G134gat), .ZN(new_n394));
  INV_X1    g193(.A(G134gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(G127gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n393), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT67), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G113gat), .B(G120gat), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n400), .A2(KEYINPUT1), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n392), .A2(G134gat), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n401), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n387), .A3(KEYINPUT3), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n404), .B1(new_n399), .B2(new_n401), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n388), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n410), .B2(new_n388), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n408), .B(new_n409), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n410), .B(new_n388), .ZN(new_n418));
  INV_X1    g217(.A(new_n409), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n374), .B(new_n417), .C1(new_n421), .C2(new_n416), .ZN(new_n422));
  INV_X1    g221(.A(new_n374), .ZN(new_n423));
  INV_X1    g222(.A(new_n417), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n416), .B1(new_n415), .B2(new_n420), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n424), .A2(new_n425), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n374), .A3(new_n427), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G197gat), .B(G204gat), .ZN(new_n434));
  INV_X1    g233(.A(G211gat), .ZN(new_n435));
  INV_X1    g234(.A(G218gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n434), .B1(KEYINPUT22), .B2(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(G211gat), .B(G218gat), .Z(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(G169gat), .A2(G176gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT23), .ZN(new_n442));
  NAND2_X1  g241(.A1(G169gat), .A2(G176gat), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(G169gat), .B2(G176gat), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT24), .ZN(new_n447));
  INV_X1    g246(.A(G183gat), .ZN(new_n448));
  INV_X1    g247(.A(G190gat), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n450), .B(new_n451), .C1(G183gat), .C2(G190gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n446), .A2(KEYINPUT64), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT25), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT64), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT25), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n446), .A3(new_n452), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT65), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT27), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(G183gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT27), .B(G183gat), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n449), .B(new_n462), .C1(new_n463), .C2(new_n460), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT28), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(G190gat), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n464), .A2(new_n465), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n441), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT26), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n443), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n441), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n455), .B(new_n459), .C1(new_n467), .C2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT29), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n475), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(KEYINPUT73), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT73), .B1(new_n472), .B2(new_n477), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n440), .B(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n440), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n472), .A2(new_n477), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n477), .B1(new_n472), .B2(new_n473), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(KEYINPUT74), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT73), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n485), .B1(new_n489), .B2(new_n478), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT74), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(new_n440), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT37), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(KEYINPUT75), .B(G8gat), .Z(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT76), .B(G36gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G64gat), .B(G92gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n482), .B(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n440), .B1(new_n484), .B2(new_n485), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n500), .A2(KEYINPUT37), .A3(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n493), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n492), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT37), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT38), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI22_X1  g305(.A1(new_n503), .A2(KEYINPUT38), .B1(new_n493), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n499), .B1(new_n504), .B2(KEYINPUT38), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n433), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT31), .B(G22gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(G228gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n390), .A2(new_n473), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n482), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT3), .B1(new_n440), .B2(new_n473), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n515), .A2(new_n388), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n208), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n208), .B1(new_n514), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n512), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n519), .ZN(new_n521));
  INV_X1    g320(.A(new_n512), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G78gat), .B(G106gat), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(new_n520), .B2(new_n523), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n504), .A2(new_n499), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n487), .A2(new_n492), .A3(new_n498), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n504), .A2(KEYINPUT30), .A3(new_n499), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n408), .B1(new_n413), .B2(new_n414), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n419), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(KEYINPUT39), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n535), .B(KEYINPUT39), .C1(new_n419), .C2(new_n418), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(new_n423), .ZN(new_n538));
  NOR2_X1   g337(.A1(KEYINPUT81), .A2(KEYINPUT40), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT81), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT40), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n533), .A2(new_n540), .A3(new_n422), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n509), .A2(new_n527), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT36), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT68), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n406), .B2(new_n472), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n455), .A2(new_n459), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n467), .A2(new_n471), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n549), .A2(new_n410), .A3(new_n550), .A4(KEYINPUT68), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n406), .A2(new_n472), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(G227gat), .A2(G233gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT33), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G15gat), .B(G43gat), .ZN(new_n556));
  INV_X1    g355(.A(G71gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT69), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G99gat), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n553), .A2(new_n554), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT32), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT71), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT32), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n555), .A2(new_n560), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT32), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n565), .B1(new_n562), .B2(KEYINPUT32), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n572));
  OAI22_X1  g371(.A1(new_n553), .A2(new_n554), .B1(new_n572), .B2(KEYINPUT34), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(KEYINPUT34), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n567), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n575), .B1(new_n567), .B2(new_n571), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n546), .B1(new_n579), .B2(KEYINPUT72), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n532), .A2(new_n531), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT77), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT77), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n532), .A2(new_n583), .A3(new_n531), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n582), .A2(new_n432), .A3(new_n530), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n525), .A2(new_n526), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n588), .B(KEYINPUT36), .C1(new_n577), .C2(new_n578), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n545), .A2(new_n580), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n578), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(new_n527), .A3(new_n576), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT35), .B1(new_n592), .B2(new_n585), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n577), .A2(new_n586), .A3(new_n578), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n433), .A2(new_n533), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT35), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT85), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT85), .B1(new_n311), .B2(new_n312), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n227), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n233), .A2(new_n310), .A3(new_n313), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n605), .B(KEYINPUT13), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT86), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n304), .A2(new_n309), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n228), .A2(new_n235), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n605), .A4(new_n603), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n604), .A2(KEYINPUT86), .A3(new_n606), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n609), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n610), .B1(new_n227), .B2(KEYINPUT17), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n233), .A2(new_n234), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n605), .B(new_n603), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT18), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n619), .A2(KEYINPUT88), .ZN(new_n620));
  XOR2_X1   g419(.A(G169gat), .B(G197gat), .Z(new_n621));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n619), .A2(KEYINPUT88), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n614), .A2(new_n620), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n609), .A2(new_n619), .A3(new_n612), .A4(new_n613), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT87), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n630), .A2(new_n631), .A3(new_n626), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n630), .B2(new_n626), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT89), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(KEYINPUT89), .B(new_n629), .C1(new_n632), .C2(new_n633), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n599), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT90), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n599), .A2(KEYINPUT90), .A3(new_n639), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n370), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n433), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT100), .B(G1gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1324gat));
  XNOR2_X1  g446(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT90), .B1(new_n599), .B2(new_n639), .ZN(new_n649));
  AOI211_X1 g448(.A(new_n641), .B(new_n638), .C1(new_n590), .C2(new_n598), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n533), .B(new_n369), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT16), .B(G8gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT102), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n648), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g455(.A(KEYINPUT103), .B(new_n648), .C1(new_n651), .C2(new_n653), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n651), .A2(G8gat), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n652), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n660), .B1(new_n651), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n644), .A2(KEYINPUT104), .A3(new_n533), .A4(new_n662), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n658), .A2(new_n659), .A3(new_n664), .A4(new_n665), .ZN(G1325gat));
  OAI21_X1  g465(.A(new_n369), .B1(new_n649), .B2(new_n650), .ZN(new_n667));
  INV_X1    g466(.A(new_n579), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n298), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n580), .A2(new_n589), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(G15gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT105), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n644), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT106), .ZN(G1326gat));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n644), .A2(new_n676), .A3(new_n586), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT107), .B1(new_n667), .B2(new_n527), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n679), .B(new_n681), .ZN(G1327gat));
  AOI21_X1  g481(.A(new_n272), .B1(new_n590), .B2(new_n598), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n368), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n334), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n634), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n685), .A2(new_n433), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G29gat), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n687), .B1(new_n642), .B2(new_n643), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n273), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n432), .A2(G29gat), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR4_X1   g496(.A1(new_n694), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n432), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n691), .B1(new_n697), .B2(new_n698), .ZN(G1328gat));
  NAND4_X1  g498(.A1(new_n693), .A2(new_n204), .A3(new_n533), .A4(new_n273), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n700), .A2(KEYINPUT46), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n533), .A3(new_n689), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G36gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(KEYINPUT46), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(G1329gat));
  NAND4_X1  g504(.A1(new_n693), .A2(new_n210), .A3(new_n579), .A4(new_n273), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n684), .B1(new_n599), .B2(new_n273), .ZN(new_n707));
  AOI211_X1 g506(.A(KEYINPUT44), .B(new_n272), .C1(new_n590), .C2(new_n598), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n670), .B(new_n689), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT47), .B1(new_n710), .B2(KEYINPUT108), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n706), .B(new_n710), .C1(KEYINPUT108), .C2(KEYINPUT47), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1330gat));
  NAND4_X1  g514(.A1(new_n693), .A2(new_n208), .A3(new_n586), .A4(new_n273), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT48), .B1(new_n716), .B2(KEYINPUT109), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n586), .B(new_n689), .C1(new_n707), .C2(new_n708), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G50gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n716), .B(new_n719), .C1(KEYINPUT109), .C2(KEYINPUT48), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1331gat));
  AOI21_X1  g522(.A(new_n634), .B1(new_n590), .B2(new_n598), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n273), .A2(new_n334), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n725), .A3(new_n368), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n432), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n282), .ZN(G1332gat));
  INV_X1    g527(.A(new_n726), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT49), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n284), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(new_n533), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT110), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n729), .A2(new_n735), .A3(new_n533), .A4(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n730), .A2(new_n284), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n729), .A2(new_n557), .A3(new_n579), .ZN(new_n740));
  INV_X1    g539(.A(new_n670), .ZN(new_n741));
  OAI21_X1  g540(.A(G71gat), .B1(new_n726), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n586), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g546(.A1(new_n333), .A2(new_n634), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n599), .A2(new_n273), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT51), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n683), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n433), .A3(new_n368), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n748), .A2(new_n368), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT112), .Z(new_n756));
  NAND3_X1  g555(.A1(new_n685), .A2(G85gat), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n249), .A2(new_n754), .B1(new_n758), .B2(new_n433), .ZN(G1336gat));
  OAI211_X1 g558(.A(new_n533), .B(new_n756), .C1(new_n707), .C2(new_n708), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n750), .A2(new_n533), .A3(new_n368), .A4(new_n752), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(G92gat), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT52), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n685), .A2(new_n670), .A3(new_n756), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G99gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n753), .A2(new_n241), .A3(new_n368), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n668), .ZN(G1338gat));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n586), .A3(new_n368), .A4(new_n752), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n242), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n685), .A2(G106gat), .A3(new_n586), .A4(new_n756), .ZN(new_n772));
  AOI211_X1 g571(.A(KEYINPUT113), .B(new_n769), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n769), .A2(KEYINPUT113), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(KEYINPUT113), .ZN(new_n775));
  AND4_X1   g574(.A1(new_n774), .A2(new_n771), .A3(new_n775), .A4(new_n772), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n773), .A2(new_n776), .ZN(G1339gat));
  NAND2_X1  g576(.A1(new_n369), .A2(new_n688), .ZN(new_n778));
  INV_X1    g577(.A(new_n353), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n341), .A2(new_n347), .A3(new_n779), .A4(new_n349), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(KEYINPUT54), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n355), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n359), .B1(new_n366), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n784), .A3(KEYINPUT55), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n784), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n782), .A2(new_n784), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n787), .A2(new_n790), .A3(new_n363), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n605), .B1(new_n611), .B2(new_n603), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n604), .A2(new_n606), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n625), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n629), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n272), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n368), .A2(new_n629), .A3(new_n795), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n792), .B2(new_n688), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(new_n799), .B2(new_n272), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n778), .B1(new_n800), .B2(new_n333), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n594), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n533), .A2(new_n432), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(G113gat), .B1(new_n804), .B2(new_n638), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n688), .A2(G113gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n804), .B2(new_n806), .ZN(G1340gat));
  INV_X1    g606(.A(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n368), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g609(.A1(new_n804), .A2(new_n334), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(new_n392), .ZN(G1342gat));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n273), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n813), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(G134gat), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT56), .B1(new_n813), .B2(G134gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(G1343gat));
  NOR3_X1   g616(.A1(new_n670), .A2(new_n432), .A3(new_n533), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n586), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  XOR2_X1   g619(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n787), .A2(new_n363), .A3(new_n791), .ZN(new_n824));
  XNOR2_X1  g623(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n788), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n824), .A2(new_n636), .A3(new_n637), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n273), .B1(new_n827), .B2(new_n798), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n334), .B1(new_n828), .B2(new_n797), .ZN(new_n829));
  AOI211_X1 g628(.A(new_n823), .B(new_n527), .C1(new_n829), .C2(new_n778), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n818), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n378), .B1(new_n832), .B2(new_n639), .ZN(new_n833));
  INV_X1    g632(.A(new_n818), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n834), .A2(new_n819), .A3(G141gat), .A4(new_n638), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT58), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n634), .B(new_n818), .C1(new_n822), .C2(new_n830), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n837), .B2(G141gat), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n833), .A2(new_n836), .B1(new_n838), .B2(new_n839), .ZN(G1344gat));
  AND3_X1   g639(.A1(new_n801), .A2(new_n586), .A3(new_n821), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n369), .A2(new_n638), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n787), .A2(new_n826), .A3(new_n363), .A4(new_n791), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n798), .B1(new_n638), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n797), .B1(new_n844), .B2(new_n272), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n842), .B1(new_n845), .B2(new_n333), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n848), .B(new_n842), .C1(new_n845), .C2(new_n333), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n586), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n841), .B1(new_n850), .B2(new_n823), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n686), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n818), .A2(KEYINPUT117), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n818), .A2(KEYINPUT117), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT59), .B(G148gat), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G148gat), .B1(new_n831), .B2(new_n686), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n834), .A2(new_n819), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n686), .A2(G148gat), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n857), .A2(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n856), .A2(new_n861), .ZN(G1345gat));
  AOI21_X1  g661(.A(G155gat), .B1(new_n859), .B2(new_n333), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n333), .A2(G155gat), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT119), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n832), .B2(new_n865), .ZN(G1346gat));
  AOI21_X1  g665(.A(G162gat), .B1(new_n859), .B2(new_n273), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n273), .A2(G162gat), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n832), .B2(new_n868), .ZN(G1347gat));
  AND2_X1   g668(.A1(new_n533), .A2(new_n432), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n802), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(G169gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n634), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n870), .B(KEYINPUT120), .Z(new_n874));
  AND2_X1   g673(.A1(new_n802), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(new_n639), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n876), .B2(new_n872), .ZN(G1348gat));
  AOI21_X1  g676(.A(G176gat), .B1(new_n871), .B2(new_n368), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n875), .A2(G176gat), .A3(new_n368), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT122), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(G1349gat));
  NAND2_X1  g682(.A1(new_n875), .A2(new_n333), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n884), .A2(G183gat), .B1(new_n885), .B2(KEYINPUT60), .ZN(new_n886));
  NAND2_X1  g685(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT124), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n463), .A3(new_n333), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n888), .B1(new_n886), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(G1350gat));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n273), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G190gat), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(KEYINPUT125), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n449), .A3(new_n273), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n893), .A2(G190gat), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(G1351gat));
  AND3_X1   g700(.A1(new_n820), .A2(new_n741), .A3(new_n870), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT126), .ZN(new_n903));
  INV_X1    g702(.A(G197gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n904), .A3(new_n634), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n874), .A2(new_n741), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n851), .A2(new_n638), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n907), .B2(new_n904), .ZN(G1352gat));
  INV_X1    g707(.A(new_n902), .ZN(new_n909));
  INV_X1    g708(.A(G204gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n368), .A2(new_n910), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n909), .A2(KEYINPUT62), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT62), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n851), .A2(new_n686), .A3(new_n906), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n912), .B(new_n913), .C1(new_n910), .C2(new_n914), .ZN(G1353gat));
  NAND3_X1  g714(.A1(new_n903), .A2(new_n435), .A3(new_n333), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n851), .A2(new_n334), .A3(new_n906), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n917), .A2(new_n918), .A3(new_n435), .ZN(new_n919));
  INV_X1    g718(.A(new_n906), .ZN(new_n920));
  INV_X1    g719(.A(new_n849), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n848), .B1(new_n829), .B2(new_n842), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n923), .B2(new_n586), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n333), .B(new_n920), .C1(new_n924), .C2(new_n841), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT63), .B1(new_n925), .B2(G211gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n916), .B1(new_n919), .B2(new_n926), .ZN(G1354gat));
  OAI211_X1 g726(.A(KEYINPUT127), .B(new_n920), .C1(new_n924), .C2(new_n841), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n929), .B1(new_n851), .B2(new_n906), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n273), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G218gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n903), .A2(new_n436), .A3(new_n273), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1355gat));
endmodule


