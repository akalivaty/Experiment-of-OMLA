

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U552 ( .A(n807), .Z(n517) );
  XNOR2_X1 U553 ( .A(n548), .B(n547), .ZN(n807) );
  NOR2_X1 U554 ( .A1(n750), .A2(n749), .ZN(n751) );
  AND2_X1 U555 ( .A1(n692), .A2(n691), .ZN(n694) );
  AND2_X2 U556 ( .A1(n534), .A2(G2105), .ZN(n907) );
  XNOR2_X1 U557 ( .A(n539), .B(G543), .ZN(n576) );
  NOR2_X1 U558 ( .A1(n638), .A2(n998), .ZN(n639) );
  INV_X1 U559 ( .A(KEYINPUT65), .ZN(n547) );
  XNOR2_X1 U560 ( .A(n603), .B(KEYINPUT93), .ZN(n604) );
  INV_X1 U561 ( .A(KEYINPUT28), .ZN(n614) );
  XNOR2_X1 U562 ( .A(n663), .B(KEYINPUT30), .ZN(n664) );
  NOR2_X1 U563 ( .A1(G1966), .A2(n713), .ZN(n683) );
  AND2_X1 U564 ( .A1(n697), .A2(n695), .ZN(n696) );
  INV_X1 U565 ( .A(KEYINPUT33), .ZN(n695) );
  INV_X1 U566 ( .A(G2104), .ZN(n524) );
  XNOR2_X1 U567 ( .A(KEYINPUT66), .B(G2104), .ZN(n527) );
  INV_X1 U568 ( .A(n1007), .ZN(n702) );
  BUF_X1 U569 ( .A(n720), .Z(n903) );
  NOR2_X1 U570 ( .A1(n635), .A2(n634), .ZN(n637) );
  XOR2_X1 U571 ( .A(KEYINPUT31), .B(n668), .Z(n518) );
  AND2_X1 U572 ( .A1(n523), .A2(n648), .ZN(n519) );
  XOR2_X1 U573 ( .A(n694), .B(n693), .Z(n520) );
  AND2_X1 U574 ( .A1(n645), .A2(n644), .ZN(n521) );
  AND2_X1 U575 ( .A1(n640), .A2(n639), .ZN(n522) );
  OR2_X1 U576 ( .A1(n646), .A2(n991), .ZN(n523) );
  INV_X1 U577 ( .A(n680), .ZN(n661) );
  OR2_X1 U578 ( .A1(n683), .A2(n662), .ZN(n663) );
  XNOR2_X1 U579 ( .A(n615), .B(n614), .ZN(n651) );
  INV_X1 U580 ( .A(KEYINPUT29), .ZN(n652) );
  INV_X1 U581 ( .A(KEYINPUT95), .ZN(n676) );
  INV_X1 U582 ( .A(KEYINPUT97), .ZN(n693) );
  XNOR2_X1 U583 ( .A(n679), .B(KEYINPUT32), .ZN(n705) );
  NAND2_X1 U584 ( .A1(G8), .A2(n660), .ZN(n713) );
  XNOR2_X1 U585 ( .A(n704), .B(KEYINPUT99), .ZN(n717) );
  NAND2_X1 U586 ( .A1(n807), .A2(G54), .ZN(n618) );
  NOR2_X1 U587 ( .A1(n717), .A2(n716), .ZN(n750) );
  XNOR2_X1 U588 ( .A(KEYINPUT71), .B(KEYINPUT14), .ZN(n632) );
  INV_X1 U589 ( .A(G2105), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n633), .B(n632), .ZN(n634) );
  AND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n720) );
  AND2_X1 U592 ( .A1(n622), .A2(n621), .ZN(n623) );
  INV_X1 U593 ( .A(KEYINPUT0), .ZN(n539) );
  OR2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n525), .B(KEYINPUT17), .ZN(n594) );
  NAND2_X1 U596 ( .A1(n637), .A2(n636), .ZN(n998) );
  BUF_X1 U597 ( .A(n594), .Z(n902) );
  BUF_X1 U598 ( .A(n601), .Z(G164) );
  INV_X1 U599 ( .A(KEYINPUT89), .ZN(n530) );
  NAND2_X1 U600 ( .A1(n524), .A2(n526), .ZN(n525) );
  NAND2_X1 U601 ( .A1(n594), .A2(G138), .ZN(n529) );
  NAND2_X1 U602 ( .A1(n720), .A2(G102), .ZN(n528) );
  NAND2_X1 U603 ( .A1(n529), .A2(n528), .ZN(n531) );
  NAND2_X1 U604 ( .A1(n530), .A2(n531), .ZN(n533) );
  NAND2_X1 U605 ( .A1(n533), .A2(n532), .ZN(n538) );
  AND2_X1 U606 ( .A1(G2104), .A2(G2105), .ZN(n906) );
  NAND2_X1 U607 ( .A1(G114), .A2(n906), .ZN(n536) );
  XOR2_X1 U608 ( .A(KEYINPUT66), .B(G2104), .Z(n534) );
  NAND2_X1 U609 ( .A1(G126), .A2(n907), .ZN(n535) );
  NAND2_X1 U610 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U611 ( .A1(n538), .A2(n537), .ZN(n601) );
  XNOR2_X1 U612 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n544) );
  NOR2_X2 U613 ( .A1(G651), .A2(G543), .ZN(n814) );
  NAND2_X1 U614 ( .A1(G90), .A2(n814), .ZN(n541) );
  INV_X1 U615 ( .A(G651), .ZN(n545) );
  NOR2_X1 U616 ( .A1(n576), .A2(n545), .ZN(n811) );
  NAND2_X1 U617 ( .A1(G77), .A2(n811), .ZN(n540) );
  NAND2_X1 U618 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U619 ( .A(n542), .B(KEYINPUT9), .ZN(n543) );
  XNOR2_X1 U620 ( .A(n544), .B(n543), .ZN(n552) );
  NOR2_X1 U621 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X2 U622 ( .A(KEYINPUT1), .B(n546), .Z(n806) );
  NAND2_X1 U623 ( .A1(G64), .A2(n806), .ZN(n550) );
  NOR2_X1 U624 ( .A1(G651), .A2(n576), .ZN(n548) );
  NAND2_X1 U625 ( .A1(G52), .A2(n517), .ZN(n549) );
  NAND2_X1 U626 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U627 ( .A1(n552), .A2(n551), .ZN(G171) );
  NAND2_X1 U628 ( .A1(G89), .A2(n814), .ZN(n553) );
  XNOR2_X1 U629 ( .A(n553), .B(KEYINPUT76), .ZN(n554) );
  XNOR2_X1 U630 ( .A(n554), .B(KEYINPUT4), .ZN(n556) );
  NAND2_X1 U631 ( .A1(G76), .A2(n811), .ZN(n555) );
  NAND2_X1 U632 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U633 ( .A(n557), .B(KEYINPUT5), .ZN(n562) );
  NAND2_X1 U634 ( .A1(G63), .A2(n806), .ZN(n559) );
  NAND2_X1 U635 ( .A1(G51), .A2(n517), .ZN(n558) );
  NAND2_X1 U636 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U637 ( .A(KEYINPUT6), .B(n560), .Z(n561) );
  NAND2_X1 U638 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U639 ( .A(n563), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U640 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U641 ( .A1(n517), .A2(G50), .ZN(n564) );
  XOR2_X1 U642 ( .A(KEYINPUT85), .B(n564), .Z(n566) );
  NAND2_X1 U643 ( .A1(n806), .A2(G62), .ZN(n565) );
  NAND2_X1 U644 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U645 ( .A(KEYINPUT86), .B(n567), .Z(n571) );
  NAND2_X1 U646 ( .A1(G88), .A2(n814), .ZN(n569) );
  NAND2_X1 U647 ( .A1(G75), .A2(n811), .ZN(n568) );
  AND2_X1 U648 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U649 ( .A1(n571), .A2(n570), .ZN(G303) );
  NAND2_X1 U650 ( .A1(G49), .A2(n517), .ZN(n573) );
  NAND2_X1 U651 ( .A1(G74), .A2(G651), .ZN(n572) );
  NAND2_X1 U652 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U653 ( .A(KEYINPUT83), .B(n574), .Z(n575) );
  NOR2_X1 U654 ( .A1(n806), .A2(n575), .ZN(n578) );
  NAND2_X1 U655 ( .A1(n576), .A2(G87), .ZN(n577) );
  NAND2_X1 U656 ( .A1(n578), .A2(n577), .ZN(G288) );
  NAND2_X1 U657 ( .A1(G73), .A2(n811), .ZN(n579) );
  XNOR2_X1 U658 ( .A(n579), .B(KEYINPUT2), .ZN(n586) );
  NAND2_X1 U659 ( .A1(G48), .A2(n517), .ZN(n581) );
  NAND2_X1 U660 ( .A1(G86), .A2(n814), .ZN(n580) );
  NAND2_X1 U661 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n806), .A2(G61), .ZN(n582) );
  XOR2_X1 U663 ( .A(KEYINPUT84), .B(n582), .Z(n583) );
  NOR2_X1 U664 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U665 ( .A1(n586), .A2(n585), .ZN(G305) );
  NAND2_X1 U666 ( .A1(n517), .A2(G47), .ZN(n588) );
  NAND2_X1 U667 ( .A1(n806), .A2(G60), .ZN(n587) );
  NAND2_X1 U668 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U669 ( .A(KEYINPUT67), .B(n589), .ZN(n593) );
  NAND2_X1 U670 ( .A1(G85), .A2(n814), .ZN(n591) );
  NAND2_X1 U671 ( .A1(G72), .A2(n811), .ZN(n590) );
  AND2_X1 U672 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n593), .A2(n592), .ZN(G290) );
  NAND2_X1 U674 ( .A1(n902), .A2(G137), .ZN(n771) );
  AND2_X1 U675 ( .A1(n771), .A2(G40), .ZN(n600) );
  NAND2_X1 U676 ( .A1(G113), .A2(n906), .ZN(n596) );
  NAND2_X1 U677 ( .A1(G125), .A2(n907), .ZN(n595) );
  AND2_X1 U678 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U679 ( .A1(G101), .A2(n720), .ZN(n597) );
  XOR2_X1 U680 ( .A(KEYINPUT23), .B(n597), .Z(n598) );
  AND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n770) );
  NAND2_X1 U682 ( .A1(n600), .A2(n770), .ZN(n718) );
  INV_X1 U683 ( .A(n718), .ZN(n602) );
  NOR2_X2 U684 ( .A1(n601), .A2(G1384), .ZN(n719) );
  NAND2_X2 U685 ( .A1(n602), .A2(n719), .ZN(n660) );
  INV_X2 U686 ( .A(n660), .ZN(n654) );
  NAND2_X1 U687 ( .A1(G2072), .A2(n654), .ZN(n605) );
  INV_X1 U688 ( .A(KEYINPUT27), .ZN(n603) );
  XNOR2_X1 U689 ( .A(n605), .B(n604), .ZN(n607) );
  AND2_X1 U690 ( .A1(n660), .A2(G1956), .ZN(n606) );
  NOR2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n647) );
  NAND2_X1 U692 ( .A1(G65), .A2(n806), .ZN(n609) );
  NAND2_X1 U693 ( .A1(G53), .A2(n517), .ZN(n608) );
  NAND2_X1 U694 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U695 ( .A1(G91), .A2(n814), .ZN(n611) );
  NAND2_X1 U696 ( .A1(G78), .A2(n811), .ZN(n610) );
  NAND2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n822) );
  NOR2_X1 U699 ( .A1(n647), .A2(n822), .ZN(n615) );
  NAND2_X1 U700 ( .A1(G92), .A2(n814), .ZN(n617) );
  NAND2_X1 U701 ( .A1(G79), .A2(n811), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n617), .A2(n616), .ZN(n620) );
  XNOR2_X1 U703 ( .A(KEYINPUT75), .B(n618), .ZN(n619) );
  NOR2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n806), .A2(G66), .ZN(n621) );
  XNOR2_X2 U706 ( .A(n623), .B(KEYINPUT15), .ZN(n991) );
  NAND2_X1 U707 ( .A1(G1348), .A2(n660), .ZN(n625) );
  NAND2_X1 U708 ( .A1(G2067), .A2(n654), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n646) );
  NAND2_X1 U710 ( .A1(n991), .A2(n646), .ZN(n640) );
  XNOR2_X1 U711 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n642) );
  NOR2_X1 U712 ( .A1(G1996), .A2(n642), .ZN(n638) );
  XNOR2_X1 U713 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G81), .A2(n814), .ZN(n626) );
  XNOR2_X1 U715 ( .A(n626), .B(KEYINPUT72), .ZN(n627) );
  XNOR2_X1 U716 ( .A(n627), .B(KEYINPUT12), .ZN(n629) );
  NAND2_X1 U717 ( .A1(G68), .A2(n811), .ZN(n628) );
  NAND2_X1 U718 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U719 ( .A(n631), .B(n630), .ZN(n635) );
  NAND2_X1 U720 ( .A1(G56), .A2(n806), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n517), .A2(G43), .ZN(n636) );
  INV_X1 U722 ( .A(G1341), .ZN(n999) );
  NAND2_X1 U723 ( .A1(n999), .A2(n642), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n641), .A2(n660), .ZN(n645) );
  AND2_X1 U725 ( .A1(G1996), .A2(n654), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n522), .A2(n521), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n647), .A2(n822), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n519), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n659) );
  OR2_X1 U732 ( .A1(n654), .A2(G1961), .ZN(n656) );
  XNOR2_X1 U733 ( .A(G2078), .B(KEYINPUT25), .ZN(n1015) );
  NAND2_X1 U734 ( .A1(n654), .A2(n1015), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n656), .A2(n655), .ZN(n665) );
  AND2_X1 U736 ( .A1(n665), .A2(G171), .ZN(n657) );
  XOR2_X1 U737 ( .A(KEYINPUT92), .B(n657), .Z(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n669) );
  NOR2_X1 U739 ( .A1(G2084), .A2(n660), .ZN(n680) );
  NAND2_X1 U740 ( .A1(n661), .A2(G8), .ZN(n662) );
  NOR2_X1 U741 ( .A1(G168), .A2(n664), .ZN(n667) );
  NOR2_X1 U742 ( .A1(G171), .A2(n665), .ZN(n666) );
  NOR2_X1 U743 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U744 ( .A1(n669), .A2(n518), .ZN(n681) );
  NAND2_X1 U745 ( .A1(n681), .A2(G286), .ZN(n675) );
  NOR2_X1 U746 ( .A1(G1971), .A2(n713), .ZN(n671) );
  NOR2_X1 U747 ( .A1(G2090), .A2(n660), .ZN(n670) );
  NOR2_X1 U748 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U749 ( .A1(n672), .A2(G303), .ZN(n673) );
  XNOR2_X1 U750 ( .A(n673), .B(KEYINPUT94), .ZN(n674) );
  NAND2_X1 U751 ( .A1(n675), .A2(n674), .ZN(n677) );
  XNOR2_X1 U752 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U753 ( .A1(n678), .A2(G8), .ZN(n679) );
  NAND2_X1 U754 ( .A1(G8), .A2(n680), .ZN(n685) );
  INV_X1 U755 ( .A(n681), .ZN(n682) );
  NOR2_X1 U756 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U757 ( .A1(n685), .A2(n684), .ZN(n706) );
  NAND2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n993) );
  AND2_X1 U759 ( .A1(n706), .A2(n993), .ZN(n686) );
  NAND2_X1 U760 ( .A1(n705), .A2(n686), .ZN(n692) );
  INV_X1 U761 ( .A(n993), .ZN(n690) );
  NOR2_X1 U762 ( .A1(G1976), .A2(G288), .ZN(n995) );
  NOR2_X1 U763 ( .A1(G1971), .A2(G303), .ZN(n687) );
  XNOR2_X1 U764 ( .A(KEYINPUT96), .B(n687), .ZN(n688) );
  NOR2_X1 U765 ( .A1(n995), .A2(n688), .ZN(n689) );
  OR2_X1 U766 ( .A1(n690), .A2(n689), .ZN(n691) );
  INV_X1 U767 ( .A(n713), .ZN(n697) );
  NAND2_X1 U768 ( .A1(n520), .A2(n696), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n995), .A2(n697), .ZN(n698) );
  NAND2_X1 U770 ( .A1(n698), .A2(KEYINPUT33), .ZN(n699) );
  NAND2_X1 U771 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U772 ( .A(n701), .B(KEYINPUT98), .ZN(n703) );
  XNOR2_X1 U773 ( .A(G1981), .B(G305), .ZN(n1007) );
  NAND2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U775 ( .A1(n706), .A2(n705), .ZN(n709) );
  NOR2_X1 U776 ( .A1(G2090), .A2(G303), .ZN(n707) );
  NAND2_X1 U777 ( .A1(G8), .A2(n707), .ZN(n708) );
  NAND2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n710), .A2(n713), .ZN(n715) );
  NOR2_X1 U780 ( .A1(G1981), .A2(G305), .ZN(n711) );
  XOR2_X1 U781 ( .A(n711), .B(KEYINPUT24), .Z(n712) );
  OR2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n765) );
  NAND2_X1 U785 ( .A1(G140), .A2(n902), .ZN(n722) );
  NAND2_X1 U786 ( .A1(G104), .A2(n903), .ZN(n721) );
  NAND2_X1 U787 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U788 ( .A(KEYINPUT34), .B(n723), .ZN(n728) );
  NAND2_X1 U789 ( .A1(G116), .A2(n906), .ZN(n725) );
  NAND2_X1 U790 ( .A1(G128), .A2(n907), .ZN(n724) );
  NAND2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U792 ( .A(n726), .B(KEYINPUT35), .Z(n727) );
  NOR2_X1 U793 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U794 ( .A(KEYINPUT36), .B(n729), .Z(n730) );
  XOR2_X1 U795 ( .A(KEYINPUT90), .B(n730), .Z(n919) );
  XNOR2_X1 U796 ( .A(KEYINPUT37), .B(G2067), .ZN(n762) );
  NOR2_X1 U797 ( .A1(n919), .A2(n762), .ZN(n963) );
  NAND2_X1 U798 ( .A1(n765), .A2(n963), .ZN(n760) );
  NAND2_X1 U799 ( .A1(G131), .A2(n902), .ZN(n732) );
  NAND2_X1 U800 ( .A1(G95), .A2(n903), .ZN(n731) );
  NAND2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n736) );
  NAND2_X1 U802 ( .A1(G107), .A2(n906), .ZN(n734) );
  NAND2_X1 U803 ( .A1(G119), .A2(n907), .ZN(n733) );
  NAND2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U805 ( .A1(n736), .A2(n735), .ZN(n914) );
  INV_X1 U806 ( .A(G1991), .ZN(n1021) );
  NOR2_X1 U807 ( .A1(n914), .A2(n1021), .ZN(n745) );
  NAND2_X1 U808 ( .A1(G141), .A2(n902), .ZN(n738) );
  NAND2_X1 U809 ( .A1(G117), .A2(n906), .ZN(n737) );
  NAND2_X1 U810 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U811 ( .A1(n903), .A2(G105), .ZN(n739) );
  XOR2_X1 U812 ( .A(KEYINPUT38), .B(n739), .Z(n740) );
  NOR2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U814 ( .A1(n907), .A2(G129), .ZN(n742) );
  NAND2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n892) );
  AND2_X1 U816 ( .A1(n892), .A2(G1996), .ZN(n744) );
  NOR2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n968) );
  INV_X1 U818 ( .A(n765), .ZN(n746) );
  NOR2_X1 U819 ( .A1(n968), .A2(n746), .ZN(n757) );
  INV_X1 U820 ( .A(n757), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n760), .A2(n747), .ZN(n748) );
  XOR2_X1 U822 ( .A(KEYINPUT91), .B(n748), .Z(n749) );
  XNOR2_X1 U823 ( .A(n751), .B(KEYINPUT100), .ZN(n753) );
  XNOR2_X1 U824 ( .A(G1986), .B(G290), .ZN(n1005) );
  NAND2_X1 U825 ( .A1(n1005), .A2(n765), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n768) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n892), .ZN(n978) );
  AND2_X1 U828 ( .A1(n1021), .A2(n914), .ZN(n970) );
  NOR2_X1 U829 ( .A1(G1986), .A2(G290), .ZN(n754) );
  XOR2_X1 U830 ( .A(n754), .B(KEYINPUT101), .Z(n755) );
  NOR2_X1 U831 ( .A1(n970), .A2(n755), .ZN(n756) );
  NOR2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U833 ( .A1(n978), .A2(n758), .ZN(n759) );
  XNOR2_X1 U834 ( .A(KEYINPUT39), .B(n759), .ZN(n761) );
  NAND2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U836 ( .A1(n919), .A2(n762), .ZN(n962) );
  NAND2_X1 U837 ( .A1(n763), .A2(n962), .ZN(n764) );
  XNOR2_X1 U838 ( .A(KEYINPUT102), .B(n764), .ZN(n766) );
  NAND2_X1 U839 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U840 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U841 ( .A(n769), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U842 ( .A1(n771), .A2(n770), .ZN(G160) );
  XOR2_X1 U843 ( .A(G2443), .B(G2446), .Z(n773) );
  XNOR2_X1 U844 ( .A(G2427), .B(G2451), .ZN(n772) );
  XNOR2_X1 U845 ( .A(n773), .B(n772), .ZN(n779) );
  XOR2_X1 U846 ( .A(G2430), .B(G2454), .Z(n775) );
  XNOR2_X1 U847 ( .A(G1341), .B(G1348), .ZN(n774) );
  XNOR2_X1 U848 ( .A(n775), .B(n774), .ZN(n777) );
  XOR2_X1 U849 ( .A(G2435), .B(G2438), .Z(n776) );
  XNOR2_X1 U850 ( .A(n777), .B(n776), .ZN(n778) );
  XOR2_X1 U851 ( .A(n779), .B(n778), .Z(n780) );
  AND2_X1 U852 ( .A1(G14), .A2(n780), .ZN(G401) );
  AND2_X1 U853 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U854 ( .A1(G135), .A2(n902), .ZN(n782) );
  NAND2_X1 U855 ( .A1(G111), .A2(n906), .ZN(n781) );
  NAND2_X1 U856 ( .A1(n782), .A2(n781), .ZN(n787) );
  NAND2_X1 U857 ( .A1(G123), .A2(n907), .ZN(n783) );
  XNOR2_X1 U858 ( .A(n783), .B(KEYINPUT18), .ZN(n785) );
  NAND2_X1 U859 ( .A1(n903), .A2(G99), .ZN(n784) );
  NAND2_X1 U860 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U861 ( .A1(n787), .A2(n786), .ZN(n966) );
  XNOR2_X1 U862 ( .A(n966), .B(G2096), .ZN(n788) );
  XNOR2_X1 U863 ( .A(n788), .B(KEYINPUT79), .ZN(n789) );
  OR2_X1 U864 ( .A1(G2100), .A2(n789), .ZN(G156) );
  INV_X1 U865 ( .A(n822), .ZN(G299) );
  INV_X1 U866 ( .A(G57), .ZN(G237) );
  INV_X1 U867 ( .A(G132), .ZN(G219) );
  INV_X1 U868 ( .A(G82), .ZN(G220) );
  NAND2_X1 U869 ( .A1(G7), .A2(G661), .ZN(n790) );
  XNOR2_X1 U870 ( .A(n790), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U871 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n792) );
  INV_X1 U872 ( .A(G223), .ZN(n849) );
  NAND2_X1 U873 ( .A1(G567), .A2(n849), .ZN(n791) );
  XNOR2_X1 U874 ( .A(n792), .B(n791), .ZN(G234) );
  INV_X1 U875 ( .A(G860), .ZN(n798) );
  NOR2_X1 U876 ( .A1(n998), .A2(n798), .ZN(n793) );
  XOR2_X1 U877 ( .A(KEYINPUT74), .B(n793), .Z(G153) );
  INV_X1 U878 ( .A(G171), .ZN(G301) );
  NAND2_X1 U879 ( .A1(G868), .A2(G301), .ZN(n795) );
  INV_X1 U880 ( .A(G868), .ZN(n833) );
  NAND2_X1 U881 ( .A1(n991), .A2(n833), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(G284) );
  NOR2_X1 U883 ( .A1(G286), .A2(n833), .ZN(n797) );
  NOR2_X1 U884 ( .A1(G868), .A2(G299), .ZN(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(G297) );
  NAND2_X1 U886 ( .A1(n798), .A2(G559), .ZN(n799) );
  INV_X1 U887 ( .A(n991), .ZN(n818) );
  NAND2_X1 U888 ( .A1(n799), .A2(n818), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n800), .B(KEYINPUT16), .ZN(n802) );
  XOR2_X1 U890 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n801) );
  XNOR2_X1 U891 ( .A(n802), .B(n801), .ZN(G148) );
  NOR2_X1 U892 ( .A1(G868), .A2(n998), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G868), .A2(n818), .ZN(n803) );
  NOR2_X1 U894 ( .A1(G559), .A2(n803), .ZN(n804) );
  NOR2_X1 U895 ( .A1(n805), .A2(n804), .ZN(G282) );
  NAND2_X1 U896 ( .A1(G67), .A2(n806), .ZN(n809) );
  NAND2_X1 U897 ( .A1(G55), .A2(n517), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U899 ( .A(KEYINPUT82), .B(n810), .Z(n813) );
  NAND2_X1 U900 ( .A1(n811), .A2(G80), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n817) );
  NAND2_X1 U902 ( .A1(G93), .A2(n814), .ZN(n815) );
  XNOR2_X1 U903 ( .A(KEYINPUT81), .B(n815), .ZN(n816) );
  OR2_X1 U904 ( .A1(n817), .A2(n816), .ZN(n832) );
  XNOR2_X1 U905 ( .A(KEYINPUT80), .B(n998), .ZN(n819) );
  NAND2_X1 U906 ( .A1(n818), .A2(G559), .ZN(n830) );
  XNOR2_X1 U907 ( .A(n819), .B(n830), .ZN(n820) );
  NOR2_X1 U908 ( .A1(G860), .A2(n820), .ZN(n821) );
  XOR2_X1 U909 ( .A(n832), .B(n821), .Z(G145) );
  INV_X1 U910 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U911 ( .A(n822), .B(n998), .ZN(n823) );
  XNOR2_X1 U912 ( .A(n823), .B(G305), .ZN(n824) );
  XOR2_X1 U913 ( .A(n824), .B(KEYINPUT87), .Z(n826) );
  XOR2_X1 U914 ( .A(n832), .B(KEYINPUT19), .Z(n825) );
  XNOR2_X1 U915 ( .A(n826), .B(n825), .ZN(n827) );
  XNOR2_X1 U916 ( .A(n827), .B(G290), .ZN(n828) );
  XNOR2_X1 U917 ( .A(n828), .B(G288), .ZN(n829) );
  XNOR2_X1 U918 ( .A(G166), .B(n829), .ZN(n922) );
  XNOR2_X1 U919 ( .A(n830), .B(n922), .ZN(n831) );
  NAND2_X1 U920 ( .A1(n831), .A2(G868), .ZN(n835) );
  NAND2_X1 U921 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U922 ( .A1(n835), .A2(n834), .ZN(G295) );
  NAND2_X1 U923 ( .A1(G2078), .A2(G2084), .ZN(n836) );
  XOR2_X1 U924 ( .A(KEYINPUT20), .B(n836), .Z(n837) );
  NAND2_X1 U925 ( .A1(G2090), .A2(n837), .ZN(n838) );
  XNOR2_X1 U926 ( .A(KEYINPUT21), .B(n838), .ZN(n839) );
  NAND2_X1 U927 ( .A1(n839), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U928 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U929 ( .A1(G220), .A2(G219), .ZN(n840) );
  XOR2_X1 U930 ( .A(KEYINPUT22), .B(n840), .Z(n841) );
  NOR2_X1 U931 ( .A1(G218), .A2(n841), .ZN(n842) );
  XNOR2_X1 U932 ( .A(KEYINPUT88), .B(n842), .ZN(n843) );
  NAND2_X1 U933 ( .A1(n843), .A2(G96), .ZN(n853) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n853), .ZN(n847) );
  NAND2_X1 U935 ( .A1(G69), .A2(G120), .ZN(n844) );
  NOR2_X1 U936 ( .A1(G237), .A2(n844), .ZN(n845) );
  NAND2_X1 U937 ( .A1(G108), .A2(n845), .ZN(n854) );
  NAND2_X1 U938 ( .A1(G567), .A2(n854), .ZN(n846) );
  NAND2_X1 U939 ( .A1(n847), .A2(n846), .ZN(n855) );
  NAND2_X1 U940 ( .A1(G483), .A2(G661), .ZN(n848) );
  NOR2_X1 U941 ( .A1(n855), .A2(n848), .ZN(n852) );
  NAND2_X1 U942 ( .A1(n852), .A2(G36), .ZN(G176) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n849), .ZN(G217) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n850) );
  NAND2_X1 U945 ( .A1(G661), .A2(n850), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n851) );
  NAND2_X1 U947 ( .A1(n852), .A2(n851), .ZN(G188) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  INV_X1 U951 ( .A(G69), .ZN(G235) );
  NOR2_X1 U952 ( .A1(n854), .A2(n853), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U954 ( .A(KEYINPUT103), .B(n855), .ZN(G319) );
  XOR2_X1 U955 ( .A(G2096), .B(G2678), .Z(n857) );
  XNOR2_X1 U956 ( .A(G2072), .B(KEYINPUT43), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n858), .B(KEYINPUT42), .Z(n860) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2090), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U961 ( .A(KEYINPUT104), .B(G2100), .Z(n862) );
  XNOR2_X1 U962 ( .A(G2078), .B(G2084), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(G227) );
  XOR2_X1 U965 ( .A(G1976), .B(G1961), .Z(n866) );
  XNOR2_X1 U966 ( .A(G1986), .B(G1956), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U968 ( .A(G1981), .B(G1966), .Z(n868) );
  XNOR2_X1 U969 ( .A(G1996), .B(G1991), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U971 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U972 ( .A(KEYINPUT105), .B(G2474), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n874) );
  XOR2_X1 U974 ( .A(G1971), .B(KEYINPUT41), .Z(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(G229) );
  NAND2_X1 U976 ( .A1(G136), .A2(n902), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G112), .A2(n906), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G124), .A2(n907), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n877), .B(KEYINPUT106), .ZN(n878) );
  XNOR2_X1 U981 ( .A(KEYINPUT44), .B(n878), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G100), .A2(n903), .ZN(n879) );
  XOR2_X1 U983 ( .A(KEYINPUT107), .B(n879), .Z(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U985 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U986 ( .A1(G118), .A2(n906), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G130), .A2(n907), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G142), .A2(n902), .ZN(n887) );
  NAND2_X1 U990 ( .A1(G106), .A2(n903), .ZN(n886) );
  NAND2_X1 U991 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n888), .Z(n889) );
  NOR2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U994 ( .A(G164), .B(n891), .ZN(n918) );
  XOR2_X1 U995 ( .A(n966), .B(G162), .Z(n894) );
  XOR2_X1 U996 ( .A(G160), .B(n892), .Z(n893) );
  XNOR2_X1 U997 ( .A(n894), .B(n893), .ZN(n901) );
  XOR2_X1 U998 ( .A(KEYINPUT112), .B(KEYINPUT110), .Z(n896) );
  XNOR2_X1 U999 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n895) );
  XNOR2_X1 U1000 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U1001 ( .A(n897), .B(KEYINPUT108), .Z(n899) );
  XNOR2_X1 U1002 ( .A(KEYINPUT111), .B(KEYINPUT113), .ZN(n898) );
  XNOR2_X1 U1003 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U1004 ( .A(n901), .B(n900), .Z(n916) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n902), .ZN(n905) );
  NAND2_X1 U1006 ( .A1(G103), .A2(n903), .ZN(n904) );
  NAND2_X1 U1007 ( .A1(n905), .A2(n904), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(G115), .A2(n906), .ZN(n909) );
  NAND2_X1 U1009 ( .A1(G127), .A2(n907), .ZN(n908) );
  NAND2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(KEYINPUT109), .B(n910), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(KEYINPUT47), .B(n911), .ZN(n912) );
  NOR2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n973) );
  XNOR2_X1 U1014 ( .A(n914), .B(n973), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n920), .B(n919), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n921), .ZN(G395) );
  XNOR2_X1 U1019 ( .A(n922), .B(KEYINPUT114), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(G171), .B(G286), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n924), .B(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n925), .B(n991), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n926), .ZN(G397) );
  NOR2_X1 U1024 ( .A1(G227), .A2(G229), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(n928), .B(n927), .ZN(n929) );
  XOR2_X1 U1027 ( .A(KEYINPUT49), .B(n929), .Z(n930) );
  NOR2_X1 U1028 ( .A1(G401), .A2(n930), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(G319), .A2(n931), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT117), .B(n932), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(G395), .A2(G397), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(G225) );
  INV_X1 U1033 ( .A(G225), .ZN(G308) );
  INV_X1 U1034 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1035 ( .A(G1348), .B(KEYINPUT59), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(n935), .B(G4), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G1341), .B(G19), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(G1981), .B(G6), .ZN(n936) );
  NOR2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n942) );
  XOR2_X1 U1041 ( .A(KEYINPUT123), .B(G1956), .Z(n940) );
  XNOR2_X1 U1042 ( .A(G20), .B(n940), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1044 ( .A(KEYINPUT60), .B(n943), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G1986), .B(KEYINPUT126), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(n944), .B(G24), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(G1971), .B(G22), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(G1976), .B(G23), .ZN(n945) );
  NOR2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1050 ( .A(n947), .B(KEYINPUT125), .ZN(n948) );
  NOR2_X1 U1051 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1052 ( .A(KEYINPUT58), .B(n950), .Z(n952) );
  XNOR2_X1 U1053 ( .A(G1961), .B(G5), .ZN(n951) );
  NOR2_X1 U1054 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(KEYINPUT124), .B(G1966), .ZN(n955) );
  XNOR2_X1 U1057 ( .A(G21), .B(n955), .ZN(n956) );
  NOR2_X1 U1058 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1059 ( .A(KEYINPUT61), .B(n958), .ZN(n960) );
  INV_X1 U1060 ( .A(G16), .ZN(n959) );
  NAND2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1062 ( .A1(n961), .A2(G11), .ZN(n990) );
  INV_X1 U1063 ( .A(n962), .ZN(n964) );
  NOR2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n972) );
  XOR2_X1 U1065 ( .A(G2084), .B(G160), .Z(n965) );
  NOR2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n983) );
  XOR2_X1 U1070 ( .A(G2072), .B(n973), .Z(n975) );
  XOR2_X1 U1071 ( .A(G164), .B(G2078), .Z(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(KEYINPUT50), .B(n976), .ZN(n981) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n979), .Z(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT52), .B(n984), .ZN(n986) );
  INV_X1 U1080 ( .A(KEYINPUT55), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n987), .A2(G29), .ZN(n988) );
  XOR2_X1 U1083 ( .A(KEYINPUT118), .B(n988), .Z(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n1041) );
  XOR2_X1 U1085 ( .A(KEYINPUT56), .B(G16), .Z(n1014) );
  XNOR2_X1 U1086 ( .A(G166), .B(G1971), .ZN(n997) );
  XOR2_X1 U1087 ( .A(G1348), .B(n991), .Z(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n1012) );
  XNOR2_X1 U1091 ( .A(n999), .B(n998), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G299), .B(G1956), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(G301), .B(G1961), .ZN(n1000) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(G168), .B(G1966), .Z(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(KEYINPUT57), .B(n1008), .Z(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1039) );
  XOR2_X1 U1103 ( .A(n1015), .B(G27), .Z(n1020) );
  XNOR2_X1 U1104 ( .A(G2067), .B(G26), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(G2072), .B(G33), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(KEYINPUT121), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(n1021), .B(G25), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(G28), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(n1023), .B(KEYINPUT120), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(G1996), .B(G32), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(n1028), .B(KEYINPUT53), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(G2084), .B(G34), .Z(n1029) );
  XNOR2_X1 U1117 ( .A(KEYINPUT54), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1034) );
  XOR2_X1 U1119 ( .A(KEYINPUT119), .B(G2090), .Z(n1032) );
  XNOR2_X1 U1120 ( .A(G35), .B(n1032), .ZN(n1033) );
  NOR2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1122 ( .A(KEYINPUT55), .B(n1035), .Z(n1036) );
  XNOR2_X1 U1123 ( .A(KEYINPUT122), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1124 ( .A1(G29), .A2(n1037), .ZN(n1038) );
  NOR2_X1 U1125 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1127 ( .A(KEYINPUT62), .B(n1042), .ZN(n1043) );
  XNOR2_X1 U1128 ( .A(KEYINPUT127), .B(n1043), .ZN(G311) );
  INV_X1 U1129 ( .A(G311), .ZN(G150) );
endmodule

