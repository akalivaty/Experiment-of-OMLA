//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT82), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G952), .ZN(new_n191));
  NAND2_X1  g005(.A1(G234), .A2(G237), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n193), .B(KEYINPUT97), .Z(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(G902), .A3(G953), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT21), .B(G898), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n199), .B(KEYINPUT98), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT84), .ZN(new_n201));
  XNOR2_X1  g015(.A(G110), .B(G122), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT6), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G101), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G116), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT2), .B(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G113), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT2), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT2), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G113), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G116), .B(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n219), .A2(new_n226), .A3(KEYINPUT68), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT68), .B1(new_n219), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n212), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n210), .A2(G101), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n231));
  INV_X1    g045(.A(G101), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n205), .A2(new_n208), .A3(new_n232), .A4(new_n209), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT4), .A4(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n210), .A2(G101), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT80), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n229), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n220), .B1(new_n225), .B2(KEYINPUT5), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n214), .B2(KEYINPUT5), .ZN(new_n241));
  OR3_X1    g055(.A1(new_n214), .A2(new_n240), .A3(KEYINPUT5), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n207), .A2(G104), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n204), .A2(G107), .ZN(new_n245));
  OAI21_X1  g059(.A(G101), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n233), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n243), .A2(new_n247), .A3(new_n226), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n201), .B(new_n203), .C1(new_n238), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n237), .A2(new_n234), .ZN(new_n250));
  INV_X1    g064(.A(new_n212), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n219), .A2(new_n226), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n219), .A2(new_n226), .A3(KEYINPUT68), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n248), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n203), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT84), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n257), .B2(new_n202), .ZN(new_n262));
  INV_X1    g076(.A(new_n202), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n263), .B1(new_n238), .B2(new_n248), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT1), .A3(G146), .ZN(new_n267));
  XNOR2_X1  g081(.A(G143), .B(G146), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G128), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G143), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(G146), .ZN(new_n273));
  AND4_X1   g087(.A1(new_n270), .A2(new_n272), .A3(new_n273), .A4(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G125), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT0), .ZN(new_n278));
  INV_X1    g092(.A(G128), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n272), .A2(new_n273), .ZN(new_n282));
  NOR2_X1   g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n268), .A2(KEYINPUT0), .A3(G128), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G125), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n277), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n190), .A2(G224), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n289), .B(new_n290), .Z(new_n291));
  NAND3_X1  g105(.A1(new_n260), .A2(new_n265), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(KEYINPUT7), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n277), .A2(new_n288), .A3(KEYINPUT7), .A4(new_n290), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n296), .B1(new_n257), .B2(new_n202), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n243), .A2(new_n226), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n233), .A2(new_n246), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(KEYINPUT85), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n202), .B(KEYINPUT8), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n299), .B2(new_n301), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n298), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n299), .A2(new_n301), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(KEYINPUT86), .A3(new_n302), .A4(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(G902), .B1(new_n297), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n311), .B(KEYINPUT87), .Z(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n292), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n313), .B1(new_n292), .B2(new_n310), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n189), .B(new_n200), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT9), .B(G234), .ZN(new_n318));
  OAI21_X1  g132(.A(G221), .B1(new_n318), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT11), .ZN(new_n321));
  INV_X1    g135(.A(G137), .ZN(new_n322));
  OAI22_X1  g136(.A1(KEYINPUT65), .A2(new_n321), .B1(new_n322), .B2(G134), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n324));
  INV_X1    g138(.A(G134), .ZN(new_n325));
  OAI22_X1  g139(.A1(new_n324), .A2(KEYINPUT11), .B1(new_n325), .B2(G137), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT65), .A4(G134), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G131), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n320), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n324), .A2(KEYINPUT11), .B1(new_n325), .B2(G137), .ZN(new_n331));
  AND4_X1   g145(.A1(KEYINPUT65), .A2(new_n321), .A3(new_n322), .A4(G134), .ZN(new_n332));
  AOI22_X1  g146(.A1(KEYINPUT65), .A2(new_n321), .B1(new_n322), .B2(G134), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT67), .A3(G131), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n329), .B(new_n331), .C1(new_n332), .C2(new_n333), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT66), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n326), .A2(new_n327), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n340), .A2(KEYINPUT66), .A3(new_n329), .A4(new_n331), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n344));
  AOI21_X1  g158(.A(G128), .B1(new_n272), .B2(new_n273), .ZN(new_n345));
  INV_X1    g159(.A(new_n267), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n268), .A2(new_n270), .A3(G128), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n267), .B(KEYINPUT81), .C1(new_n268), .C2(G128), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT10), .B1(new_n350), .B2(new_n247), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n275), .A2(new_n352), .A3(new_n300), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n212), .A2(new_n286), .A3(new_n285), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n237), .B2(new_n234), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n343), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n351), .A2(new_n353), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n330), .A2(new_n335), .B1(new_n339), .B2(new_n341), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n190), .A2(G227), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT79), .ZN(new_n363));
  XNOR2_X1  g177(.A(G110), .B(G140), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n357), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n350), .A2(new_n247), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n275), .A2(new_n300), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT12), .B1(new_n370), .B2(new_n343), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n343), .A3(KEYINPUT12), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n356), .A2(new_n351), .A3(new_n353), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n372), .A2(new_n373), .B1(new_n374), .B2(new_n360), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n367), .B(G469), .C1(new_n375), .C2(new_n366), .ZN(new_n376));
  INV_X1    g190(.A(G469), .ZN(new_n377));
  INV_X1    g191(.A(G902), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NOR4_X1   g195(.A1(new_n356), .A2(new_n343), .A3(new_n351), .A4(new_n353), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n360), .B1(new_n358), .B2(new_n359), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n365), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n373), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n361), .B(new_n366), .C1(new_n385), .C2(new_n371), .ZN(new_n386));
  AOI211_X1 g200(.A(G469), .B(G902), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n319), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n279), .A2(G143), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n325), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G128), .B(G143), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n393), .B2(new_n389), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n325), .ZN(new_n395));
  XNOR2_X1  g209(.A(G116), .B(G122), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n207), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n266), .A2(G128), .ZN(new_n399));
  OAI21_X1  g213(.A(G134), .B1(new_n390), .B2(new_n399), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n395), .A2(new_n400), .B1(new_n396), .B2(new_n207), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT94), .ZN(new_n402));
  INV_X1    g216(.A(G122), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(G116), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT14), .B1(new_n403), .B2(G116), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n215), .A3(G122), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(G107), .C1(KEYINPUT94), .C2(new_n407), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n401), .A2(new_n409), .A3(KEYINPUT95), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT95), .B1(new_n401), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n398), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G217), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n318), .A2(new_n413), .A3(G953), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n398), .B(new_n414), .C1(new_n410), .C2(new_n411), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT96), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT96), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n412), .A2(new_n419), .A3(new_n415), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n378), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n422), .A2(KEYINPUT15), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n421), .B(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n425));
  NOR2_X1   g239(.A1(G475), .A2(G902), .ZN(new_n426));
  XNOR2_X1  g240(.A(G113), .B(G122), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(new_n204), .ZN(new_n428));
  INV_X1    g242(.A(G237), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n190), .A3(G214), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n266), .ZN(new_n431));
  NOR2_X1   g245(.A1(G237), .A2(G953), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(G143), .A3(G214), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(KEYINPUT88), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(KEYINPUT18), .A2(G131), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n435), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n431), .A2(KEYINPUT88), .A3(new_n437), .A4(new_n433), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G140), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n276), .B2(KEYINPUT74), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT74), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(G125), .A3(G140), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(G146), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(G125), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n276), .A2(G140), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(new_n271), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n439), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT89), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT89), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n439), .A2(new_n452), .A3(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n431), .A2(new_n433), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G131), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n431), .A2(new_n329), .A3(new_n433), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT91), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n441), .A2(KEYINPUT19), .A3(new_n443), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT19), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n445), .A2(new_n446), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n461), .B1(new_n465), .B2(G146), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n462), .A2(KEYINPUT91), .A3(new_n464), .A4(new_n271), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n441), .A2(KEYINPUT16), .A3(new_n443), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT16), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n445), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G146), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n456), .A2(KEYINPUT90), .A3(new_n457), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n460), .A2(new_n468), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n428), .B1(new_n454), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n456), .A2(new_n477), .A3(new_n457), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n469), .A2(new_n271), .A3(new_n471), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n455), .A2(KEYINPUT17), .A3(G131), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n478), .A2(new_n479), .A3(new_n473), .A4(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(KEYINPUT89), .B(new_n448), .C1(new_n436), .C2(new_n438), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n452), .B1(new_n439), .B2(new_n449), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n428), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n425), .B(new_n426), .C1(new_n476), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT92), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n475), .B1(new_n482), .B2(new_n483), .ZN(new_n488));
  INV_X1    g302(.A(new_n428), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n484), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n425), .A4(new_n426), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n426), .B1(new_n476), .B2(new_n485), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT20), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n428), .B1(new_n454), .B2(new_n481), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n378), .B1(new_n497), .B2(new_n485), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G475), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n424), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n317), .A2(new_n388), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n254), .A2(new_n255), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  INV_X1    g317(.A(new_n287), .ZN(new_n504));
  XOR2_X1   g318(.A(G134), .B(G137), .Z(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G131), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n269), .B2(new_n274), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n339), .B2(new_n341), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n343), .A2(new_n504), .B1(new_n508), .B2(KEYINPUT69), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n345), .A2(new_n346), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n510), .A2(new_n348), .B1(G131), .B2(new_n505), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n342), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT69), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n503), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n287), .A2(KEYINPUT64), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT64), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n285), .A2(new_n286), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n503), .B(new_n512), .C1(new_n360), .C2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n502), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT31), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n343), .A2(new_n504), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT66), .B1(new_n328), .B2(new_n329), .ZN(new_n525));
  INV_X1    g339(.A(new_n341), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n511), .B(KEYINPUT69), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n227), .B2(new_n228), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n255), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n524), .A2(new_n514), .A3(new_n527), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n432), .A2(G210), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT27), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT26), .B(G101), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n522), .A2(new_n523), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n502), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n527), .B1(new_n360), .B2(new_n287), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT30), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n540), .B1(new_n543), .B2(new_n520), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT31), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  INV_X1    g359(.A(new_n536), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n529), .A2(new_n530), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n512), .B1(new_n360), .B2(new_n287), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT72), .B(new_n512), .C1(new_n360), .C2(new_n287), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT28), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n512), .B1(new_n360), .B2(new_n519), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n502), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n554), .B1(new_n532), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n546), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n539), .A2(new_n545), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(G472), .A2(G902), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT32), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n541), .A2(new_n547), .A3(new_n542), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n546), .B1(new_n544), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n532), .A2(new_n556), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n553), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n287), .B1(new_n336), .B2(new_n342), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n549), .B1(new_n568), .B2(new_n508), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n531), .A3(new_n551), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT28), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n536), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT29), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n565), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n531), .B1(new_n509), .B2(new_n514), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT28), .B1(new_n576), .B2(new_n564), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n577), .A2(KEYINPUT29), .A3(new_n536), .A4(new_n572), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n378), .ZN(new_n579));
  OAI21_X1  g393(.A(G472), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n559), .A2(KEYINPUT32), .A3(new_n560), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n563), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n413), .B1(G234), .B2(new_n378), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT73), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT22), .B(G137), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n585), .B(new_n586), .Z(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n473), .A2(new_n447), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT77), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT23), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n213), .B2(G128), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n279), .A2(KEYINPUT23), .A3(G119), .ZN(new_n593));
  INV_X1    g407(.A(G110), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n213), .A2(G128), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT76), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n279), .A2(G119), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT24), .B(G110), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n596), .B2(KEYINPUT76), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n590), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n596), .A2(KEYINPUT76), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n605), .A2(KEYINPUT77), .A3(new_n597), .A4(new_n602), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n589), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT78), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n473), .A2(new_n479), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n600), .A2(new_n601), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(G110), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT75), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n610), .A2(KEYINPUT75), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n607), .A2(new_n608), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n588), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n620), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n608), .A2(new_n607), .B1(new_n616), .B2(new_n617), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n587), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(new_n624), .A3(new_n378), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT25), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n584), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n621), .A2(new_n624), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n583), .A2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n501), .A2(new_n582), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  NAND2_X1  g450(.A1(KEYINPUT99), .A2(G472), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n559), .A2(new_n378), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n559), .B2(new_n378), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n319), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n361), .B1(new_n385), .B2(new_n371), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n365), .B1(new_n374), .B2(new_n360), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n642), .A2(new_n365), .B1(new_n643), .B2(new_n357), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n379), .B1(new_n644), .B2(G469), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n384), .A2(new_n386), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n377), .A3(new_n378), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n641), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n629), .A2(new_n648), .A3(new_n632), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n496), .A2(new_n499), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n418), .A2(new_n652), .A3(new_n420), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n416), .A2(KEYINPUT33), .A3(new_n417), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(G478), .A3(new_n378), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n421), .A2(new_n422), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n651), .A2(new_n200), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n314), .B1(new_n316), .B2(KEYINPUT100), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n292), .A2(new_n660), .A3(new_n310), .A4(new_n313), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n188), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n658), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n658), .B2(new_n662), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n650), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NAND2_X1  g482(.A1(new_n495), .A2(new_n486), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n499), .ZN(new_n670));
  INV_X1    g484(.A(new_n200), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n670), .A2(new_n424), .A3(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n662), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n650), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NAND2_X1  g490(.A1(new_n622), .A2(new_n623), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n588), .A2(KEYINPUT36), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n631), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n629), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n501), .A2(new_n640), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  XOR2_X1   g498(.A(new_n194), .B(KEYINPUT102), .Z(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n685), .B1(new_n686), .B2(new_n196), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n670), .A2(new_n424), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n582), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n662), .A2(new_n681), .A3(new_n648), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n279), .ZN(G30));
  XOR2_X1   g506(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n687), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n648), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT40), .Z(new_n696));
  NOR2_X1   g510(.A1(new_n315), .A2(new_n316), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT38), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n424), .A2(new_n188), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n699), .A2(new_n651), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n681), .ZN(new_n703));
  NAND2_X1  g517(.A1(G472), .A2(G902), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n546), .B1(new_n576), .B2(new_n564), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n544), .A2(new_n537), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n563), .A2(new_n710), .A3(new_n581), .A4(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n696), .A2(new_n702), .A3(new_n703), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  AOI221_X4 g528(.A(new_n687), .B1(new_n655), .B2(new_n656), .C1(new_n496), .C2(new_n499), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n582), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n690), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n271), .ZN(G48));
  NAND2_X1  g532(.A1(KEYINPUT105), .A2(G469), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n646), .B2(new_n378), .ZN(new_n720));
  INV_X1    g534(.A(new_n719), .ZN(new_n721));
  AOI211_X1 g535(.A(G902), .B(new_n721), .C1(new_n384), .C2(new_n386), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n722), .A3(new_n641), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n633), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n582), .B(new_n725), .C1(new_n664), .C2(new_n665), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND3_X1  g542(.A1(new_n673), .A2(new_n582), .A3(new_n725), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  INV_X1    g544(.A(new_n500), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n681), .A2(new_n731), .A3(new_n200), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n659), .A2(new_n661), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n733), .A2(new_n734), .A3(new_n189), .A4(new_n723), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n733), .B1(new_n662), .B2(new_n723), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n582), .B(new_n732), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  NOR4_X1   g552(.A1(new_n720), .A2(new_n722), .A3(new_n671), .A4(new_n641), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n700), .A2(new_n734), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(G472), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n559), .B2(new_n378), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n536), .B1(new_n577), .B2(new_n572), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n523), .B1(new_n522), .B2(new_n538), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n547), .B1(new_n541), .B2(new_n542), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n571), .B1(new_n747), .B2(new_n532), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n546), .B1(new_n748), .B2(new_n552), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT107), .A3(new_n545), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n746), .A2(new_n539), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n742), .B1(new_n751), .B2(new_n560), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n740), .A2(new_n634), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  NAND2_X1  g568(.A1(new_n750), .A2(new_n539), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT107), .B1(new_n749), .B2(new_n545), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n560), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n559), .A2(new_n378), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(G472), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n681), .A3(new_n715), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n662), .A2(new_n733), .A3(new_n723), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n734), .A2(new_n189), .A3(new_n723), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT106), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n760), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n276), .ZN(G27));
  INV_X1    g579(.A(new_n316), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n314), .A3(new_n189), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n388), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n582), .A2(new_n634), .A3(new_n715), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n687), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n651), .A2(new_n657), .A3(new_n772), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n773), .A2(new_n767), .A3(new_n388), .A4(new_n770), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n563), .A2(KEYINPUT108), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT32), .B1(new_n559), .B2(new_n560), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n580), .B(new_n581), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n774), .B(new_n634), .C1(new_n775), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n771), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT109), .B(G131), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G33));
  NAND4_X1  g596(.A1(new_n582), .A2(new_n634), .A3(new_n688), .A4(new_n768), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n644), .A2(KEYINPUT45), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT110), .Z(new_n786));
  NOR2_X1   g600(.A1(new_n644), .A2(KEYINPUT45), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n377), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n379), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(KEYINPUT46), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n647), .B1(new_n789), .B2(KEYINPUT46), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n319), .B(new_n694), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n651), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n657), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT43), .Z(new_n796));
  INV_X1    g610(.A(new_n640), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(new_n681), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n767), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n796), .A2(KEYINPUT44), .A3(new_n797), .A4(new_n681), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n793), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NOR4_X1   g618(.A1(new_n582), .A2(new_n634), .A3(new_n773), .A4(new_n767), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n319), .B1(new_n790), .B2(new_n791), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(KEYINPUT47), .B(new_n319), .C1(new_n790), .C2(new_n791), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n805), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  INV_X1    g626(.A(new_n808), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n720), .A2(new_n722), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n641), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n809), .A3(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n796), .A2(new_n685), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n752), .A2(new_n634), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n767), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n757), .A2(new_n681), .A3(new_n759), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n724), .A2(new_n767), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n801), .A2(new_n723), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n712), .A2(new_n826), .A3(new_n633), .A4(new_n194), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n794), .A3(new_n655), .A4(new_n656), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n824), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n825), .B2(new_n828), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n724), .B2(new_n189), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n723), .A2(KEYINPUT115), .A3(new_n188), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n698), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n819), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n831), .B1(new_n819), .B2(new_n835), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n830), .A2(new_n838), .A3(KEYINPUT118), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT118), .B1(new_n830), .B2(new_n838), .ZN(new_n840));
  OAI211_X1 g654(.A(KEYINPUT51), .B(new_n821), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n836), .A2(KEYINPUT116), .A3(new_n837), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n830), .A3(new_n821), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n778), .A2(new_n775), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n633), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n817), .A2(new_n849), .A3(new_n823), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT48), .Z(new_n851));
  NAND3_X1  g665(.A1(new_n827), .A2(new_n651), .A3(new_n657), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n763), .A2(new_n761), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n191), .B(new_n852), .C1(new_n819), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n841), .A2(new_n847), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n690), .B1(new_n689), .B2(new_n716), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n764), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n700), .A2(new_n734), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n648), .A2(new_n772), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n860), .A2(new_n703), .A3(new_n712), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT52), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n690), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n865), .B(new_n582), .C1(new_n688), .C2(new_n715), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n822), .B(new_n715), .C1(new_n735), .C2(new_n736), .ZN(new_n867));
  AND4_X1   g681(.A1(KEYINPUT52), .A2(new_n866), .A3(new_n867), .A4(new_n863), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT114), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n859), .A2(KEYINPUT52), .A3(new_n863), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n867), .A3(new_n863), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n752), .A2(new_n681), .A3(new_n715), .A4(new_n768), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n424), .A2(new_n499), .A3(new_n669), .A4(new_n772), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n767), .A2(new_n878), .A3(new_n388), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n582), .A2(new_n879), .A3(new_n681), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n783), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n657), .B1(new_n496), .B2(new_n499), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n731), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n317), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n640), .A2(new_n883), .A3(new_n649), .A4(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n885), .A2(new_n635), .A3(new_n682), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n780), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n726), .A2(new_n737), .A3(new_n729), .A4(new_n753), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT112), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n725), .A2(new_n582), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n891), .A2(new_n673), .B1(new_n818), .B2(new_n740), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(KEYINPUT112), .A3(new_n726), .A4(new_n737), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT113), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n887), .A2(new_n890), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n890), .A3(new_n893), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT113), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n876), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT53), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n870), .A2(new_n873), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n897), .A2(new_n900), .A3(new_n895), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n899), .A2(KEYINPUT54), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n888), .A2(new_n900), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n904), .A2(new_n887), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n901), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n898), .B2(new_n900), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n903), .B1(new_n909), .B2(KEYINPUT54), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n857), .A2(new_n910), .B1(G952), .B2(G953), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n634), .A2(new_n189), .A3(new_n319), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT111), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n814), .B(KEYINPUT49), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n698), .A2(new_n914), .ZN(new_n915));
  OR4_X1    g729(.A1(new_n712), .A2(new_n913), .A3(new_n795), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n916), .ZN(G75));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n897), .A2(new_n895), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n864), .A2(new_n868), .A3(KEYINPUT114), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n874), .B1(new_n870), .B2(new_n873), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n900), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n378), .B1(new_n923), .B2(new_n906), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n918), .B1(new_n924), .B2(new_n312), .ZN(new_n925));
  NOR4_X1   g739(.A1(new_n908), .A2(KEYINPUT119), .A3(new_n378), .A4(new_n313), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n260), .A2(new_n265), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n291), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n925), .A2(new_n926), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n190), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT56), .B1(new_n924), .B2(new_n312), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n929), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n932), .A2(new_n936), .ZN(G51));
  XNOR2_X1  g751(.A(new_n379), .B(KEYINPUT120), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT57), .Z(new_n939));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n908), .A2(new_n940), .ZN(new_n941));
  AOI211_X1 g755(.A(KEYINPUT54), .B(new_n907), .C1(new_n898), .C2(new_n900), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n646), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n924), .A2(new_n786), .A3(new_n788), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n933), .B1(new_n944), .B2(new_n945), .ZN(G54));
  NAND2_X1  g760(.A1(KEYINPUT58), .A2(G475), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n924), .A2(new_n491), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n491), .B1(new_n924), .B2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n933), .ZN(G60));
  NOR2_X1   g765(.A1(new_n941), .A2(new_n942), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT59), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n653), .A2(new_n654), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n934), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  AOI22_X1  g771(.A1(new_n910), .A2(new_n955), .B1(new_n653), .B2(new_n654), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n909), .A2(new_n679), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n630), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n908), .B2(new_n961), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n934), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n934), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G66));
  INV_X1    g784(.A(G224), .ZN(new_n971));
  OAI21_X1  g785(.A(G953), .B1(new_n197), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT121), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n890), .A2(new_n893), .A3(new_n886), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n975), .B2(G953), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n927), .B1(G898), .B2(new_n190), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G69));
  NOR2_X1   g792(.A1(new_n515), .A2(new_n521), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n465), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n859), .B(KEYINPUT122), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n713), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n984), .A3(new_n713), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n811), .A2(new_n803), .ZN(new_n986));
  INV_X1    g800(.A(new_n883), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n987), .A2(KEYINPUT123), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(KEYINPUT123), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n695), .A2(new_n767), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n582), .A3(new_n634), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n983), .A2(new_n985), .A3(new_n986), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n980), .B1(new_n993), .B2(new_n190), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n793), .A2(new_n860), .A3(new_n849), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n995), .A2(new_n780), .A3(new_n783), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n986), .A2(new_n981), .A3(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(G953), .ZN(new_n998));
  NAND2_X1  g812(.A1(G900), .A2(G953), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n980), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n994), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(G227), .ZN(new_n1002));
  OAI21_X1  g816(.A(G953), .B1(new_n1002), .B2(new_n686), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1001), .B(new_n1003), .ZN(G72));
  XOR2_X1   g818(.A(new_n704), .B(KEYINPUT63), .Z(new_n1005));
  OAI21_X1  g819(.A(new_n1005), .B1(new_n993), .B2(new_n974), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n522), .A2(new_n532), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT124), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1008), .A2(new_n546), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n997), .B2(new_n974), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n546), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT125), .Z(new_n1013));
  AOI21_X1  g827(.A(new_n933), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT126), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n707), .B1(new_n565), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1007), .A2(KEYINPUT126), .A3(new_n546), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n899), .A2(new_n902), .A3(new_n1005), .A4(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1010), .A2(new_n1014), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(KEYINPUT127), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT127), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1010), .A2(new_n1014), .A3(new_n1022), .A4(new_n1019), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(G57));
endmodule


