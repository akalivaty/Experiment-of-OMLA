//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(G355));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G116), .A2(G270), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT66), .B(G238), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n211), .B1(G68), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT67), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n214), .A2(new_n216), .B1(G1), .B2(G20), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G20), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n220), .B1(new_n221), .B2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n223), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n217), .A2(new_n218), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR4_X1   g0032(.A1(new_n219), .A2(new_n227), .A3(new_n228), .A4(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G232), .A3(G1698), .ZN(new_n255));
  AND3_X1   g0055(.A1(KEYINPUT75), .A2(G33), .A3(G97), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT75), .B1(G33), .B2(G97), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI211_X1 g0061(.A(G226), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n255), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n272), .A3(G274), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n268), .B(G274), .C1(G41), .C2(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT69), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n271), .A2(G238), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n267), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(new_n267), .B2(new_n276), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT14), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(G179), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n267), .A2(new_n276), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n267), .A2(new_n276), .A3(new_n277), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT14), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(G169), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT76), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(G68), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT12), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n203), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n230), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G77), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n230), .A2(new_n251), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n295), .B1(new_n296), .B2(new_n297), .C1(new_n201), .C2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n231), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT11), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(KEYINPUT11), .A3(new_n301), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n292), .A2(new_n231), .A3(new_n300), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n268), .A2(G20), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(G68), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT77), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT77), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n303), .B2(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n290), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n280), .A2(G190), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n287), .A2(G200), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(new_n310), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n254), .A2(G1698), .ZN(new_n322));
  INV_X1    g0122(.A(G223), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n322), .A2(new_n323), .B1(new_n297), .B2(new_n254), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n254), .A2(G222), .A3(new_n259), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n266), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n274), .B(new_n272), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(G226), .B2(new_n271), .ZN(new_n329));
  AOI21_X1  g0129(.A(G169), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT8), .B(G58), .ZN(new_n331));
  INV_X1    g0131(.A(G150), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n331), .A2(new_n296), .B1(new_n332), .B2(new_n298), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n204), .A2(G20), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(KEYINPUT70), .B(new_n301), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n201), .B1(new_n268), .B2(G20), .ZN(new_n337));
  INV_X1    g0137(.A(new_n292), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n306), .A2(new_n337), .B1(new_n201), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n334), .B1(new_n332), .B2(new_n298), .C1(new_n296), .C2(new_n331), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT70), .B1(new_n341), .B2(new_n301), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n330), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT71), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT71), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n330), .B2(new_n343), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n327), .A2(new_n329), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n345), .B(new_n347), .C1(G179), .C2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n254), .A2(G232), .A3(new_n259), .ZN(new_n350));
  INV_X1    g0150(.A(G107), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n350), .B1(new_n351), .B2(new_n254), .C1(new_n322), .C2(new_n212), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n266), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n328), .B1(G244), .B2(new_n271), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n353), .A2(KEYINPUT72), .A3(G190), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n301), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n356), .A2(G77), .A3(new_n292), .A4(new_n307), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G20), .A2(G77), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n360), .B1(new_n331), .B2(new_n298), .C1(new_n296), .C2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n301), .B1(new_n297), .B2(new_n338), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n355), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n353), .B2(new_n354), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT72), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n353), .A2(new_n354), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n366), .A2(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n368), .A2(new_n281), .B1(new_n359), .B2(new_n363), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n353), .A2(new_n372), .A3(new_n354), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n364), .A2(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n348), .A2(new_n369), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n365), .B1(new_n327), .B2(new_n329), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT9), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n343), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT9), .B1(new_n340), .B2(new_n342), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT74), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT10), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n377), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n377), .B2(new_n381), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n349), .B(new_n374), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n288), .B1(new_n280), .B2(G179), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n314), .B1(new_n389), .B2(new_n282), .ZN(new_n390));
  INV_X1    g0190(.A(new_n320), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT78), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT81), .ZN(new_n393));
  OAI211_X1 g0193(.A(G223), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n394));
  OAI211_X1 g0194(.A(G226), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n266), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n265), .A2(G232), .A3(new_n269), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT80), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n265), .A2(new_n269), .A3(KEYINPUT80), .A4(G232), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n273), .A2(new_n275), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n398), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n365), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n401), .A2(new_n402), .B1(new_n273), .B2(new_n275), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n369), .A3(new_n398), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n260), .A2(new_n261), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n410), .B2(new_n230), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n253), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(G68), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n202), .A2(new_n203), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G58), .A2(G68), .ZN(new_n416));
  OAI21_X1  g0216(.A(G20), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n230), .A2(new_n251), .A3(G159), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n356), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n252), .A2(new_n230), .A3(new_n253), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n203), .B1(new_n424), .B2(new_n412), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n417), .A2(new_n418), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n421), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n307), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n331), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n430), .A2(new_n305), .B1(new_n431), .B2(new_n292), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT79), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT79), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n434), .B1(new_n431), .B2(new_n292), .C1(new_n430), .C2(new_n305), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n420), .A2(new_n427), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n409), .A2(new_n436), .A3(KEYINPUT17), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT17), .B1(new_n409), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n393), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n405), .A2(new_n281), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n407), .A2(new_n372), .A3(new_n398), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n442), .A2(new_n436), .A3(KEYINPUT18), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n407), .A2(new_n372), .A3(new_n398), .ZN(new_n445));
  AOI21_X1  g0245(.A(G169), .B1(new_n407), .B2(new_n398), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n433), .A2(new_n435), .ZN(new_n448));
  INV_X1    g0248(.A(new_n426), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT16), .B1(new_n414), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n418), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n301), .B1(new_n425), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n448), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n444), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n443), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT17), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n407), .A2(new_n369), .A3(new_n398), .ZN(new_n457));
  AOI21_X1  g0257(.A(G200), .B1(new_n407), .B2(new_n398), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n456), .B1(new_n459), .B2(new_n453), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n409), .A2(new_n436), .A3(KEYINPUT17), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(KEYINPUT81), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n439), .A2(new_n455), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AND4_X1   g0264(.A1(new_n321), .A2(new_n387), .A3(new_n392), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(G41), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  INV_X1    g0272(.A(new_n231), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n470), .A2(new_n472), .B1(new_n473), .B2(new_n264), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n268), .A2(G45), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n468), .B2(new_n469), .ZN(new_n476));
  INV_X1    g0276(.A(G274), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n473), .B2(new_n264), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n474), .A2(G270), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G257), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n480));
  OAI211_X1 g0280(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n252), .A2(G303), .A3(new_n253), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n266), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n268), .A2(G33), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n306), .A2(G116), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n338), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n300), .A2(new_n231), .B1(G20), .B2(new_n488), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  INV_X1    g0291(.A(G97), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n491), .B(new_n230), .C1(G33), .C2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT20), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n490), .A2(KEYINPUT20), .A3(new_n493), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n487), .B(new_n489), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n485), .A2(new_n496), .A3(KEYINPUT21), .A4(G169), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT84), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n281), .B1(new_n479), .B2(new_n484), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(KEYINPUT84), .A3(KEYINPUT21), .A4(new_n496), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n496), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT21), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n479), .A2(G179), .A3(new_n484), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n496), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n496), .B1(new_n485), .B2(G200), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n369), .B2(new_n485), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n502), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n306), .A2(new_n486), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT25), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n292), .B2(G107), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n292), .A2(new_n513), .A3(G107), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT88), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(KEYINPUT88), .B(new_n513), .C1(new_n292), .C2(G107), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n512), .A2(G107), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n230), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT22), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n254), .A2(new_n523), .A3(new_n230), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n230), .A2(G33), .A3(G116), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT86), .B1(new_n528), .B2(KEYINPUT23), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n230), .A2(G107), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n526), .B(new_n527), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT85), .B1(new_n351), .B2(G20), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n532), .A2(KEYINPUT86), .A3(KEYINPUT23), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n525), .A2(new_n534), .A3(KEYINPUT87), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(KEYINPUT24), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT87), .B1(new_n525), .B2(new_n534), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n356), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n520), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n474), .A2(G264), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n476), .A2(new_n478), .ZN(new_n545));
  OAI211_X1 g0345(.A(G250), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G294), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n259), .B1(new_n252), .B2(new_n253), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(KEYINPUT89), .A3(G257), .ZN(new_n550));
  OAI211_X1 g0350(.A(G257), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT89), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n548), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n544), .B(new_n545), .C1(new_n554), .C2(new_n265), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n281), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n546), .A2(new_n547), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT89), .B1(new_n549), .B2(G257), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n551), .A2(new_n552), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n266), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n561), .A2(new_n372), .A3(new_n545), .A4(new_n544), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n543), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n555), .A2(new_n365), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n561), .A2(new_n369), .A3(new_n545), .A4(new_n544), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n543), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n265), .A2(G250), .A3(new_n475), .ZN(new_n569));
  OR2_X1    g0369(.A1(G238), .A2(G1698), .ZN(new_n570));
  INV_X1    g0370(.A(G244), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G1698), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n572), .C1(new_n260), .C2(new_n261), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G116), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n569), .B1(new_n575), .B2(new_n266), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT83), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n265), .A2(G274), .A3(new_n472), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT82), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n478), .A2(new_n580), .A3(new_n472), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n576), .A2(new_n577), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n577), .B1(new_n576), .B2(new_n582), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n281), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n254), .A2(new_n230), .A3(G68), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n296), .A2(new_n492), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(KEYINPUT19), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT19), .B1(new_n256), .B2(new_n257), .ZN(new_n589));
  INV_X1    g0389(.A(G87), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n589), .A2(new_n230), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n301), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n361), .A2(new_n338), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n594), .C1(new_n361), .C2(new_n511), .ZN(new_n595));
  INV_X1    g0395(.A(new_n569), .ZN(new_n596));
  NOR2_X1   g0396(.A1(G238), .A2(G1698), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n571), .B2(G1698), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n598), .A2(new_n254), .B1(G33), .B2(G116), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(new_n265), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n580), .B1(new_n478), .B2(new_n472), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n580), .A2(new_n265), .A3(G274), .A4(new_n472), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT83), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n576), .A2(new_n577), .A3(new_n582), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n372), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n585), .A2(new_n595), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(G200), .B1(new_n583), .B2(new_n584), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n512), .A2(G87), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n593), .A2(new_n594), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(G190), .A3(new_n605), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n298), .A2(new_n297), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT6), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n492), .A2(new_n351), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n591), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n351), .A2(KEYINPUT6), .A3(G97), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n613), .B1(new_n618), .B2(G20), .ZN(new_n619));
  OAI21_X1  g0419(.A(G107), .B1(new_n411), .B2(new_n413), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n301), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n292), .A2(G97), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n511), .B2(new_n492), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(G244), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT4), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n491), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n266), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n470), .A2(new_n472), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(G257), .A3(new_n265), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n545), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n634), .A2(new_n638), .A3(G179), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n281), .B1(new_n634), .B2(new_n638), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n627), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n625), .B1(new_n621), .B2(new_n301), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n634), .A2(new_n638), .A3(new_n369), .ZN(new_n643));
  AOI21_X1  g0443(.A(G200), .B1(new_n634), .B2(new_n638), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n607), .A2(new_n612), .A3(new_n641), .A4(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n465), .A2(new_n510), .A3(new_n568), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT90), .ZN(G372));
  INV_X1    g0449(.A(new_n349), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n371), .A2(new_n373), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n390), .B1(new_n320), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n439), .A2(new_n462), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n455), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n384), .A2(new_n385), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n465), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n502), .B(new_n506), .C1(new_n543), .C2(new_n563), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n641), .A2(new_n645), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n543), .A2(new_n567), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n576), .A2(new_n582), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G200), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n611), .A2(new_n610), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n281), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n606), .A2(new_n595), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT91), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n639), .B2(new_n640), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n634), .A2(new_n638), .A3(G179), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n637), .B1(new_n266), .B2(new_n633), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n670), .B(KEYINPUT91), .C1(new_n281), .C2(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n669), .A2(new_n627), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n667), .A2(new_n664), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT26), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n634), .A2(new_n638), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G169), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n642), .B1(new_n677), .B2(new_n670), .ZN(new_n678));
  AND4_X1   g0478(.A1(KEYINPUT26), .A2(new_n607), .A3(new_n612), .A4(new_n678), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n665), .B(new_n667), .C1(new_n675), .C2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n657), .B1(new_n658), .B2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n502), .A2(new_n506), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n268), .A2(new_n230), .A3(G13), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n525), .A2(new_n534), .A3(KEYINPUT87), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n693), .A2(new_n540), .A3(new_n541), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n301), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n519), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n556), .A2(new_n562), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n690), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n661), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n564), .A2(new_n690), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT92), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT92), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(new_n705), .A3(new_n702), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n692), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n699), .A2(new_n690), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT93), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n701), .A2(new_n705), .A3(new_n702), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n705), .B1(new_n701), .B2(new_n702), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n691), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  INV_X1    g0513(.A(new_n708), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n710), .A2(new_n711), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n496), .A2(new_n690), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n510), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n684), .B2(new_n718), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n716), .A2(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n225), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n591), .A2(new_n590), .A3(new_n488), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT94), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n726), .A2(new_n728), .A3(new_n268), .ZN(new_n729));
  INV_X1    g0529(.A(new_n229), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n726), .ZN(new_n731));
  XNOR2_X1  g0531(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  INV_X1    g0534(.A(new_n690), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n680), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n669), .A2(new_n627), .A3(new_n672), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n667), .A2(new_n664), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT26), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT26), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n607), .A2(new_n612), .A3(new_n678), .A4(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n665), .A2(new_n667), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n734), .B1(new_n742), .B2(new_n735), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n568), .A2(new_n647), .A3(new_n510), .A4(new_n735), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n671), .A2(new_n604), .A3(new_n605), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n505), .A2(new_n544), .A3(new_n561), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n583), .A2(new_n584), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n544), .B1(new_n554), .B2(new_n265), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n479), .A2(new_n484), .A3(G179), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n750), .A2(new_n753), .A3(KEYINPUT30), .A4(new_n671), .ZN(new_n754));
  AOI21_X1  g0554(.A(G179), .B1(new_n576), .B2(new_n582), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n676), .A2(new_n555), .A3(new_n485), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n749), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n690), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT31), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n745), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G330), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n744), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n733), .B1(new_n765), .B2(G1), .ZN(G364));
  INV_X1    g0566(.A(new_n721), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n230), .A2(G13), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT96), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(KEYINPUT97), .A3(new_n471), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n268), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT97), .B1(new_n769), .B2(new_n471), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n726), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G330), .B2(new_n720), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n231), .B1(G20), .B2(new_n281), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n725), .A2(new_n254), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(G45), .B2(new_n229), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G45), .B2(new_n248), .ZN(new_n784));
  NAND3_X1  g0584(.A1(G355), .A2(new_n225), .A3(new_n254), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G116), .B2(new_n225), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n781), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n774), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n230), .A2(G179), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n365), .A2(G190), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT100), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(KEYINPUT100), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n230), .A2(new_n372), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n796), .A2(KEYINPUT98), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT98), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n795), .A2(G107), .B1(G77), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n789), .A2(new_n797), .ZN(new_n803));
  INV_X1    g0603(.A(G159), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT101), .ZN(new_n808));
  AND3_X1   g0608(.A1(new_n796), .A2(new_n808), .A3(new_n790), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(new_n796), .B2(new_n790), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n802), .B(new_n807), .C1(new_n203), .C2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n789), .A2(G190), .A3(G200), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n796), .A2(G190), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n365), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n254), .B1(new_n590), .B2(new_n813), .C1(new_n816), .C2(new_n201), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n369), .A2(G179), .A3(G200), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n230), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n492), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n814), .A2(G200), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n202), .ZN(new_n823));
  NOR4_X1   g0623(.A1(new_n812), .A2(new_n817), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT102), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n821), .A2(G322), .ZN(new_n827));
  INV_X1    g0627(.A(new_n803), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n254), .B1(new_n828), .B2(G329), .ZN(new_n829));
  INV_X1    g0629(.A(G294), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n830), .B2(new_n819), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n827), .B(new_n831), .C1(G326), .C2(new_n815), .ZN(new_n832));
  INV_X1    g0632(.A(new_n813), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT103), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(KEYINPUT103), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G303), .B1(G311), .B2(new_n801), .ZN(new_n838));
  INV_X1    g0638(.A(new_n811), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT33), .B(G317), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n795), .A2(G283), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n832), .A2(new_n838), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n825), .A2(KEYINPUT102), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n826), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n788), .B1(new_n845), .B2(new_n780), .ZN(new_n846));
  INV_X1    g0646(.A(new_n779), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n720), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n776), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  NOR2_X1   g0650(.A1(new_n651), .A2(new_n690), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n359), .A2(new_n363), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n690), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n364), .B2(new_n370), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n852), .B1(new_n856), .B2(new_n652), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n681), .B2(new_n690), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n374), .A2(new_n735), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n675), .A2(new_n679), .ZN(new_n860));
  INV_X1    g0660(.A(new_n659), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n661), .A2(new_n641), .A3(new_n645), .A4(new_n664), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n667), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n859), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n774), .B1(new_n865), .B2(new_n763), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n763), .B2(new_n865), .ZN(new_n867));
  INV_X1    g0667(.A(new_n774), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n780), .A2(new_n777), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n297), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n837), .A2(G107), .B1(G283), .B2(new_n839), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n795), .A2(G87), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n871), .B(new_n872), .C1(new_n488), .C2(new_n800), .ZN(new_n873));
  INV_X1    g0673(.A(G311), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n410), .B1(new_n803), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(G303), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n822), .A2(new_n830), .B1(new_n816), .B2(new_n876), .ZN(new_n877));
  NOR4_X1   g0677(.A1(new_n873), .A2(new_n820), .A3(new_n875), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n795), .A2(G68), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n836), .B2(new_n201), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT104), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  INV_X1    g0683(.A(G132), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n254), .B1(new_n803), .B2(new_n884), .C1(new_n819), .C2(new_n202), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(G137), .A2(new_n815), .B1(new_n821), .B2(G143), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n887), .B1(new_n800), .B2(new_n804), .C1(new_n332), .C2(new_n811), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT34), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n878), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n780), .ZN(new_n891));
  INV_X1    g0691(.A(new_n857), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n870), .B1(new_n890), .B2(new_n891), .C1(new_n892), .C2(new_n778), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n867), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(G384));
  INV_X1    g0695(.A(KEYINPUT109), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n760), .A2(new_n761), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n699), .A2(new_n661), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n898), .A2(new_n646), .A3(new_n509), .A4(new_n690), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n745), .A2(KEYINPUT109), .A3(new_n760), .A4(new_n761), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n465), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT110), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n315), .A2(new_n690), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n316), .A2(new_n904), .A3(new_n320), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n315), .B(new_n690), .C1(new_n391), .C2(new_n290), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n857), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n900), .A2(new_n907), .A3(new_n901), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT106), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n447), .A2(new_n453), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n409), .A2(new_n436), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  INV_X1    g0712(.A(new_n688), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n453), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT105), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(KEYINPUT105), .A3(KEYINPUT37), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n914), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n463), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n921), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n909), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n921), .A2(new_n923), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n908), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT107), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n918), .A2(new_n933), .A3(new_n915), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n910), .A2(new_n911), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n935), .A2(KEYINPUT107), .A3(new_n912), .A4(new_n914), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT18), .B1(new_n442), .B2(new_n436), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n447), .A2(new_n444), .A3(new_n453), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n460), .A2(new_n937), .A3(new_n938), .A4(new_n461), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n922), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n934), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n928), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n930), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT40), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n932), .A2(KEYINPUT40), .B1(new_n908), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(G330), .B1(new_n903), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n903), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT111), .Z(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n926), .A2(new_n931), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n905), .A2(new_n906), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n864), .B2(new_n852), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT39), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n943), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n929), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n390), .A2(new_n735), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n688), .B1(new_n443), .B2(new_n454), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n953), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT108), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n953), .A2(KEYINPUT108), .A3(new_n959), .A4(new_n960), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n465), .B1(new_n736), .B2(new_n743), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n657), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n965), .B(new_n967), .Z(new_n968));
  AOI22_X1  g0768(.A1(new_n949), .A2(new_n968), .B1(G1), .B2(new_n769), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n949), .B2(new_n968), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n618), .A2(KEYINPUT35), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n618), .A2(KEYINPUT35), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n231), .A2(new_n230), .A3(new_n488), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT36), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n415), .A2(new_n229), .A3(new_n297), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n203), .A2(G50), .ZN(new_n977));
  OAI211_X1 g0777(.A(G1), .B(new_n223), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n970), .A2(new_n975), .A3(new_n978), .ZN(G367));
  NOR3_X1   g0779(.A1(new_n237), .A2(new_n725), .A3(new_n254), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n781), .B1(new_n225), .B2(new_n361), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n774), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n811), .A2(new_n804), .B1(new_n800), .B2(new_n201), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT115), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n819), .A2(new_n203), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(G143), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(new_n987), .B2(new_n816), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G150), .B2(new_n821), .ZN(new_n989));
  INV_X1    g0789(.A(G137), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n254), .B1(new_n803), .B2(new_n990), .C1(new_n202), .C2(new_n813), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n795), .B2(G77), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n983), .A2(KEYINPUT115), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n984), .A2(new_n989), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n837), .A2(KEYINPUT46), .A3(G116), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n813), .A2(new_n488), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(KEYINPUT46), .B2(new_n996), .C1(new_n830), .C2(new_n811), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT114), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n794), .A2(new_n492), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G303), .A2(new_n821), .B1(new_n815), .B2(G311), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n254), .B1(new_n828), .B2(G317), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n351), .C2(new_n819), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n999), .B(new_n1002), .C1(G283), .C2(new_n801), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n997), .A2(KEYINPUT114), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n994), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n982), .B1(new_n1007), .B2(new_n780), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n610), .A2(new_n735), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1009), .A2(new_n595), .A3(new_n606), .A4(new_n666), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n738), .B2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1008), .B1(new_n847), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n660), .B1(new_n642), .B2(new_n735), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n673), .A2(new_n690), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n707), .A2(KEYINPUT93), .A3(new_n708), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n716), .A2(KEYINPUT45), .A3(new_n1015), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1015), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n709), .A2(new_n715), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT44), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n709), .A2(KEYINPUT44), .A3(new_n715), .A4(new_n1023), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1022), .A2(new_n1028), .A3(new_n723), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n723), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n717), .B(new_n691), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(new_n767), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(new_n764), .ZN(new_n1034));
  AOI21_X1  g0834(.A(KEYINPUT113), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1027), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT45), .B1(new_n716), .B2(new_n1015), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1019), .B(new_n1023), .C1(new_n709), .C2(new_n715), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1036), .A2(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n722), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1022), .A2(new_n1028), .A3(new_n723), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1041), .A2(KEYINPUT113), .A3(new_n1042), .A4(new_n1034), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n765), .B1(new_n1035), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n726), .B(KEYINPUT41), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n773), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n707), .A2(new_n1015), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT42), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n641), .B1(new_n1023), .B2(new_n699), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1050), .B1(new_n735), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(KEYINPUT112), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT112), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1056), .A3(new_n1053), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n722), .A2(new_n1015), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n1052), .A2(new_n1053), .A3(new_n1061), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1058), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1060), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1012), .B1(new_n1048), .B2(new_n1066), .ZN(G387));
  NOR3_X1   g0867(.A1(new_n1034), .A2(G41), .A3(new_n725), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1033), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1068), .B1(new_n765), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n773), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n710), .A2(new_n711), .A3(new_n847), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n254), .B1(new_n828), .B2(G326), .ZN(new_n1073));
  INV_X1    g0873(.A(G283), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n819), .A2(new_n1074), .B1(new_n813), .B2(new_n830), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G317), .A2(new_n821), .B1(new_n815), .B2(G322), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n800), .B2(new_n876), .C1(new_n874), .C2(new_n811), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT49), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1073), .B1(new_n488), .B2(new_n794), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n819), .A2(new_n361), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G159), .B2(new_n815), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n201), .B2(new_n822), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n999), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n813), .A2(new_n297), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n410), .B(new_n1088), .C1(G150), .C2(new_n828), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n839), .A2(new_n431), .B1(new_n801), .B2(G68), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1082), .A2(new_n1083), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n780), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n241), .A2(new_n471), .A3(new_n254), .ZN(new_n1094));
  OR3_X1    g0894(.A1(new_n331), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT50), .B1(new_n331), .B2(G50), .ZN(new_n1096));
  AOI21_X1  g0896(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n728), .B1(new_n1098), .B2(new_n410), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(new_n725), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n781), .B1(new_n351), .B2(new_n225), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1093), .B(new_n774), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1070), .B1(new_n1071), .B2(new_n1033), .C1(new_n1072), .C2(new_n1103), .ZN(G393));
  NAND3_X1  g0904(.A1(new_n1041), .A2(new_n1042), .A3(new_n1034), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT113), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1043), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1108), .B(new_n726), .C1(new_n1031), .C2(new_n1034), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1110), .A2(KEYINPUT116), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1071), .B1(new_n1110), .B2(KEYINPUT116), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1015), .A2(new_n847), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT117), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G150), .A2(new_n815), .B1(new_n821), .B2(G159), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT51), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n872), .B1(new_n800), .B2(new_n331), .C1(new_n201), .C2(new_n811), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n819), .A2(new_n297), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n254), .B1(new_n803), .B2(new_n987), .C1(new_n203), .C2(new_n813), .ZN(new_n1119));
  OR4_X1    g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n410), .B1(new_n813), .B2(new_n1074), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G322), .B2(new_n828), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n830), .B2(new_n800), .C1(new_n794), .C2(new_n351), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT118), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n811), .A2(new_n876), .B1(new_n488), .B2(new_n819), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G311), .A2(new_n821), .B1(new_n815), .B2(G317), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT52), .Z(new_n1128));
  OAI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n891), .B1(new_n1120), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n781), .B1(new_n492), .B2(new_n225), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n245), .B2(new_n782), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1130), .A2(new_n868), .A3(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1111), .A2(new_n1112), .B1(new_n1114), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1109), .A2(new_n1134), .ZN(G390));
  OAI21_X1  g0935(.A(KEYINPUT119), .B1(new_n952), .B2(new_n958), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n955), .A2(new_n956), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT119), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n851), .B1(new_n680), .B2(new_n859), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1138), .B(new_n957), .C1(new_n1139), .C2(new_n951), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n856), .A2(new_n652), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n739), .A2(new_n741), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n735), .B(new_n1142), .C1(new_n863), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n852), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n951), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n943), .A3(new_n957), .ZN(new_n1148));
  INV_X1    g0948(.A(G330), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT31), .B1(new_n757), .B2(new_n690), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1149), .B(new_n857), .C1(new_n1152), .C2(new_n745), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1146), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1141), .A2(new_n1148), .A3(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n465), .A2(new_n900), .A3(G330), .A4(new_n901), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n966), .A2(new_n1156), .A3(new_n657), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n762), .A2(G330), .A3(new_n892), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n951), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n900), .A2(G330), .A3(new_n907), .A4(new_n901), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1139), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n900), .A2(G330), .A3(new_n892), .A4(new_n901), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n951), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1145), .B1(new_n1153), .B2(new_n1146), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1157), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n943), .A2(new_n957), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n957), .B1(new_n1139), .B2(new_n951), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(KEYINPUT119), .A2(new_n1171), .B1(new_n955), .B2(new_n956), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1170), .B1(new_n1172), .B2(new_n1140), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1155), .B(new_n1168), .C1(new_n1173), .C2(new_n1160), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1174), .A2(new_n726), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT120), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1157), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1141), .A2(new_n1148), .A3(new_n1154), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1160), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1176), .B(new_n1179), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1155), .B1(new_n1173), .B2(new_n1160), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1176), .B1(new_n1184), .B2(new_n1179), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1175), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1137), .A2(new_n777), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n837), .A2(G87), .B1(G97), .B2(new_n801), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n879), .C1(new_n351), .C2(new_n811), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n254), .B(new_n1118), .C1(G294), .C2(new_n828), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n488), .B2(new_n822), .C1(new_n1074), .C2(new_n816), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n813), .A2(new_n332), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1192), .A2(new_n1193), .B1(new_n815), .B2(G128), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n804), .B2(new_n819), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1195));
  XOR2_X1   g0995(.A(KEYINPUT54), .B(G143), .Z(new_n1196));
  AOI22_X1  g0996(.A1(new_n839), .A2(G137), .B1(new_n801), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(G125), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n254), .B1(new_n803), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G132), .B2(new_n821), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1197), .B(new_n1200), .C1(new_n201), .C2(new_n794), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1189), .A2(new_n1191), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1202), .A2(new_n780), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n868), .B(new_n1203), .C1(new_n331), .C2(new_n869), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT122), .Z(new_n1205));
  NAND2_X1  g1005(.A1(new_n1187), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1184), .B2(new_n1071), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1186), .A2(new_n1208), .ZN(G378));
  NOR2_X1   g1009(.A1(new_n343), .A2(new_n688), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n656), .A2(new_n349), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1211), .B1(new_n656), .B2(new_n349), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  OR3_X1    g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1216), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n908), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT40), .B1(new_n950), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(G330), .B1(new_n944), .B2(new_n908), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1220), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n943), .A2(KEYINPUT40), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1149), .B1(new_n1225), .B2(new_n1221), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n1219), .C1(KEYINPUT40), .C2(new_n932), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n965), .A2(new_n1228), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n963), .A2(new_n1224), .A3(new_n964), .A4(new_n1227), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n773), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n868), .B1(new_n201), .B2(new_n869), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n819), .A2(new_n332), .ZN(new_n1233));
  INV_X1    g1033(.A(G128), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n822), .A2(new_n1234), .B1(new_n816), .B2(new_n1198), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(new_n833), .C2(new_n1196), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n884), .B2(new_n811), .C1(new_n990), .C2(new_n800), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1238));
  AOI211_X1 g1038(.A(G33), .B(G41), .C1(new_n828), .C2(G124), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n794), .B2(new_n804), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1237), .B2(KEYINPUT59), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n795), .A2(G58), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n410), .A2(new_n467), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1243), .B(new_n1088), .C1(G283), .C2(new_n828), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n986), .B1(new_n816), .B2(new_n488), .C1(new_n351), .C2(new_n822), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n811), .A2(new_n492), .B1(new_n800), .B2(new_n361), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1238), .A2(new_n1241), .B1(KEYINPUT58), .B2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1243), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1248), .B2(KEYINPUT58), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1251), .A2(KEYINPUT123), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(KEYINPUT123), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1249), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1232), .B1(new_n891), .B2(new_n1254), .C1(new_n1219), .C2(new_n778), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1231), .A2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n965), .A2(new_n1228), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n963), .A2(new_n964), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT57), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(new_n1229), .A3(KEYINPUT57), .A4(new_n1230), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n726), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1256), .B1(new_n1261), .B2(new_n1263), .ZN(G375));
  INV_X1    g1064(.A(new_n1177), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1157), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n1047), .A3(new_n1179), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n951), .A2(new_n777), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n254), .B1(new_n803), .B2(new_n1234), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n816), .A2(new_n884), .B1(new_n201), .B2(new_n819), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(G137), .C2(new_n821), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n837), .A2(G159), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n839), .A2(new_n1196), .B1(new_n801), .B2(G150), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1271), .A2(new_n1242), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n837), .A2(G97), .B1(new_n795), .B2(G77), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n811), .A2(new_n488), .B1(new_n800), .B2(new_n351), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(KEYINPUT124), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(KEYINPUT124), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n822), .A2(new_n1074), .B1(new_n816), .B2(new_n830), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n410), .B1(new_n803), .B2(new_n876), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1279), .A2(new_n1084), .A3(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1275), .A2(new_n1277), .A3(new_n1278), .A4(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n891), .B1(new_n1274), .B2(new_n1282), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n868), .B(new_n1283), .C1(new_n203), .C2(new_n869), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1177), .A2(new_n773), .B1(new_n1268), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1267), .A2(new_n1285), .ZN(G381));
  XOR2_X1   g1086(.A(G375), .B(KEYINPUT125), .Z(new_n1287));
  INV_X1    g1087(.A(G390), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1185), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1182), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1207), .B1(new_n1290), .B2(new_n1175), .ZN(new_n1291));
  NOR4_X1   g1091(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1288), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  OR3_X1    g1093(.A1(new_n1287), .A2(G387), .A3(new_n1293), .ZN(G407));
  NAND2_X1  g1094(.A1(new_n689), .A2(G213), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1291), .A2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G407), .B(G213), .C1(new_n1287), .C2(new_n1297), .ZN(G409));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1266), .B1(new_n1300), .B2(new_n1168), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1265), .A2(KEYINPUT60), .A3(new_n1157), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n726), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1285), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n894), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(G384), .A3(new_n1285), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1296), .A2(G2897), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1305), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G378), .B(new_n1256), .C1(new_n1261), .C2(new_n1263), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1260), .A2(new_n1229), .A3(new_n1047), .A4(new_n1230), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(new_n1231), .A3(new_n1255), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1291), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1296), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1299), .B1(new_n1312), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1307), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT63), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(G387), .A2(new_n1288), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(G393), .B(new_n849), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1046), .B1(new_n1108), .B2(new_n765), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1065), .B1(new_n1324), .B2(new_n773), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n1012), .A3(G390), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1322), .A2(new_n1323), .A3(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1323), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1325), .A2(new_n1012), .A3(G390), .ZN(new_n1329));
  AOI21_X1  g1129(.A(G390), .B1(new_n1325), .B2(new_n1012), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1328), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1317), .A2(KEYINPUT63), .A3(new_n1319), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1321), .A2(new_n1327), .A3(new_n1331), .A4(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1327), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(new_n1295), .A3(new_n1319), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(KEYINPUT62), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1295), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1311), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1308), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1338), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1317), .A2(new_n1343), .A3(new_n1319), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1337), .A2(new_n1342), .A3(new_n1344), .A4(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1334), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1333), .A2(new_n1347), .ZN(G405));
  NAND2_X1  g1148(.A1(G375), .A2(new_n1291), .ZN(new_n1349));
  AND3_X1   g1149(.A1(new_n1349), .A2(new_n1313), .A3(new_n1307), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1307), .B1(new_n1349), .B2(new_n1313), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1334), .A2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1331), .A2(new_n1352), .A3(new_n1327), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(G402));
endmodule


