//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G20), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n212), .B1(new_n216), .B2(new_n217), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT67), .ZN(new_n247));
  OR2_X1    g0047(.A1(new_n247), .A2(KEYINPUT10), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n208), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n213), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n250), .B1(new_n206), .B2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n256), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n214), .B1(new_n208), .B2(G33), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n252), .B1(G50), .B2(new_n253), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  XOR2_X1   g0066(.A(new_n266), .B(KEYINPUT9), .Z(new_n267));
  OAI21_X1  g0067(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G274), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n272), .A2(new_n269), .A3(new_n219), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G222), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G223), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n279), .B1(new_n280), .B2(new_n277), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  AOI211_X1 g0083(.A(new_n271), .B(new_n273), .C1(new_n283), .C2(new_n272), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G190), .ZN(new_n285));
  INV_X1    g0085(.A(G200), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(new_n284), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n248), .B1(new_n267), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n247), .A2(KEYINPUT10), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  OAI211_X1 g0091(.A(G1), .B(G13), .C1(new_n257), .C2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G223), .A2(G1698), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n219), .B2(G1698), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n257), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT72), .A2(G33), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(KEYINPUT3), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n275), .A2(G33), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n294), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G87), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n292), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G179), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n292), .A2(G232), .A3(new_n268), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n304), .A2(KEYINPUT73), .A3(new_n270), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT73), .B1(new_n304), .B2(new_n270), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n270), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n302), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n259), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(G20), .B1(new_n314), .B2(new_n201), .ZN(new_n315));
  INV_X1    g0115(.A(G159), .ZN(new_n316));
  INV_X1    g0116(.A(new_n262), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(G20), .B1(new_n298), .B2(new_n299), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n313), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT72), .A2(G33), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT72), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n274), .B1(new_n324), .B2(KEYINPUT3), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT7), .B1(new_n325), .B2(G20), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n318), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT16), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT16), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT3), .B1(new_n296), .B2(new_n297), .ZN(new_n330));
  OAI211_X1 g0130(.A(KEYINPUT7), .B(new_n207), .C1(new_n330), .C2(new_n276), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n320), .B1(new_n277), .B2(G20), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n313), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n329), .B1(new_n333), .B2(new_n318), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n328), .A2(new_n250), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n256), .A2(new_n260), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n253), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n251), .B2(new_n336), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n312), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT18), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n338), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n265), .B1(new_n327), .B2(KEYINPUT16), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(new_n334), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n302), .A2(G190), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n307), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT74), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT74), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n307), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n286), .B1(new_n302), .B2(new_n310), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT17), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n344), .A2(new_n351), .A3(KEYINPUT17), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(KEYINPUT75), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT75), .ZN(new_n356));
  INV_X1    g0156(.A(new_n354), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n352), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n341), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n284), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n266), .C1(G169), .C2(new_n284), .ZN(new_n362));
  INV_X1    g0162(.A(G244), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n272), .A2(new_n269), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n277), .A2(G232), .A3(new_n278), .ZN(new_n365));
  INV_X1    g0165(.A(G107), .ZN(new_n366));
  INV_X1    g0166(.A(G238), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n365), .B1(new_n366), .B2(new_n277), .C1(new_n281), .C2(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n271), .B(new_n364), .C1(new_n368), .C2(new_n272), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n369), .A2(new_n360), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n251), .A2(G77), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n254), .A2(new_n317), .B1(new_n207), .B2(new_n280), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT15), .B(G87), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n258), .B2(new_n374), .ZN(new_n375));
  OAI221_X1 g0175(.A(new_n371), .B1(G77), .B2(new_n253), .C1(new_n265), .C2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n369), .B2(G169), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n369), .B2(G190), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n286), .B2(new_n369), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n290), .A2(new_n359), .A3(new_n362), .A4(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n258), .A2(G77), .B1(G20), .B2(new_n313), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n202), .B2(new_n317), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n385), .A2(new_n250), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n386), .A2(KEYINPUT11), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(KEYINPUT11), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT12), .B1(new_n253), .B2(G68), .ZN(new_n389));
  OR3_X1    g0189(.A1(new_n253), .A2(KEYINPUT12), .A3(G68), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n251), .A2(G68), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT71), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT14), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT13), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT69), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n299), .A2(new_n397), .A3(G226), .A4(new_n278), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n398), .A2(KEYINPUT68), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(KEYINPUT68), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n299), .A2(new_n397), .A3(G232), .A4(G1698), .ZN(new_n402));
  INV_X1    g0202(.A(G97), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n257), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n396), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n406), .B1(new_n399), .B2(new_n400), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT69), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n409), .A3(new_n272), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n272), .A2(new_n269), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n271), .B1(new_n411), .B2(G238), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n395), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n409), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n272), .B1(new_n408), .B2(KEYINPUT69), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n395), .B(new_n412), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n394), .B(G169), .C1(new_n413), .C2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(G179), .A3(new_n416), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n416), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n394), .B1(new_n423), .B2(G169), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n393), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n413), .A2(new_n417), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n392), .B1(new_n426), .B2(G190), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT70), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n423), .B2(G200), .ZN(new_n429));
  AOI211_X1 g0229(.A(KEYINPUT70), .B(new_n286), .C1(new_n420), .C2(new_n416), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n383), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT24), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n299), .A2(new_n397), .ZN(new_n435));
  INV_X1    g0235(.A(G87), .ZN(new_n436));
  OR4_X1    g0236(.A1(KEYINPUT22), .A2(new_n435), .A3(G20), .A4(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n298), .A2(new_n207), .A3(G87), .A4(new_n299), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT84), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT22), .B1(new_n438), .B2(KEYINPUT84), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT85), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(KEYINPUT85), .B(new_n437), .C1(new_n440), .C2(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n366), .A2(G20), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT23), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n296), .A2(new_n297), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G116), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n451), .B2(G20), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n434), .B1(new_n446), .B2(new_n453), .ZN(new_n454));
  AOI211_X1 g0254(.A(KEYINPUT24), .B(new_n452), .C1(new_n444), .C2(new_n445), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n250), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT86), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n366), .B1(new_n457), .B2(KEYINPUT25), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n253), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n457), .B2(KEYINPUT25), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n457), .A3(KEYINPUT25), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT77), .B1(new_n257), .B2(G1), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT77), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n206), .A3(G33), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n465), .A3(new_n253), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n250), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n461), .A2(new_n462), .B1(new_n467), .B2(G107), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n473), .A2(G264), .A3(new_n292), .ZN(new_n474));
  MUX2_X1   g0274(.A(G250), .B(G257), .S(G1698), .Z(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(new_n298), .A3(new_n299), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n450), .A2(G294), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n478), .B2(new_n272), .ZN(new_n479));
  INV_X1    g0279(.A(G274), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n473), .A2(new_n272), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G190), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(G200), .B2(new_n483), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n456), .A2(new_n468), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n331), .A2(new_n332), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n366), .A2(KEYINPUT6), .A3(G97), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n403), .A2(new_n366), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n490), .B1(new_n493), .B2(KEYINPUT6), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n265), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n253), .A2(G97), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT76), .ZN(new_n498));
  INV_X1    g0298(.A(new_n467), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n403), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n277), .A2(G250), .A3(G1698), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n363), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(new_n278), .A3(new_n299), .A4(new_n397), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n298), .A2(G244), .A3(new_n278), .A4(new_n299), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n508), .A2(KEYINPUT78), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n503), .B1(new_n508), .B2(KEYINPUT78), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n272), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n473), .A2(new_n292), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n481), .B1(new_n514), .B2(G257), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n512), .A2(new_n360), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT78), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n325), .A2(new_n517), .A3(G244), .A4(new_n278), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n508), .A2(KEYINPUT78), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n503), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n292), .B1(new_n520), .B2(new_n507), .ZN(new_n521));
  INV_X1    g0321(.A(new_n515), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n309), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n501), .A2(new_n516), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n512), .A2(G190), .A3(new_n515), .ZN(new_n525));
  OAI21_X1  g0325(.A(G200), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n496), .A2(new_n500), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n525), .A2(new_n526), .A3(new_n530), .A4(new_n527), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n524), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n487), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(G264), .A2(G1698), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n298), .A2(new_n299), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT82), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n298), .A2(new_n537), .A3(new_n299), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n435), .A2(G303), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n298), .A2(G257), .A3(new_n278), .A4(new_n299), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT81), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n325), .A2(KEYINPUT81), .A3(G257), .A4(new_n278), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n539), .A2(new_n540), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n272), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n482), .B1(new_n221), .B2(new_n513), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n253), .A2(G116), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n467), .B2(G116), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n506), .B(new_n207), .C1(G33), .C2(new_n403), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n250), .B(new_n552), .C1(new_n207), .C2(G116), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT20), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n549), .A2(KEYINPUT21), .A3(G169), .A4(new_n557), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n360), .B(new_n547), .C1(new_n545), .C2(new_n272), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n557), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT83), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n558), .A2(new_n560), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT83), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(G169), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n547), .B1(new_n545), .B2(new_n272), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n557), .B1(new_n549), .B2(G200), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n484), .B2(new_n549), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n562), .A2(new_n564), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n374), .A2(new_n253), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n298), .A2(new_n207), .A3(G68), .A4(new_n299), .ZN(new_n573));
  XNOR2_X1  g0373(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n258), .A2(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(G20), .B1(new_n574), .B2(new_n404), .ZN(new_n578));
  NOR3_X1   g0378(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n573), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n572), .B1(new_n580), .B2(new_n250), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n373), .B2(new_n499), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n206), .A2(G45), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G250), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n272), .A2(new_n584), .B1(new_n480), .B2(new_n583), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n324), .A2(new_n220), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G238), .A2(G1698), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n363), .B2(G1698), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n587), .B1(new_n325), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n586), .B1(new_n590), .B2(new_n292), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n309), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n298), .A3(new_n299), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n451), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n585), .B1(new_n594), .B2(new_n272), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n360), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n582), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n591), .A2(G200), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(G190), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n467), .A2(G87), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n598), .A2(new_n581), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n456), .A2(new_n468), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n483), .A2(G169), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n360), .B2(new_n483), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n433), .A2(new_n533), .A3(new_n571), .A4(new_n606), .ZN(G372));
  NAND2_X1  g0407(.A1(new_n431), .A2(new_n378), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n425), .B1(new_n358), .B2(new_n355), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n290), .B1(new_n609), .B2(new_n341), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n610), .A2(new_n362), .ZN(new_n611));
  INV_X1    g0411(.A(new_n445), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT84), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n325), .A2(new_n613), .A3(new_n207), .A4(G87), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(KEYINPUT22), .A3(new_n439), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT85), .B1(new_n615), .B2(new_n437), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n453), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT24), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n446), .A2(new_n434), .A3(new_n453), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n265), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n468), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n605), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n568), .A2(new_n558), .A3(new_n560), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n598), .A2(new_n599), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n581), .A2(KEYINPUT87), .A3(new_n600), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT87), .B1(new_n581), .B2(new_n600), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n629), .A2(new_n597), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n625), .A2(new_n532), .A3(new_n487), .A4(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n597), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n597), .A2(new_n601), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n524), .A2(new_n633), .A3(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n512), .A2(new_n515), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n527), .B1(new_n635), .B2(new_n309), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n636), .A2(new_n516), .A3(new_n629), .A4(new_n597), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n634), .A2(KEYINPUT88), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n524), .A2(new_n640), .A3(KEYINPUT26), .A4(new_n633), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n632), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n631), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n433), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n611), .A2(new_n644), .ZN(G369));
  INV_X1    g0445(.A(G330), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n207), .A2(G13), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n206), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT89), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT27), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(G213), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n557), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n571), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n656), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n623), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n646), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n603), .A2(new_n655), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n661), .A2(new_n487), .B1(new_n603), .B2(new_n605), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n622), .A2(new_n655), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n660), .A2(KEYINPUT90), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT90), .B1(new_n660), .B2(new_n664), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n661), .A2(new_n487), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n622), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n564), .A2(new_n562), .A3(new_n568), .ZN(new_n671));
  INV_X1    g0471(.A(new_n655), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n663), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n668), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n210), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n579), .A2(new_n220), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n217), .B2(new_n679), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n533), .A2(new_n571), .A3(new_n606), .A4(new_n672), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n479), .A2(new_n595), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n521), .A2(new_n687), .A3(new_n522), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n559), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n546), .A2(G179), .A3(new_n548), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(KEYINPUT91), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n686), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT30), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n686), .B(new_n695), .C1(new_n690), .C2(new_n692), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n591), .A2(new_n360), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n483), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n635), .A2(new_n549), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n694), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n700), .A2(new_n701), .A3(new_n655), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n700), .B2(new_n655), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n685), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n655), .B1(new_n631), .B2(new_n642), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n622), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n533), .B(new_n630), .C1(new_n709), .C2(new_n671), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n501), .A2(new_n516), .A3(new_n523), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n711), .A2(new_n602), .A3(KEYINPUT26), .ZN(new_n712));
  AOI211_X1 g0512(.A(new_n632), .B(new_n712), .C1(KEYINPUT26), .C2(new_n637), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n655), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n705), .B(new_n708), .C1(new_n707), .C2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n684), .B1(new_n716), .B2(G1), .ZN(G364));
  AOI21_X1  g0517(.A(new_n206), .B1(new_n647), .B2(G45), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n678), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n660), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n561), .B1(new_n558), .B2(new_n560), .ZN(new_n723));
  INV_X1    g0523(.A(new_n568), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n570), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n659), .B1(new_n726), .B2(new_n658), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n721), .B1(G330), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n720), .B(KEYINPUT93), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n210), .A2(new_n277), .ZN(new_n730));
  INV_X1    g0530(.A(G355), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(G116), .B2(new_n210), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n677), .A2(new_n325), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n217), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n734), .B1(new_n469), .B2(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n242), .A2(new_n469), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n732), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n213), .B1(G20), .B2(new_n309), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n729), .B1(new_n738), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n207), .A2(new_n484), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n360), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n207), .A2(G190), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n747), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G322), .A2(new_n749), .B1(new_n752), .B2(G311), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n360), .A2(new_n286), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n750), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(KEYINPUT33), .B(G317), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n756), .A2(new_n757), .B1(new_n760), .B2(G329), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n753), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n286), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n750), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n277), .B(new_n762), .C1(G283), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n758), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G294), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n746), .A2(new_n754), .ZN(new_n771));
  INV_X1    g0571(.A(G326), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT94), .ZN(new_n774));
  INV_X1    g0574(.A(G303), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n746), .A2(new_n763), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT95), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(KEYINPUT95), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n766), .B(new_n774), .C1(new_n775), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n764), .A2(new_n366), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n277), .B1(new_n748), .B2(new_n259), .ZN(new_n782));
  INV_X1    g0582(.A(new_n776), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n781), .B(new_n782), .C1(G87), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n768), .A2(G97), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n759), .A2(new_n316), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n755), .A2(new_n313), .B1(new_n751), .B2(new_n280), .ZN(new_n788));
  INV_X1    g0588(.A(new_n771), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(G50), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n780), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n745), .B1(new_n792), .B2(new_n742), .ZN(new_n793));
  INV_X1    g0593(.A(new_n741), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n727), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n728), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n379), .A2(KEYINPUT100), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT100), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n378), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n801), .A2(new_n381), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n487), .A2(new_n532), .A3(new_n630), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n623), .B1(new_n603), .B2(new_n605), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n634), .A2(KEYINPUT88), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n637), .A2(new_n638), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n806), .A2(new_n641), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n597), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n802), .B(new_n672), .C1(new_n805), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n655), .A2(new_n376), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n798), .A2(new_n381), .A3(new_n811), .A4(new_n800), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n378), .A2(new_n655), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n810), .B1(new_n706), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n720), .B1(new_n815), .B2(new_n705), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n705), .B2(new_n815), .ZN(new_n817));
  INV_X1    g0617(.A(new_n742), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n435), .B1(new_n779), .B2(new_n366), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT96), .Z(new_n820));
  NOR2_X1   g0620(.A1(new_n764), .A2(new_n436), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G311), .B2(new_n760), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n822), .B1(new_n770), .B2(new_n748), .C1(new_n775), .C2(new_n771), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n785), .B1(new_n220), .B2(new_n751), .C1(new_n824), .C2(new_n755), .ZN(new_n825));
  OR3_X1    g0625(.A1(new_n820), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  INV_X1    g0627(.A(G150), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n771), .A2(new_n827), .B1(new_n755), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT97), .Z(new_n830));
  INV_X1    g0630(.A(G143), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n831), .B2(new_n748), .C1(new_n316), .C2(new_n751), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT34), .Z(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n325), .B1(new_n834), .B2(new_n759), .C1(new_n769), .C2(new_n259), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n779), .A2(new_n202), .B1(new_n313), .B2(new_n764), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(KEYINPUT98), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(KEYINPUT98), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n826), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT99), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n818), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  INV_X1    g0642(.A(new_n729), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n742), .A2(new_n739), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(new_n280), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n842), .B(new_n845), .C1(new_n740), .C2(new_n814), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n817), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  NOR2_X1   g0648(.A1(new_n647), .A2(new_n206), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n708), .B1(new_n714), .B2(new_n707), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n433), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n851), .A2(new_n611), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n335), .A2(new_n338), .ZN(new_n854));
  INV_X1    g0654(.A(new_n653), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n344), .A2(new_n351), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(new_n344), .C2(new_n312), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n339), .B(KEYINPUT18), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n357), .A2(new_n352), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n853), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n857), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n343), .B1(KEYINPUT16), .B2(new_n327), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n866), .A2(new_n338), .B1(new_n312), .B2(new_n653), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n858), .B2(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n338), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n855), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT38), .B(new_n869), .C1(new_n359), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n869), .B1(new_n359), .B2(new_n871), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n853), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n425), .A2(new_n655), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n875), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n801), .A2(new_n655), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n810), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n877), .A2(new_n872), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n393), .A2(new_n655), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n432), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n425), .A2(new_n431), .A3(new_n886), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n884), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n341), .A2(new_n653), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n881), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n852), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n433), .A2(new_n704), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT101), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n888), .A2(new_n889), .B1(new_n813), .B2(new_n812), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n704), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n864), .B2(new_n872), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n885), .A2(new_n704), .A3(new_n897), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n898), .A2(new_n900), .B1(new_n901), .B2(new_n899), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n646), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n896), .B2(new_n902), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n849), .B1(new_n894), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n894), .B2(new_n904), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n908));
  NOR4_X1   g0708(.A1(new_n907), .A2(new_n908), .A3(new_n216), .A4(new_n220), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT36), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n735), .B(G77), .C1(new_n259), .C2(new_n313), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n202), .A2(G68), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n206), .B(G13), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n906), .A2(new_n914), .ZN(G367));
  OR2_X1    g0715(.A1(new_n627), .A2(new_n628), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n630), .B1(new_n916), .B2(new_n672), .ZN(new_n917));
  OR3_X1    g0717(.A1(new_n916), .A2(new_n672), .A3(new_n597), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT43), .B1(new_n919), .B2(KEYINPUT102), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT102), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n917), .A2(new_n922), .A3(new_n918), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n921), .B1(new_n920), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT104), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n926), .A2(new_n927), .B1(KEYINPUT43), .B2(new_n919), .ZN(new_n928));
  INV_X1    g0728(.A(new_n663), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n670), .A2(new_n929), .A3(new_n674), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n532), .B1(new_n527), .B2(new_n672), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n524), .A2(new_n655), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT42), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT42), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n664), .A2(new_n936), .A3(new_n674), .A4(new_n933), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n529), .A2(new_n531), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n711), .B1(new_n622), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n672), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n935), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n928), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n667), .A2(new_n933), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n926), .A2(new_n927), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n928), .A2(new_n667), .A3(new_n933), .A4(new_n941), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n678), .B(KEYINPUT41), .Z(new_n950));
  INV_X1    g0750(.A(KEYINPUT45), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n929), .B(new_n933), .C1(new_n662), .C2(new_n673), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(KEYINPUT105), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(KEYINPUT105), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT105), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n675), .A2(new_n956), .A3(new_n933), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n952), .A2(KEYINPUT105), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n957), .A2(KEYINPUT45), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT44), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n675), .B2(new_n933), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n929), .B1(new_n662), .B2(new_n673), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(KEYINPUT44), .A3(new_n934), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n955), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n667), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n668), .A2(new_n955), .A3(new_n959), .A4(new_n964), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n727), .A2(G330), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n673), .B1(new_n662), .B2(new_n663), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(KEYINPUT106), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n968), .B1(KEYINPUT106), .B2(new_n969), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n930), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n969), .A2(KEYINPUT106), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n660), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n975), .A2(new_n664), .A3(new_n674), .A4(new_n970), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n715), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n966), .A2(new_n967), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n950), .B1(new_n978), .B2(new_n716), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n949), .B1(new_n979), .B2(new_n719), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n743), .B1(new_n210), .B2(new_n373), .C1(new_n734), .C2(new_n238), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n729), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT46), .B1(new_n783), .B2(G116), .ZN(new_n983));
  INV_X1    g0783(.A(new_n325), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n770), .B2(new_n755), .C1(new_n775), .C2(new_n748), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(G107), .C2(new_n768), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n765), .A2(G97), .ZN(new_n987));
  INV_X1    g0787(.A(G311), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n988), .B2(new_n771), .ZN(new_n989));
  INV_X1    g0789(.A(G317), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n751), .A2(new_n824), .B1(new_n759), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(KEYINPUT46), .A2(G116), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n986), .B(new_n992), .C1(new_n779), .C2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT107), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n771), .A2(new_n831), .B1(new_n776), .B2(new_n259), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n435), .B(new_n996), .C1(G150), .C2(new_n749), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n764), .A2(new_n280), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n755), .A2(new_n316), .B1(new_n751), .B2(new_n202), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(G137), .C2(new_n760), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n768), .A2(G68), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT108), .Z(new_n1003));
  NAND2_X1  g0803(.A1(new_n995), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT109), .Z(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n982), .B1(new_n794), .B2(new_n919), .C1(new_n1006), .C2(new_n818), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n980), .A2(new_n1007), .ZN(G387));
  NOR2_X1   g0808(.A1(new_n977), .A2(new_n679), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n973), .A2(new_n976), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n716), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n719), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n783), .A2(G294), .B1(new_n768), .B2(G283), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G322), .A2(new_n789), .B1(new_n756), .B2(G311), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n775), .B2(new_n751), .C1(new_n990), .C2(new_n748), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT48), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n1016), .B2(new_n1015), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT49), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n764), .A2(new_n220), .B1(new_n759), .B2(new_n772), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1019), .A2(new_n325), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n783), .A2(G77), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n374), .A2(new_n768), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1022), .A2(new_n987), .A3(new_n325), .A4(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n336), .A2(new_n755), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n771), .A2(new_n316), .B1(new_n751), .B2(new_n313), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n748), .A2(new_n202), .B1(new_n759), .B2(new_n828), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n742), .B1(new_n1021), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n235), .A2(new_n469), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n254), .A2(G50), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT50), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(G45), .B(new_n680), .C1(G68), .C2(G77), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n734), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1030), .B1(new_n1036), .B2(KEYINPUT110), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(KEYINPUT110), .B2(new_n1036), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(G107), .B2(new_n210), .C1(new_n681), .C2(new_n730), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n843), .B1(new_n1039), .B2(new_n743), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1029), .B(new_n1040), .C1(new_n664), .C2(new_n794), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1012), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1011), .A2(new_n1042), .ZN(G393));
  NAND2_X1  g0843(.A1(new_n966), .A2(new_n967), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n934), .A2(new_n741), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n743), .B1(new_n403), .B2(new_n210), .C1(new_n734), .C2(new_n245), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n729), .A2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n771), .A2(new_n990), .B1(new_n748), .B2(new_n988), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G303), .A2(new_n756), .B1(new_n752), .B2(G294), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G283), .A2(new_n783), .B1(new_n760), .B2(G322), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n277), .B(new_n781), .C1(G116), .C2(new_n768), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n821), .B(new_n984), .C1(G143), .C2(new_n760), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n756), .A2(G50), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n313), .B2(new_n776), .C1(new_n254), .C2(new_n751), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n768), .A2(G77), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1055), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n771), .A2(new_n828), .B1(new_n748), .B2(new_n316), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT51), .Z(new_n1062));
  OAI21_X1  g0862(.A(new_n1054), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1048), .B1(new_n1063), .B2(new_n742), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1045), .A2(new_n719), .B1(new_n1046), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n977), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1044), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n678), .A3(new_n978), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n1068), .ZN(G390));
  INV_X1    g0869(.A(KEYINPUT111), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n425), .A2(new_n431), .A3(new_n886), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n886), .B1(new_n425), .B2(new_n431), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n810), .B2(new_n883), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1070), .B1(new_n1074), .B2(new_n880), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n882), .B1(new_n706), .B2(new_n802), .ZN(new_n1076));
  OAI211_X1 g0876(.A(KEYINPUT111), .B(new_n879), .C1(new_n1076), .C2(new_n1073), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n875), .A2(new_n878), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n882), .B1(new_n714), .B2(new_n802), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n879), .B(new_n873), .C1(new_n1080), .C2(new_n1073), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n704), .A2(G330), .A3(new_n814), .A4(new_n890), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1079), .A2(new_n1083), .A3(new_n1081), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n719), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n843), .B1(new_n336), .B2(new_n844), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT113), .Z(new_n1089));
  OAI21_X1  g0889(.A(new_n277), .B1(new_n748), .B2(new_n834), .ZN(new_n1090));
  INV_X1    g0890(.A(G128), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n771), .A2(new_n1091), .B1(new_n755), .B2(new_n827), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(G159), .C2(new_n768), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n776), .A2(new_n828), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT54), .B(G143), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n202), .A2(new_n764), .B1(new_n751), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G125), .B2(new_n760), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1093), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n771), .A2(new_n824), .B1(new_n755), .B2(new_n366), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n277), .B(new_n1100), .C1(G68), .C2(new_n765), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1059), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G97), .A2(new_n752), .B1(new_n760), .B2(G294), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n220), .B2(new_n748), .C1(new_n779), .C2(new_n436), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1099), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n742), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1089), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT114), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1078), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n740), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1087), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n479), .A2(new_n595), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n512), .A2(new_n1113), .A3(new_n515), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(KEYINPUT91), .B2(new_n691), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n559), .A2(new_n689), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT92), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n699), .B1(new_n1117), .B2(new_n695), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n696), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n655), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT31), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n700), .A2(new_n701), .A3(new_n655), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n646), .B1(new_n1123), .B2(new_n685), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n433), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n851), .A2(new_n611), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n704), .A2(G330), .A3(new_n814), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1073), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1128), .A2(new_n1080), .A3(KEYINPUT112), .A4(new_n1083), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT112), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1076), .B1(new_n1128), .B2(new_n1083), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1126), .B(new_n1129), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n679), .B1(new_n1112), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1129), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n890), .B1(new_n1124), .B2(new_n814), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n884), .B1(new_n1138), .B2(new_n1084), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1136), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1140), .A2(new_n1085), .A3(new_n1086), .A4(new_n1126), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1111), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(G378));
  INV_X1    g0943(.A(KEYINPUT57), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1126), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1079), .A2(new_n1083), .A3(new_n1081), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1083), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1145), .B1(new_n1148), .B2(new_n1140), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n898), .A2(new_n900), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n901), .A2(new_n899), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n893), .B1(new_n1152), .B2(new_n646), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT117), .ZN(new_n1154));
  XOR2_X1   g0954(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n290), .A2(new_n362), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n266), .A3(new_n855), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT116), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n855), .A2(new_n266), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n290), .A2(new_n362), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1159), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1156), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1155), .A3(new_n1162), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1154), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n881), .A2(new_n891), .A3(new_n892), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n902), .A2(new_n1169), .A3(G330), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1153), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1168), .B1(new_n1153), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1144), .B1(new_n1149), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1168), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n902), .A2(new_n1169), .A3(G330), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1169), .B1(new_n902), .B2(G330), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1153), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1134), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(KEYINPUT57), .C1(new_n1181), .C2(new_n1145), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1174), .A2(new_n678), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n718), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n739), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G77), .A2(new_n783), .B1(new_n752), .B2(new_n374), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n765), .A2(G58), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n749), .A2(G107), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n1001), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G97), .A2(new_n756), .B1(new_n760), .B2(G283), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n220), .B2(new_n771), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n984), .A2(new_n291), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT115), .B(KEYINPUT58), .Z(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1193), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G125), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n771), .A2(new_n1200), .B1(new_n755), .B2(new_n834), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1096), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n783), .A2(new_n1202), .B1(new_n752), .B2(G137), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1091), .B2(new_n748), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1201), .B(new_n1204), .C1(G150), .C2(new_n768), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n765), .A2(G159), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n760), .C2(G124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1199), .B1(new_n1196), .B2(new_n1194), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n742), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n719), .B(new_n678), .C1(new_n202), .C2(new_n844), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1186), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1184), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1183), .A2(new_n1217), .ZN(G375));
  OAI21_X1  g1018(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1145), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n950), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(new_n1221), .A3(new_n1134), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT118), .Z(new_n1223));
  NAND2_X1  g1023(.A1(new_n1073), .A2(new_n739), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n742), .A2(G68), .A3(new_n739), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n789), .A2(G132), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT119), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n777), .A2(G159), .A3(new_n778), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n752), .A2(G150), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G137), .A2(new_n749), .B1(new_n760), .B2(G128), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n756), .A2(new_n1202), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n768), .A2(G50), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1232), .A2(new_n1188), .A3(new_n1233), .A4(new_n325), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G294), .A2(new_n789), .B1(new_n756), .B2(G116), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n998), .A2(new_n277), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1023), .A3(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G107), .A2(new_n752), .B1(new_n760), .B2(G303), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n824), .B2(new_n748), .C1(new_n779), .C2(new_n403), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1231), .A2(new_n1234), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1225), .B(new_n843), .C1(new_n742), .C2(new_n1240), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1140), .A2(new_n719), .B1(new_n1224), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1223), .A2(new_n1242), .ZN(G381));
  AND2_X1   g1043(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n847), .A3(new_n1245), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(G381), .A2(G387), .A3(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT120), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1217), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1141), .A2(new_n1126), .B1(new_n1179), .B2(new_n1178), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n679), .B1(new_n1250), .B2(KEYINPUT57), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1249), .B1(new_n1251), .B2(new_n1174), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1142), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1248), .A2(new_n1253), .ZN(G407));
  OAI211_X1 g1054(.A(G407), .B(G213), .C1(G343), .C2(new_n1253), .ZN(G409));
  INV_X1    g1055(.A(KEYINPUT127), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT125), .B1(G387), .B2(new_n1244), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n796), .B1(new_n1011), .B2(new_n1042), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1245), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(G390), .A2(new_n980), .A3(new_n1007), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G390), .B1(new_n980), .B2(new_n1007), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n1257), .A2(new_n1260), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G387), .A2(new_n1244), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1265), .A2(KEYINPUT125), .A3(new_n1261), .A4(new_n1259), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1264), .A2(KEYINPUT126), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT126), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1142), .B1(new_n1183), .B2(new_n1217), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT121), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1184), .B2(new_n1216), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n719), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(KEYINPUT121), .A3(new_n1215), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1180), .B(new_n1221), .C1(new_n1181), .C2(new_n1145), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1142), .A2(new_n1273), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n654), .A2(G213), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1271), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1139), .A2(new_n1131), .A3(new_n1130), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1126), .B1(new_n1281), .B2(new_n1129), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(KEYINPUT60), .B2(new_n1134), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1219), .A2(KEYINPUT60), .A3(new_n1145), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n678), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G384), .B(new_n1242), .C1(new_n1283), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT122), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1134), .A2(KEYINPUT60), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1220), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n678), .A3(new_n1284), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1291), .A2(KEYINPUT122), .A3(G384), .A4(new_n1242), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1242), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n847), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1288), .A2(new_n1292), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1270), .B1(new_n1280), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1288), .A2(new_n1292), .A3(new_n1294), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(new_n1271), .A2(new_n1279), .A3(new_n1297), .A4(KEYINPUT62), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n654), .A2(G213), .A3(G2897), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1297), .A2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1288), .A2(new_n1292), .A3(new_n1294), .A4(new_n1301), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1300), .B1(new_n1305), .B2(new_n1280), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1269), .B1(new_n1299), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT124), .B1(new_n1305), .B2(new_n1280), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1278), .B(new_n1277), .C1(new_n1252), .C2(new_n1142), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT124), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1310), .A2(new_n1311), .A3(new_n1303), .A4(new_n1304), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G375), .A2(G378), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1314), .A2(new_n1315), .A3(KEYINPUT63), .A4(new_n1295), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1264), .A2(new_n1300), .A3(new_n1266), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1271), .A2(new_n1279), .A3(new_n1297), .ZN(new_n1318));
  XOR2_X1   g1118(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1316), .B(new_n1317), .C1(new_n1318), .C2(new_n1320), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1313), .A2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1256), .B1(new_n1308), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1318), .A2(new_n1270), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1314), .A2(new_n1315), .A3(new_n1295), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1327));
  OAI22_X1  g1127(.A1(new_n1327), .A2(new_n1306), .B1(new_n1268), .B2(new_n1267), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1325), .A2(new_n1319), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1329), .A2(new_n1309), .A3(new_n1330), .A4(new_n1312), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1328), .A2(KEYINPUT127), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1323), .A2(new_n1332), .ZN(G405));
  NAND2_X1  g1133(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(new_n1297), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1253), .A2(new_n1314), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1335), .B(new_n1336), .ZN(G402));
endmodule


