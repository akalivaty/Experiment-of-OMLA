

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  AND2_X1 U324 ( .A1(n398), .A2(n397), .ZN(n399) );
  INV_X1 U325 ( .A(n529), .ZN(n397) );
  XNOR2_X1 U326 ( .A(n355), .B(G29GAT), .ZN(n356) );
  XNOR2_X1 U327 ( .A(KEYINPUT38), .B(n451), .ZN(n502) );
  NOR2_X1 U328 ( .A1(n566), .A2(n570), .ZN(n568) );
  XOR2_X1 U329 ( .A(n301), .B(n300), .Z(n292) );
  XOR2_X1 U330 ( .A(G99GAT), .B(G85GAT), .Z(n413) );
  INV_X1 U331 ( .A(KEYINPUT72), .ZN(n422) );
  XNOR2_X1 U332 ( .A(n531), .B(KEYINPUT93), .ZN(n398) );
  INV_X1 U333 ( .A(KEYINPUT54), .ZN(n470) );
  XNOR2_X1 U334 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U335 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U336 ( .A(n470), .B(KEYINPUT121), .ZN(n471) );
  XNOR2_X1 U337 ( .A(n425), .B(n424), .ZN(n429) );
  NOR2_X1 U338 ( .A1(n586), .A2(n411), .ZN(n412) );
  XNOR2_X1 U339 ( .A(n468), .B(n467), .ZN(n549) );
  XOR2_X1 U340 ( .A(n309), .B(n308), .Z(n477) );
  XOR2_X1 U341 ( .A(n454), .B(KEYINPUT41), .Z(n556) );
  XNOR2_X1 U342 ( .A(n365), .B(n364), .ZN(n519) );
  XNOR2_X1 U343 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n452) );
  XNOR2_X1 U345 ( .A(n481), .B(n480), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(G29GAT), .B(G43GAT), .Z(n294) );
  XNOR2_X1 U348 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n435) );
  XOR2_X1 U350 ( .A(n413), .B(G218GAT), .Z(n297) );
  XNOR2_X1 U351 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n295), .B(G162GAT), .ZN(n343) );
  XNOR2_X1 U353 ( .A(G134GAT), .B(n343), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U355 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n299) );
  NAND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U358 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n303) );
  XNOR2_X1 U359 ( .A(G106GAT), .B(G92GAT), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n304), .B(KEYINPUT75), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n292), .B(n305), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n435), .B(n306), .ZN(n309) );
  XNOR2_X1 U364 ( .A(G36GAT), .B(G190GAT), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n307), .B(KEYINPUT76), .ZN(n368) );
  INV_X1 U366 ( .A(n368), .ZN(n308) );
  XNOR2_X1 U367 ( .A(KEYINPUT36), .B(n477), .ZN(n586) );
  XOR2_X1 U368 ( .A(G211GAT), .B(G78GAT), .Z(n311) );
  XNOR2_X1 U369 ( .A(G183GAT), .B(G71GAT), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U371 ( .A(n312), .B(G155GAT), .Z(n314) );
  XOR2_X1 U372 ( .A(KEYINPUT69), .B(G1GAT), .Z(n447) );
  XNOR2_X1 U373 ( .A(n447), .B(G22GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n319) );
  XNOR2_X1 U375 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n315), .B(KEYINPUT13), .ZN(n414) );
  XOR2_X1 U377 ( .A(G15GAT), .B(G127GAT), .Z(n386) );
  XOR2_X1 U378 ( .A(n414), .B(n386), .Z(n317) );
  NAND2_X1 U379 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U380 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U381 ( .A(n319), .B(n318), .Z(n327) );
  XOR2_X1 U382 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n321) );
  XNOR2_X1 U383 ( .A(G8GAT), .B(G64GAT), .ZN(n320) );
  XNOR2_X1 U384 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U385 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n323) );
  XNOR2_X1 U386 ( .A(KEYINPUT77), .B(KEYINPUT12), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n559) );
  INV_X1 U390 ( .A(n559), .ZN(n582) );
  XOR2_X1 U391 ( .A(G141GAT), .B(G22GAT), .Z(n434) );
  XOR2_X1 U392 ( .A(KEYINPUT83), .B(KEYINPUT23), .Z(n329) );
  XNOR2_X1 U393 ( .A(KEYINPUT85), .B(KEYINPUT22), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U395 ( .A(n434), .B(n330), .Z(n332) );
  NAND2_X1 U396 ( .A1(G228GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U397 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U398 ( .A(G204GAT), .B(KEYINPUT24), .Z(n334) );
  XNOR2_X1 U399 ( .A(KEYINPUT86), .B(KEYINPUT84), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U401 ( .A(n336), .B(n335), .Z(n341) );
  XOR2_X1 U402 ( .A(G211GAT), .B(KEYINPUT21), .Z(n338) );
  XNOR2_X1 U403 ( .A(G197GAT), .B(G218GAT), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n338), .B(n337), .ZN(n376) );
  XNOR2_X1 U405 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n339) );
  XNOR2_X1 U406 ( .A(n339), .B(KEYINPUT2), .ZN(n361) );
  XNOR2_X1 U407 ( .A(n376), .B(n361), .ZN(n340) );
  XNOR2_X1 U408 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U409 ( .A(n343), .B(n342), .ZN(n345) );
  XNOR2_X1 U410 ( .A(G106GAT), .B(G78GAT), .ZN(n344) );
  XOR2_X1 U411 ( .A(n344), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U412 ( .A(n345), .B(n431), .ZN(n474) );
  XNOR2_X1 U413 ( .A(KEYINPUT28), .B(n474), .ZN(n494) );
  XOR2_X1 U414 ( .A(KEYINPUT87), .B(KEYINPUT4), .Z(n347) );
  XNOR2_X1 U415 ( .A(KEYINPUT5), .B(KEYINPUT88), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n347), .B(n346), .ZN(n365) );
  XOR2_X1 U417 ( .A(G148GAT), .B(G162GAT), .Z(n349) );
  XNOR2_X1 U418 ( .A(G141GAT), .B(G127GAT), .ZN(n348) );
  XNOR2_X1 U419 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U420 ( .A(KEYINPUT89), .B(G57GAT), .Z(n351) );
  XNOR2_X1 U421 ( .A(G1GAT), .B(G120GAT), .ZN(n350) );
  XNOR2_X1 U422 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U423 ( .A(n353), .B(n352), .Z(n359) );
  XNOR2_X1 U424 ( .A(G113GAT), .B(G134GAT), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n354), .B(KEYINPUT0), .ZN(n383) );
  XOR2_X1 U426 ( .A(G85GAT), .B(n383), .Z(n357) );
  NAND2_X1 U427 ( .A1(G225GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U428 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U429 ( .A(n360), .B(KEYINPUT6), .Z(n363) );
  XNOR2_X1 U430 ( .A(n361), .B(KEYINPUT1), .ZN(n362) );
  XNOR2_X1 U431 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U432 ( .A(G169GAT), .B(G8GAT), .Z(n436) );
  XOR2_X1 U433 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n370) );
  XOR2_X1 U434 ( .A(G64GAT), .B(G92GAT), .Z(n367) );
  XNOR2_X1 U435 ( .A(G176GAT), .B(G204GAT), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n430) );
  XNOR2_X1 U437 ( .A(n430), .B(n368), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U439 ( .A(n436), .B(n371), .Z(n373) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U442 ( .A(G183GAT), .B(KEYINPUT17), .Z(n375) );
  XNOR2_X1 U443 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n382) );
  XOR2_X1 U445 ( .A(n382), .B(n376), .Z(n377) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n522) );
  XNOR2_X1 U447 ( .A(KEYINPUT27), .B(n522), .ZN(n404) );
  NAND2_X1 U448 ( .A1(n519), .A2(n404), .ZN(n379) );
  XOR2_X1 U449 ( .A(KEYINPUT92), .B(n379), .Z(n547) );
  NAND2_X1 U450 ( .A1(n494), .A2(n547), .ZN(n531) );
  XOR2_X1 U451 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n381) );
  XNOR2_X1 U452 ( .A(G169GAT), .B(G99GAT), .ZN(n380) );
  XNOR2_X1 U453 ( .A(n381), .B(n380), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n383), .B(n382), .ZN(n394) );
  XOR2_X1 U455 ( .A(KEYINPUT80), .B(KEYINPUT20), .Z(n385) );
  XNOR2_X1 U456 ( .A(KEYINPUT65), .B(G176GAT), .ZN(n384) );
  XNOR2_X1 U457 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U458 ( .A(G120GAT), .B(G71GAT), .Z(n421) );
  XOR2_X1 U459 ( .A(G190GAT), .B(n421), .Z(n388) );
  XNOR2_X1 U460 ( .A(G43GAT), .B(n386), .ZN(n387) );
  XNOR2_X1 U461 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U462 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U463 ( .A1(G227GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U464 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U465 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n396), .B(n395), .ZN(n529) );
  XOR2_X1 U467 ( .A(KEYINPUT94), .B(n399), .Z(n410) );
  INV_X1 U468 ( .A(n519), .ZN(n408) );
  NAND2_X1 U469 ( .A1(n529), .A2(n522), .ZN(n400) );
  NAND2_X1 U470 ( .A1(n400), .A2(n474), .ZN(n401) );
  XNOR2_X1 U471 ( .A(n401), .B(KEYINPUT25), .ZN(n402) );
  XNOR2_X1 U472 ( .A(n402), .B(KEYINPUT95), .ZN(n406) );
  NOR2_X1 U473 ( .A1(n474), .A2(n529), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n403), .B(KEYINPUT26), .ZN(n572) );
  NAND2_X1 U475 ( .A1(n404), .A2(n572), .ZN(n405) );
  NAND2_X1 U476 ( .A1(n406), .A2(n405), .ZN(n407) );
  NAND2_X1 U477 ( .A1(n408), .A2(n407), .ZN(n409) );
  NAND2_X1 U478 ( .A1(n410), .A2(n409), .ZN(n483) );
  NAND2_X1 U479 ( .A1(n582), .A2(n483), .ZN(n411) );
  XNOR2_X1 U480 ( .A(KEYINPUT37), .B(n412), .ZN(n518) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n418) );
  INV_X1 U482 ( .A(n418), .ZN(n416) );
  AND2_X1 U483 ( .A1(G230GAT), .A2(G233GAT), .ZN(n417) );
  INV_X1 U484 ( .A(n417), .ZN(n415) );
  NAND2_X1 U485 ( .A1(n416), .A2(n415), .ZN(n420) );
  NAND2_X1 U486 ( .A1(n418), .A2(n417), .ZN(n419) );
  NAND2_X1 U487 ( .A1(n420), .A2(n419), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n421), .B(KEYINPUT73), .ZN(n423) );
  XOR2_X1 U489 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n427) );
  XNOR2_X1 U490 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n454) );
  XNOR2_X1 U495 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U497 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n439) );
  NAND2_X1 U498 ( .A1(G229GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U500 ( .A(n441), .B(n440), .Z(n446) );
  XOR2_X1 U501 ( .A(KEYINPUT67), .B(G113GAT), .Z(n443) );
  XNOR2_X1 U502 ( .A(G197GAT), .B(G15GAT), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n444), .B(KEYINPUT30), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n448) );
  XOR2_X1 U506 ( .A(n448), .B(n447), .Z(n450) );
  XNOR2_X1 U507 ( .A(G36GAT), .B(G50GAT), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n574) );
  INV_X1 U509 ( .A(n574), .ZN(n550) );
  NAND2_X1 U510 ( .A1(n454), .A2(n550), .ZN(n485) );
  NOR2_X1 U511 ( .A1(n518), .A2(n485), .ZN(n451) );
  NAND2_X1 U512 ( .A1(n502), .A2(n529), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n522), .B(KEYINPUT120), .ZN(n469) );
  INV_X1 U514 ( .A(n477), .ZN(n561) );
  XNOR2_X1 U515 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n574), .A2(n556), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U518 ( .A1(n559), .A2(n457), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT109), .ZN(n459) );
  NOR2_X1 U520 ( .A1(n561), .A2(n459), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT47), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n586), .A2(n582), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n461), .B(KEYINPUT45), .ZN(n462) );
  NAND2_X1 U524 ( .A1(n462), .A2(n454), .ZN(n463) );
  XOR2_X1 U525 ( .A(KEYINPUT110), .B(n463), .Z(n464) );
  NAND2_X1 U526 ( .A1(n464), .A2(n574), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n466), .A2(n465), .ZN(n468) );
  XNOR2_X1 U528 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n469), .A2(n549), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(n473) );
  NOR2_X1 U531 ( .A1(n519), .A2(n473), .ZN(n573) );
  NAND2_X1 U532 ( .A1(n573), .A2(n474), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n475), .B(KEYINPUT55), .ZN(n476) );
  NAND2_X1 U534 ( .A1(n476), .A2(n529), .ZN(n570) );
  NOR2_X1 U535 ( .A1(n477), .A2(n570), .ZN(n481) );
  XNOR2_X1 U536 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n479) );
  INV_X1 U537 ( .A(G190GAT), .ZN(n478) );
  XOR2_X1 U538 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n488) );
  NOR2_X1 U539 ( .A1(n561), .A2(n582), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n482), .B(KEYINPUT16), .ZN(n484) );
  NAND2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n505) );
  NOR2_X1 U542 ( .A1(n485), .A2(n505), .ZN(n486) );
  XNOR2_X1 U543 ( .A(KEYINPUT96), .B(n486), .ZN(n495) );
  NAND2_X1 U544 ( .A1(n495), .A2(n519), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n489), .ZN(G1324GAT) );
  NAND2_X1 U547 ( .A1(n495), .A2(n522), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n490), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U550 ( .A1(n495), .A2(n529), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(n493), .ZN(G1326GAT) );
  INV_X1 U553 ( .A(n494), .ZN(n526) );
  NAND2_X1 U554 ( .A1(n495), .A2(n526), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U556 ( .A1(n502), .A2(n519), .ZN(n499) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT99), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n497), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U560 ( .A1(n502), .A2(n522), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(KEYINPUT100), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT101), .Z(n504) );
  NAND2_X1 U564 ( .A1(n502), .A2(n526), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT102), .Z(n507) );
  XOR2_X1 U567 ( .A(n556), .B(KEYINPUT103), .Z(n566) );
  INV_X1 U568 ( .A(n566), .ZN(n534) );
  NAND2_X1 U569 ( .A1(n574), .A2(n534), .ZN(n517) );
  NOR2_X1 U570 ( .A1(n505), .A2(n517), .ZN(n514) );
  NAND2_X1 U571 ( .A1(n514), .A2(n519), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n509) );
  XOR2_X1 U573 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  XOR2_X1 U575 ( .A(G64GAT), .B(KEYINPUT105), .Z(n511) );
  NAND2_X1 U576 ( .A1(n514), .A2(n522), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n529), .A2(n514), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(KEYINPUT106), .ZN(n513) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U582 ( .A1(n514), .A2(n526), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  XOR2_X1 U584 ( .A(G85GAT), .B(KEYINPUT107), .Z(n521) );
  NOR2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n525) );
  NAND2_X1 U586 ( .A1(n525), .A2(n519), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n522), .A2(n525), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n529), .A2(n525), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT111), .Z(n533) );
  NAND2_X1 U596 ( .A1(n529), .A2(n549), .ZN(n530) );
  NOR2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n543), .A2(n550), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n536) );
  NAND2_X1 U601 ( .A1(n543), .A2(n534), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT112), .Z(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n540) );
  NAND2_X1 U607 ( .A1(n543), .A2(n559), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U611 ( .A1(n543), .A2(n561), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n546), .ZN(G1343GAT) );
  XOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT117), .Z(n552) );
  AND2_X1 U615 ( .A1(n572), .A2(n547), .ZN(n548) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n555) );
  INV_X1 U617 ( .A(n555), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n562), .A2(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(n558), .B(n557), .Z(G1345GAT) );
  NAND2_X1 U625 ( .A1(n562), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT119), .Z(n564) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n574), .A2(n570), .ZN(n565) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n565), .Z(G1348GAT) );
  XNOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n582), .A2(n570), .ZN(n571) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n571), .Z(G1350GAT) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n585) );
  NOR2_X1 U638 ( .A1(n574), .A2(n585), .ZN(n579) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n454), .A2(n585), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(G218GAT), .B(n589), .Z(G1355GAT) );
endmodule

