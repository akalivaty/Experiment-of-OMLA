//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT24), .B(G110), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT79), .B1(new_n193), .B2(new_n195), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n200));
  INV_X1    g014(.A(new_n190), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n200), .B(new_n192), .C1(new_n201), .C2(KEYINPUT23), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n198), .A2(new_n199), .B1(G110), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT16), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n209), .B(KEYINPUT80), .C1(KEYINPUT16), .C2(new_n206), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT80), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n208), .A3(new_n211), .A4(KEYINPUT16), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n204), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT16), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT80), .B1(new_n206), .B2(KEYINPUT16), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n204), .B(new_n212), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n203), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  OAI22_X1  g034(.A1(new_n202), .A2(G110), .B1(new_n194), .B2(new_n196), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n206), .A2(new_n208), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n204), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G137), .ZN(new_n226));
  INV_X1    g040(.A(G221), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n227), .A2(new_n187), .A3(G953), .ZN(new_n228));
  XOR2_X1   g042(.A(new_n226), .B(new_n228), .Z(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n218), .A2(KEYINPUT81), .A3(new_n224), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT81), .B1(new_n218), .B2(new_n224), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n230), .B1(new_n234), .B2(new_n229), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT25), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n188), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  INV_X1    g054(.A(new_n230), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n225), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n231), .ZN(new_n244));
  INV_X1    g058(.A(new_n229), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n241), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n240), .B1(new_n246), .B2(G902), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n235), .A2(KEYINPUT25), .A3(new_n236), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT82), .ZN(new_n249));
  AOI21_X1  g063(.A(G902), .B1(new_n187), .B2(G217), .ZN(new_n250));
  XOR2_X1   g064(.A(new_n250), .B(KEYINPUT83), .Z(new_n251));
  AOI22_X1  g065(.A1(new_n239), .A2(new_n249), .B1(new_n251), .B2(new_n235), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n254));
  INV_X1    g068(.A(G237), .ZN(new_n255));
  INV_X1    g069(.A(G953), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n255), .A2(new_n256), .A3(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n254), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT29), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT77), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n191), .A2(G116), .ZN(new_n264));
  INV_X1    g078(.A(G116), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G119), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT2), .B(G113), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G143), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT64), .B1(new_n270), .B2(G146), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(new_n204), .A3(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(G146), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT1), .B1(new_n270), .B2(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G128), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n204), .A2(G143), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n279), .A2(new_n280), .A3(new_n274), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  INV_X1    g098(.A(G137), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G134), .ZN(new_n286));
  INV_X1    g100(.A(G134), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G137), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT11), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n287), .B2(G137), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(KEYINPUT11), .A3(G134), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n291), .A2(new_n292), .A3(new_n288), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT66), .B(G131), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n269), .B1(new_n283), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n291), .A2(new_n292), .A3(new_n288), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G131), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n294), .A2(new_n291), .A3(new_n292), .A4(new_n288), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(KEYINPUT0), .A2(G128), .ZN(new_n301));
  NOR2_X1   g115(.A1(KEYINPUT0), .A2(G128), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(G143), .B(G146), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n275), .A2(new_n303), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n263), .B(KEYINPUT28), .C1(new_n296), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n283), .A2(new_n295), .ZN(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G119), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(new_n268), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT71), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n262), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n306), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n281), .B1(new_n275), .B2(new_n277), .ZN(new_n316));
  INV_X1    g130(.A(new_n289), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n299), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n310), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n312), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n263), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n311), .A2(KEYINPUT71), .A3(new_n312), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(KEYINPUT77), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT68), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n316), .B2(new_n318), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n283), .A2(new_n295), .A3(KEYINPUT68), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n306), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n300), .A2(KEYINPUT67), .A3(new_n305), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n332), .A3(new_n310), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n328), .A2(new_n332), .A3(KEYINPUT75), .A4(new_n310), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n300), .A2(KEYINPUT67), .A3(new_n305), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT67), .B1(new_n300), .B2(new_n305), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n326), .B(new_n327), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n339), .A2(new_n340), .A3(new_n269), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(new_n339), .B2(new_n269), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n335), .B(new_n336), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AOI211_X1 g157(.A(new_n261), .B(new_n324), .C1(new_n343), .C2(KEYINPUT28), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT78), .B1(new_n344), .B2(G902), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n346));
  INV_X1    g160(.A(new_n260), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(KEYINPUT30), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT30), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT65), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n300), .B1(new_n305), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n305), .A2(new_n350), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n349), .B(new_n308), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n310), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n333), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n347), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n308), .B1(new_n351), .B2(new_n352), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n269), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n312), .B1(new_n333), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n321), .A2(new_n322), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT70), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n260), .B(new_n361), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n346), .B(new_n356), .C1(new_n363), .C2(KEYINPUT73), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT74), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n356), .A2(new_n346), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n359), .A2(new_n360), .ZN(new_n368));
  INV_X1    g182(.A(new_n362), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT73), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n367), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n343), .A2(KEYINPUT28), .ZN(new_n376));
  INV_X1    g190(.A(new_n324), .ZN(new_n377));
  INV_X1    g191(.A(new_n261), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n236), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n345), .A2(new_n366), .A3(new_n375), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G472), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT72), .B1(new_n368), .B2(new_n369), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT72), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n385), .B(new_n362), .C1(new_n359), .C2(new_n360), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n348), .A2(new_n353), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n355), .B1(new_n387), .B2(new_n269), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT31), .B1(new_n388), .B2(new_n260), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT31), .ZN(new_n390));
  NOR4_X1   g204(.A1(new_n354), .A2(new_n390), .A3(new_n355), .A4(new_n347), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n384), .B(new_n386), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(G472), .A2(G902), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT32), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT32), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n253), .B1(new_n383), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G214), .B1(G237), .B2(G902), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT9), .B(G234), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n227), .B1(new_n402), .B2(new_n236), .ZN(new_n403));
  INV_X1    g217(.A(G104), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT3), .B1(new_n404), .B2(G107), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n406));
  INV_X1    g220(.A(G107), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(G104), .ZN(new_n408));
  INV_X1    g222(.A(G101), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(G107), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n405), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n407), .A3(G104), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT85), .B1(new_n404), .B2(G107), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n407), .A2(G104), .ZN(new_n415));
  OAI211_X1 g229(.A(G101), .B(new_n413), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n276), .A2(G128), .B1(new_n280), .B2(new_n274), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n411), .B(new_n416), .C1(new_n417), .C2(new_n281), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n411), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n420), .B2(new_n283), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n300), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(KEYINPUT12), .A3(new_n300), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT10), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT86), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n418), .A2(new_n430), .A3(new_n427), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n300), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n416), .A2(new_n411), .A3(KEYINPUT87), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT87), .B1(new_n416), .B2(new_n411), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT10), .B(new_n283), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n405), .A2(new_n408), .A3(new_n410), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G101), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT4), .A3(new_n411), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n440), .A3(G101), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n305), .A3(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n432), .A2(new_n433), .A3(new_n436), .A4(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G110), .B(G140), .ZN(new_n444));
  INV_X1    g258(.A(G227), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G953), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n444), .B(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n426), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n418), .A2(new_n430), .A3(new_n427), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n430), .B1(new_n418), .B2(new_n427), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n436), .A2(new_n442), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n300), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n448), .B1(new_n454), .B2(new_n443), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n449), .B1(new_n455), .B2(KEYINPUT88), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n426), .A2(new_n443), .A3(new_n457), .A4(new_n448), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G469), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n236), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n236), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n454), .A2(new_n443), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n448), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n426), .B2(new_n443), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT84), .B1(new_n426), .B2(new_n443), .ZN(new_n467));
  OAI22_X1  g281(.A1(new_n464), .A2(new_n466), .B1(new_n467), .B2(new_n448), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n462), .B1(new_n468), .B2(G469), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n403), .B1(new_n461), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G210), .B1(G237), .B2(G902), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n316), .A2(new_n207), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n207), .B2(new_n305), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n256), .A2(G224), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT92), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n473), .B(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n439), .A2(new_n269), .A3(new_n441), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G122), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n267), .A2(new_n268), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT5), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n191), .A3(G116), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT89), .ZN(new_n482));
  INV_X1    g296(.A(G113), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n309), .B2(KEYINPUT5), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n479), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n485), .B(new_n486), .C1(new_n435), .C2(new_n434), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n419), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n416), .A2(new_n411), .A3(KEYINPUT87), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n486), .B1(new_n492), .B2(new_n485), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n477), .B(new_n478), .C1(new_n488), .C2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n477), .B1(new_n488), .B2(new_n493), .ZN(new_n495));
  INV_X1    g309(.A(new_n478), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT91), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n494), .A2(KEYINPUT6), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n477), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n485), .B1(new_n435), .B2(new_n434), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT90), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n502), .B2(new_n487), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n503), .A2(new_n504), .A3(new_n497), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n476), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT93), .B(new_n476), .C1(new_n499), .C2(new_n505), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n474), .B1(new_n473), .B2(KEYINPUT94), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n511), .B(KEYINPUT7), .C1(KEYINPUT94), .C2(new_n474), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n485), .A2(new_n419), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n478), .B(KEYINPUT8), .Z(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n485), .A2(new_n419), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n474), .A2(KEYINPUT7), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n515), .A2(new_n516), .B1(new_n473), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n494), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n236), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n471), .B1(new_n510), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n471), .ZN(new_n524));
  AOI211_X1 g338(.A(new_n524), .B(new_n521), .C1(new_n508), .C2(new_n509), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n400), .B(new_n470), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n294), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT95), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT96), .B1(new_n528), .B2(G143), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n255), .A2(new_n256), .A3(G214), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(KEYINPUT96), .A2(G143), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n530), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n527), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n530), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT96), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(KEYINPUT95), .B2(new_n270), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n541), .B2(new_n533), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n294), .A3(new_n531), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n536), .A2(new_n543), .A3(new_n537), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n538), .A2(new_n216), .A3(new_n220), .A4(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(G113), .B(G122), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(new_n404), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n542), .A2(KEYINPUT97), .A3(new_n531), .ZN(new_n548));
  AND2_X1   g362(.A1(KEYINPUT18), .A2(G131), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n222), .B(new_n204), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n549), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n545), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n547), .B1(new_n545), .B2(new_n553), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n236), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G475), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT20), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n536), .A2(new_n543), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n222), .A2(KEYINPUT98), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT19), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n220), .B(new_n560), .C1(new_n562), .C2(G146), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n553), .ZN(new_n564));
  INV_X1    g378(.A(new_n547), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n554), .ZN(new_n567));
  NOR2_X1   g381(.A1(G475), .A2(G902), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n559), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  AOI211_X1 g384(.A(KEYINPUT20), .B(new_n570), .C1(new_n566), .C2(new_n554), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n558), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n558), .B(KEYINPUT99), .C1(new_n569), .C2(new_n571), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(G234), .A2(G237), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(G952), .A3(new_n256), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(G902), .A3(G953), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT21), .B(G898), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G116), .B(G122), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(new_n407), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n270), .A2(G128), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n189), .A2(G143), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n287), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT13), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n588), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n587), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT100), .B1(new_n593), .B2(KEYINPUT13), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n587), .A2(new_n595), .A3(new_n591), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n592), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n586), .B(new_n590), .C1(new_n597), .C2(new_n287), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n589), .B(new_n287), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n585), .A2(new_n407), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n265), .A2(KEYINPUT14), .A3(G122), .ZN(new_n601));
  INV_X1    g415(.A(new_n585), .ZN(new_n602));
  OAI211_X1 g416(.A(G107), .B(new_n601), .C1(new_n602), .C2(KEYINPUT14), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n402), .A2(G217), .A3(new_n256), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n598), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n598), .B2(new_n604), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n236), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G478), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(KEYINPUT15), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n598), .A2(new_n604), .ZN(new_n613));
  INV_X1    g427(.A(new_n605), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n615), .B2(new_n606), .ZN(new_n616));
  INV_X1    g430(.A(new_n611), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n576), .A2(new_n584), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n526), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n399), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  OAI211_X1 g438(.A(new_n400), .B(new_n584), .C1(new_n523), .C2(new_n525), .ZN(new_n625));
  INV_X1    g439(.A(new_n576), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n610), .A2(new_n236), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n616), .B2(new_n610), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT33), .B1(new_n607), .B2(new_n608), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n615), .A2(new_n630), .A3(new_n606), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n631), .A3(G478), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT102), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n625), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n384), .A2(new_n386), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n388), .A2(new_n260), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n390), .ZN(new_n640));
  INV_X1    g454(.A(new_n391), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(G472), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n394), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n252), .A2(new_n470), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n637), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n392), .A2(new_n236), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n648), .A2(G472), .B1(new_n393), .B2(new_n392), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n649), .A2(KEYINPUT101), .A3(new_n252), .A4(new_n470), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n636), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  OR2_X1    g467(.A1(new_n569), .A2(new_n571), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n619), .A3(new_n558), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n625), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n647), .A3(new_n650), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NAND2_X1  g473(.A1(new_n239), .A2(new_n249), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n245), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n234), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n251), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(new_n584), .A3(new_n620), .A4(new_n576), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n526), .A3(new_n645), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  AOI22_X1  g482(.A1(new_n382), .A2(G472), .B1(new_n395), .B2(new_n397), .ZN(new_n669));
  INV_X1    g483(.A(new_n470), .ZN(new_n670));
  INV_X1    g484(.A(new_n664), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n509), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n495), .A2(KEYINPUT6), .A3(new_n498), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n504), .B1(new_n503), .B2(new_n478), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n503), .A2(new_n497), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT93), .B1(new_n677), .B2(new_n476), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n522), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n524), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n510), .A2(new_n471), .A3(new_n522), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n400), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n578), .B(KEYINPUT103), .Z(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n685), .B1(new_n686), .B2(new_n581), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n683), .A2(new_n655), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n672), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XOR2_X1   g504(.A(new_n687), .B(KEYINPUT39), .Z(new_n691));
  NAND2_X1  g505(.A1(new_n470), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT40), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT38), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n682), .B(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n354), .A2(new_n355), .A3(new_n347), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n362), .B2(new_n343), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n398), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n574), .A2(new_n619), .A3(new_n575), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n702), .A2(new_n400), .A3(new_n671), .A4(new_n703), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n695), .A2(new_n696), .A3(new_n698), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n270), .ZN(G45));
  NAND2_X1  g520(.A1(new_n383), .A2(new_n398), .ZN(new_n707));
  INV_X1    g521(.A(new_n683), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n671), .A2(new_n670), .ZN(new_n709));
  INV_X1    g523(.A(new_n687), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n634), .A2(new_n574), .A3(new_n575), .A4(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n707), .A2(new_n708), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  AOI21_X1  g528(.A(new_n460), .B1(new_n459), .B2(new_n236), .ZN(new_n715));
  AOI211_X1 g529(.A(G469), .B(G902), .C1(new_n456), .C2(new_n458), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n715), .A2(new_n716), .A3(new_n403), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n399), .A2(new_n636), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND4_X1  g534(.A1(new_n656), .A2(new_n707), .A3(new_n252), .A4(new_n717), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NAND3_X1  g536(.A1(new_n682), .A2(new_n400), .A3(new_n717), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n665), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n707), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  OAI211_X1 g541(.A(new_n703), .B(new_n400), .C1(new_n523), .C2(new_n525), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n389), .A2(new_n391), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n369), .B1(new_n376), .B2(new_n377), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n393), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n252), .B(new_n731), .C1(new_n643), .C2(new_n644), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n717), .A2(new_n584), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n728), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(G122), .Z(G24));
  OAI21_X1  g549(.A(new_n731), .B1(new_n643), .B2(new_n644), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n736), .A2(new_n671), .A3(new_n711), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n724), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT105), .B(G125), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G27));
  AND4_X1   g554(.A1(new_n400), .A2(new_n680), .A3(new_n470), .A4(new_n681), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n707), .A2(new_n252), .A3(new_n712), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n399), .A2(KEYINPUT42), .A3(new_n712), .A4(new_n741), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NOR2_X1   g561(.A1(new_n655), .A2(new_n687), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n707), .A2(new_n252), .A3(new_n748), .A4(new_n741), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  INV_X1    g564(.A(new_n400), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n682), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n576), .A2(new_n634), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT43), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n576), .A2(new_n755), .A3(new_n634), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n645), .A3(new_n664), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n752), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n761), .B1(KEYINPUT108), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(G469), .B1(new_n468), .B2(KEYINPUT45), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n764), .A2(KEYINPUT106), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n764), .A2(KEYINPUT106), .B1(KEYINPUT45), .B2(new_n468), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n462), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n768));
  OR3_X1    g582(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT46), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n716), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n768), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n403), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n772), .A2(new_n773), .A3(new_n691), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n763), .B(new_n774), .C1(KEYINPUT108), .C2(new_n762), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n773), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n772), .A2(KEYINPUT47), .A3(new_n773), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n707), .A2(new_n252), .A3(new_n711), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n752), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NOR2_X1   g598(.A1(new_n619), .A2(new_n687), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n654), .A2(KEYINPUT109), .A3(new_n558), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n620), .A2(new_n710), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n572), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n400), .A2(new_n790), .A3(new_n680), .A4(new_n681), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n707), .A2(new_n709), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT110), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n707), .A2(new_n794), .A3(new_n791), .A4(new_n709), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n737), .A2(new_n741), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n749), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n746), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n625), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n576), .A2(new_n634), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n620), .B2(new_n576), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n647), .A2(new_n650), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n721), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n669), .A2(new_n723), .A3(new_n665), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n806), .A2(new_n666), .A3(new_n734), .ZN(new_n807));
  INV_X1    g621(.A(new_n717), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n669), .A2(new_n253), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n809), .A2(new_n636), .B1(new_n622), .B2(new_n399), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT111), .B1(new_n800), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n718), .A2(new_n721), .A3(new_n804), .A4(new_n623), .ZN(new_n813));
  INV_X1    g627(.A(new_n734), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n708), .A2(new_n725), .A3(new_n470), .A4(new_n649), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n726), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT111), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n798), .B1(new_n793), .B2(new_n795), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n746), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n664), .A2(new_n620), .A3(new_n576), .A4(new_n687), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n708), .A2(new_n702), .A3(new_n822), .A4(new_n470), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n689), .A2(new_n713), .A3(new_n738), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT52), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n672), .A2(new_n688), .B1(new_n724), .B2(new_n737), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n713), .A4(new_n823), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n821), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(KEYINPUT112), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n829), .B1(new_n812), .B2(new_n820), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(KEYINPUT53), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  INV_X1    g651(.A(new_n826), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n832), .B1(new_n838), .B2(KEYINPUT52), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n825), .A3(new_n828), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n840), .A2(new_n811), .A3(new_n800), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n833), .A2(new_n836), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n832), .B1(new_n826), .B2(new_n827), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n835), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n835), .A2(KEYINPUT53), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n715), .A2(new_n716), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n773), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n779), .A2(new_n780), .A3(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n757), .A2(new_n684), .A3(new_n732), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(new_n752), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n398), .A2(new_n252), .A3(new_n701), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n808), .A2(new_n682), .A3(new_n751), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n626), .A2(new_n634), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n857), .A2(new_n579), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n736), .A2(new_n671), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n758), .A2(new_n858), .A3(new_n685), .A4(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n861), .B1(new_n860), .B2(new_n863), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n808), .A2(new_n400), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n698), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n853), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n868), .B1(new_n698), .B2(new_n869), .ZN(new_n872));
  OAI211_X1 g686(.A(KEYINPUT115), .B(KEYINPUT50), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT115), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT50), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n855), .A2(new_n867), .A3(new_n873), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(G952), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n878), .B(G953), .C1(new_n853), .C2(new_n724), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n857), .A2(new_n579), .A3(new_n858), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n635), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n399), .A2(new_n758), .A3(new_n685), .A4(new_n858), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT113), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n855), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n876), .A2(new_n873), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n852), .A2(KEYINPUT113), .A3(new_n854), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n860), .A2(new_n863), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n892), .B2(new_n866), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n843), .A2(new_n847), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n878), .A2(new_n256), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n849), .A2(KEYINPUT49), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n849), .A2(KEYINPUT49), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n773), .A2(new_n400), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n753), .A4(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n698), .A3(new_n857), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT117), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n896), .A2(KEYINPUT117), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(G75));
  INV_X1    g720(.A(new_n833), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n836), .A2(new_n842), .ZN(new_n908));
  OAI211_X1 g722(.A(G210), .B(G902), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n677), .B(new_n476), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n909), .B2(new_n910), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n256), .A2(G952), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(G51));
  XNOR2_X1  g731(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n462), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n831), .A2(new_n832), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n841), .B1(new_n920), .B2(new_n834), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n837), .B1(new_n921), .B2(new_n833), .ZN(new_n922));
  INV_X1    g736(.A(new_n843), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n459), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n921), .A2(new_n833), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n765), .A2(new_n766), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT120), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(G902), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n916), .B1(new_n925), .B2(new_n929), .ZN(G54));
  AND2_X1   g744(.A1(KEYINPUT58), .A2(G475), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n926), .A2(G902), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n554), .A3(new_n566), .ZN(new_n933));
  INV_X1    g747(.A(new_n916), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n926), .A2(G902), .A3(new_n567), .A4(new_n931), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G60));
  XOR2_X1   g750(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n627), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n843), .B2(new_n847), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n629), .A2(new_n631), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT121), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n934), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n941), .A2(new_n938), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n922), .B2(new_n923), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT123), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n947), .B(new_n944), .C1(new_n922), .C2(new_n923), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n943), .B1(new_n946), .B2(new_n948), .ZN(G63));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT60), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n662), .B(new_n952), .C1(new_n907), .C2(new_n908), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n921), .B2(new_n833), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n953), .B(new_n934), .C1(new_n954), .C2(new_n235), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n907), .A2(new_n908), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n246), .B1(new_n958), .B2(new_n951), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n959), .A2(KEYINPUT61), .A3(new_n934), .A4(new_n953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n957), .A2(new_n960), .ZN(G66));
  INV_X1    g775(.A(G224), .ZN(new_n962));
  OAI21_X1  g776(.A(G953), .B1(new_n582), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n817), .B2(G953), .ZN(new_n964));
  INV_X1    g778(.A(new_n677), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(G898), .B2(new_n256), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT124), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n964), .B(new_n967), .ZN(G69));
  XOR2_X1   g782(.A(new_n562), .B(KEYINPUT125), .Z(new_n969));
  XOR2_X1   g783(.A(new_n387), .B(new_n969), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n826), .A2(new_n713), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n705), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT62), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n775), .A2(new_n783), .ZN(new_n975));
  INV_X1    g789(.A(new_n399), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n803), .A2(new_n752), .A3(new_n470), .A4(new_n691), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n974), .B(new_n975), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n971), .B1(new_n978), .B2(new_n256), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n774), .A2(new_n399), .A3(new_n708), .A4(new_n703), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n826), .A2(new_n713), .A3(new_n749), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n975), .A2(new_n746), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n256), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n256), .A2(G900), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT126), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n979), .B1(new_n971), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(G953), .B1(new_n445), .B2(new_n686), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n978), .B2(new_n811), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n992), .B(new_n260), .C1(new_n355), .C2(new_n354), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n991), .B1(new_n982), .B2(new_n811), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n354), .A2(new_n355), .A3(new_n260), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n916), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n845), .A2(new_n846), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n699), .A2(KEYINPUT127), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(new_n356), .Z(new_n1000));
  AND2_X1   g814(.A1(new_n1000), .A2(new_n991), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n997), .B1(new_n998), .B2(new_n1001), .ZN(G57));
endmodule


