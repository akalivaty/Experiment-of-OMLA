//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882;
  OR2_X1    g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR3_X1   g004(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT85), .B(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  OAI221_X1 g007(.A(new_n202), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n205), .B1(new_n202), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT84), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G155gat), .B2(G162gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT84), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n217), .A2(KEYINPUT80), .ZN(new_n218));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(KEYINPUT80), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G211gat), .B(G218gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n216), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G228gat), .ZN(new_n230));
  INV_X1    g029(.A(G233gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n209), .A2(new_n215), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n225), .B1(new_n233), .B2(KEYINPUT3), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT89), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n229), .B(new_n232), .C1(new_n224), .C2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n234), .A2(new_n223), .ZN(new_n237));
  OAI22_X1  g036(.A1(new_n228), .A2(new_n237), .B1(new_n230), .B2(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G22gat), .ZN(new_n240));
  INV_X1    g039(.A(G22gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n241), .A3(new_n238), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G78gat), .B(G106gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT31), .B(G50gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n239), .A2(new_n248), .A3(G22gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n246), .A2(new_n248), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n240), .A2(new_n242), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT27), .B(G183gat), .ZN(new_n253));
  INV_X1    g052(.A(G190gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(KEYINPUT28), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT27), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(G183gat), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n257), .A2(new_n259), .A3(new_n262), .A4(new_n254), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n263), .A2(KEYINPUT69), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT69), .B1(new_n263), .B2(new_n264), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n255), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n272), .B1(KEYINPUT26), .B2(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n275), .A2(KEYINPUT26), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n270), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(KEYINPUT70), .B(new_n255), .C1(new_n265), .C2(new_n266), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n269), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n270), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G183gat), .B2(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n284), .A2(new_n275), .B1(new_n270), .B2(new_n281), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n271), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT25), .B1(new_n275), .B2(new_n284), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT65), .B(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(KEYINPUT23), .A3(new_n273), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(new_n286), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n293), .B2(KEYINPUT25), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n280), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G127gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G134gat), .ZN(new_n297));
  INV_X1    g096(.A(G134gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G127gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  XOR2_X1   g101(.A(G113gat), .B(G120gat), .Z(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n301), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n302), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT71), .B(G134gat), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n307), .A2(G127gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n297), .B(KEYINPUT72), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n280), .A2(new_n313), .A3(new_n294), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G227gat), .A2(G233gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n316), .B(KEYINPUT64), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT32), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n315), .A2(new_n318), .B1(new_n319), .B2(KEYINPUT33), .ZN(new_n320));
  XNOR2_X1  g119(.A(G71gat), .B(G99gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G15gat), .B(G43gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  OAI21_X1  g124(.A(KEYINPUT76), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n280), .A2(new_n313), .A3(new_n294), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n313), .B1(new_n280), .B2(new_n294), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT33), .ZN(new_n330));
  OAI22_X1  g129(.A1(new_n329), .A2(new_n317), .B1(KEYINPUT32), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332));
  INV_X1    g131(.A(new_n325), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n318), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(KEYINPUT33), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n336), .A2(KEYINPUT32), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n312), .A2(new_n314), .A3(new_n316), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT34), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT34), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n312), .A2(new_n343), .A3(new_n314), .A4(new_n317), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT77), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347));
  INV_X1    g146(.A(new_n316), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n327), .A2(new_n328), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n347), .B(new_n344), .C1(new_n349), .C2(new_n343), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n340), .A2(new_n351), .A3(KEYINPUT78), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n338), .B1(new_n326), .B2(new_n334), .ZN(new_n353));
  INV_X1    g152(.A(new_n350), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n347), .B1(new_n342), .B2(new_n344), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT78), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n346), .A2(new_n357), .A3(new_n350), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n252), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G226gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(new_n231), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n362), .B1(new_n295), .B2(new_n225), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n295), .A2(new_n362), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n223), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(KEYINPUT81), .ZN(new_n367));
  INV_X1    g166(.A(new_n362), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n280), .B2(new_n294), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n363), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n366), .B1(new_n372), .B2(new_n223), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  INV_X1    g173(.A(G92gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT82), .B(G64gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  AOI21_X1  g177(.A(KEYINPUT30), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n370), .B1(new_n295), .B2(new_n362), .ZN(new_n380));
  AOI211_X1 g179(.A(KEYINPUT81), .B(new_n368), .C1(new_n280), .C2(new_n294), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n280), .B2(new_n294), .ZN(new_n382));
  OAI22_X1  g181(.A1(new_n380), .A2(new_n381), .B1(new_n362), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n224), .ZN(new_n384));
  INV_X1    g183(.A(new_n378), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n366), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n373), .A2(KEYINPUT30), .A3(new_n378), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n385), .B1(new_n384), .B2(new_n366), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(KEYINPUT83), .A3(KEYINPUT30), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n379), .B(new_n387), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT88), .B(KEYINPUT6), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT4), .B1(new_n311), .B2(new_n233), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n216), .A2(new_n397), .A3(new_n310), .A4(new_n305), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n216), .A2(new_n310), .A3(new_n305), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n216), .A2(new_n227), .B1(new_n310), .B2(new_n305), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n311), .A2(new_n233), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n400), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n311), .A2(KEYINPUT86), .A3(new_n233), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n402), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(new_n412), .A3(KEYINPUT5), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n396), .A2(new_n398), .B1(new_n404), .B2(new_n405), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT5), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n401), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G57gat), .B(G85gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT87), .B(KEYINPUT0), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n395), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n417), .A2(new_n423), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n360), .A2(new_n393), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n379), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT83), .B1(new_n391), .B2(KEYINPUT30), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n363), .A2(new_n224), .A3(new_n369), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n224), .B2(new_n383), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433));
  NOR4_X1   g232(.A1(new_n432), .A2(new_n389), .A3(new_n433), .A4(new_n385), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n429), .B(new_n386), .C1(new_n430), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n425), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n394), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT93), .B1(new_n417), .B2(new_n423), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n439));
  AOI211_X1 g238(.A(new_n439), .B(new_n422), .C1(new_n413), .C2(new_n416), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n437), .B1(new_n441), .B2(new_n424), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n435), .A2(KEYINPUT35), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n428), .A2(KEYINPUT35), .B1(new_n444), .B2(new_n360), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT36), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n446), .A2(KEYINPUT36), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n353), .A2(new_n356), .A3(new_n358), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n356), .B1(new_n358), .B2(new_n353), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n447), .B(new_n448), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n352), .A2(new_n359), .A3(new_n446), .A4(KEYINPUT36), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n414), .A2(new_n401), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n422), .B1(new_n454), .B2(KEYINPUT39), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n455), .A2(KEYINPUT91), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n402), .B1(new_n410), .B2(new_n411), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(KEYINPUT92), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(KEYINPUT92), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(KEYINPUT39), .A3(new_n454), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(KEYINPUT91), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n441), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n456), .A2(KEYINPUT40), .A3(new_n460), .A4(new_n461), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n252), .B1(new_n466), .B2(new_n435), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n468), .B(new_n385), .C1(new_n432), .C2(KEYINPUT37), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT94), .B1(new_n372), .B2(new_n224), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n364), .A2(new_n224), .A3(new_n365), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n383), .A2(new_n472), .A3(new_n223), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(KEYINPUT37), .B2(new_n474), .ZN(new_n475));
  OAI221_X1 g274(.A(new_n437), .B1(new_n432), .B2(new_n385), .C1(new_n441), .C2(new_n424), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT95), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n432), .A2(KEYINPUT37), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n385), .B1(new_n432), .B2(KEYINPUT37), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT38), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n474), .A2(KEYINPUT37), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n385), .A2(KEYINPUT37), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT38), .B1(new_n386), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n442), .A2(new_n391), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n477), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n453), .B1(new_n467), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n387), .B1(new_n390), .B2(new_n392), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(new_n427), .A3(new_n429), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n252), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n445), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT16), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(G1gat), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(G1gat), .B2(new_n495), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n498), .B(G8gat), .Z(new_n499));
  INV_X1    g298(.A(KEYINPUT21), .ZN(new_n500));
  XOR2_X1   g299(.A(G57gat), .B(G64gat), .Z(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT9), .ZN(new_n502));
  XOR2_X1   g301(.A(G71gat), .B(G78gat), .Z(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n503), .A2(KEYINPUT99), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(KEYINPUT99), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n499), .B1(new_n500), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(G183gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n500), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G231gat), .A2(G233gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G127gat), .B(G155gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G211gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n515), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G43gat), .B(G50gat), .Z(new_n521));
  OR2_X1    g320(.A1(new_n521), .A2(KEYINPUT96), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(KEYINPUT96), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT15), .A3(new_n523), .ZN(new_n524));
  OR3_X1    g323(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n521), .A2(new_n528), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT98), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT97), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n525), .A2(new_n534), .A3(new_n526), .ZN(new_n535));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  OAI211_X1 g335(.A(KEYINPUT97), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI22_X1  g337(.A1(new_n532), .A2(new_n533), .B1(new_n524), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT17), .ZN(new_n540));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  INV_X1    g341(.A(G99gat), .ZN(new_n543));
  INV_X1    g342(.A(G106gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT8), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n542), .B(new_n545), .C1(G85gat), .C2(G92gat), .ZN(new_n546));
  XOR2_X1   g345(.A(G99gat), .B(G106gat), .Z(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT101), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n540), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n550), .ZN(new_n553));
  AND2_X1   g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n539), .A2(new_n553), .B1(KEYINPUT41), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT102), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n554), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT100), .ZN(new_n563));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n561), .A2(new_n565), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n520), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n550), .B(new_n509), .Z(new_n570));
  NOR2_X1   g369(.A1(new_n550), .A2(new_n509), .ZN(new_n571));
  MUX2_X1   g370(.A(new_n570), .B(new_n571), .S(KEYINPUT10), .Z(new_n572));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n570), .A2(new_n573), .ZN(new_n575));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576));
  INV_X1    g375(.A(G204gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT103), .B(G176gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OR3_X1    g380(.A1(new_n574), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT104), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n574), .B2(new_n575), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n494), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n499), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n539), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n590), .B1(new_n540), .B2(new_n499), .ZN(new_n591));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT18), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n591), .A2(KEYINPUT18), .A3(new_n592), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n539), .B(new_n589), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n592), .B(KEYINPUT13), .Z(new_n596));
  AOI211_X1 g395(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598));
  INV_X1    g397(.A(G197gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT11), .B(G169gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n597), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n426), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G1gat), .ZN(G1324gat));
  INV_X1    g409(.A(KEYINPUT42), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT16), .B(G8gat), .ZN(new_n612));
  OR4_X1    g411(.A1(new_n611), .A2(new_n607), .A3(new_n393), .A4(new_n612), .ZN(new_n613));
  OR3_X1    g412(.A1(new_n607), .A2(KEYINPUT105), .A3(new_n393), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT105), .B1(new_n607), .B2(new_n393), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n611), .B1(new_n616), .B2(G8gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n612), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n613), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT106), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(G1325gat));
  NAND2_X1  g420(.A1(new_n352), .A2(new_n359), .ZN(new_n622));
  AOI21_X1  g421(.A(G15gat), .B1(new_n608), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n453), .A2(G15gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT107), .Z(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n608), .B2(new_n625), .ZN(G1326gat));
  INV_X1    g425(.A(new_n252), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n607), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT43), .B(G22gat), .Z(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT108), .B(KEYINPUT109), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n628), .B(new_n631), .ZN(G1327gat));
  INV_X1    g431(.A(KEYINPUT110), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n566), .A2(new_n567), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n489), .A2(new_n467), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n451), .A2(new_n452), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n493), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n444), .A2(new_n360), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n627), .B1(new_n449), .B2(new_n450), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT35), .B1(new_n639), .B2(new_n492), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n634), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n633), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n494), .C2(new_n634), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT35), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n435), .A2(new_n426), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n360), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n491), .A2(new_n647), .A3(new_n429), .A4(new_n442), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n639), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT111), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT111), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n640), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT44), .B1(new_n655), .B2(new_n637), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n568), .A2(KEYINPUT112), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n566), .A2(KEYINPUT112), .A3(new_n567), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n646), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n520), .ZN(new_n662));
  INV_X1    g461(.A(new_n606), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n662), .A2(new_n663), .A3(new_n585), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G29gat), .B1(new_n665), .B2(new_n427), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n642), .A2(new_n664), .ZN(new_n667));
  INV_X1    g466(.A(G29gat), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n426), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT45), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(new_n670), .ZN(G1328gat));
  OAI21_X1  g470(.A(G36gat), .B1(new_n665), .B2(new_n393), .ZN(new_n672));
  INV_X1    g471(.A(G36gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n667), .A2(new_n673), .A3(new_n435), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT46), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(G1329gat));
  INV_X1    g475(.A(KEYINPUT47), .ZN(new_n677));
  OAI21_X1  g476(.A(G43gat), .B1(new_n665), .B2(new_n636), .ZN(new_n678));
  INV_X1    g477(.A(G43gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n667), .A2(new_n679), .A3(new_n622), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n677), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n678), .A2(KEYINPUT113), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(KEYINPUT113), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT114), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n680), .B1(new_n684), .B2(KEYINPUT47), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n680), .A2(new_n684), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n681), .B1(new_n686), .B2(new_n687), .ZN(G1330gat));
  NAND3_X1  g487(.A1(new_n661), .A2(new_n252), .A3(new_n664), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n627), .A2(G50gat), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n689), .A2(G50gat), .B1(new_n667), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g491(.A1(new_n655), .A2(new_n637), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n693), .A2(new_n569), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n606), .A2(new_n586), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n427), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT115), .B(G57gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1332gat));
  NOR2_X1   g498(.A1(new_n696), .A2(new_n393), .ZN(new_n700));
  NOR2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  AND2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n700), .B2(new_n701), .ZN(G1333gat));
  OAI21_X1  g503(.A(G71gat), .B1(new_n696), .B2(new_n636), .ZN(new_n705));
  INV_X1    g504(.A(G71gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n622), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n696), .B2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g508(.A1(new_n696), .A2(new_n627), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(G78gat), .Z(G1335gat));
  INV_X1    g510(.A(KEYINPUT116), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n662), .A2(new_n606), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n585), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n661), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n644), .A2(new_n645), .B1(new_n659), .B2(new_n656), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT116), .B1(new_n718), .B2(new_n714), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G85gat), .B1(new_n721), .B2(new_n427), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n693), .A2(new_n568), .A3(new_n713), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT51), .Z(new_n724));
  NOR3_X1   g523(.A1(new_n586), .A2(G85gat), .A3(new_n427), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT117), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(new_n727), .ZN(G1336gat));
  AND4_X1   g527(.A1(new_n375), .A2(new_n724), .A3(new_n435), .A4(new_n585), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n718), .A2(new_n714), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n375), .B1(new_n730), .B2(new_n435), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n729), .A2(KEYINPUT52), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n435), .B1(new_n717), .B2(new_n720), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n729), .B1(new_n733), .B2(G92gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(G1337gat));
  AND2_X1   g535(.A1(new_n724), .A2(new_n585), .ZN(new_n737));
  AOI21_X1  g536(.A(G99gat), .B1(new_n737), .B2(new_n622), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n636), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G99gat), .ZN(G1338gat));
  INV_X1    g539(.A(new_n730), .ZN(new_n741));
  OAI21_X1  g540(.A(G106gat), .B1(new_n741), .B2(new_n627), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n544), .A3(new_n252), .A4(new_n585), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n627), .B1(new_n716), .B2(new_n719), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n746), .B2(new_n544), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n747), .A2(KEYINPUT118), .A3(KEYINPUT53), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT118), .B1(new_n747), .B2(KEYINPUT53), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(G1339gat));
  NOR2_X1   g549(.A1(new_n591), .A2(new_n592), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n595), .A2(new_n596), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n602), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT120), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n605), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n580), .B1(new_n574), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT54), .B1(new_n572), .B2(new_n573), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n574), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT119), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763));
  OR3_X1    g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n763), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n761), .B2(new_n763), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n764), .A2(new_n582), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n757), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n659), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n767), .B1(new_n604), .B2(new_n605), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n757), .A2(new_n586), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n657), .A2(new_n658), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n662), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n587), .A2(new_n606), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n639), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n426), .A3(new_n393), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n663), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g578(.A1(new_n777), .A2(new_n586), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g580(.A1(new_n777), .A2(new_n520), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT121), .B(G127gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1342gat));
  NOR2_X1   g583(.A1(new_n777), .A2(new_n634), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n307), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT56), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(new_n788), .A3(new_n307), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n787), .B(new_n789), .C1(new_n298), .C2(new_n785), .ZN(G1343gat));
  OAI21_X1  g589(.A(new_n634), .B1(new_n770), .B2(new_n771), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n662), .B1(new_n769), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n252), .B1(new_n792), .B2(new_n774), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT57), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(new_n252), .C1(new_n773), .C2(new_n774), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n453), .A2(new_n427), .A3(new_n435), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n794), .A2(new_n796), .A3(new_n606), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT122), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n798), .A2(new_n799), .A3(G141gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n798), .B2(G141gat), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n775), .A2(new_n627), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n802), .A2(new_n208), .A3(new_n606), .A4(new_n797), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n800), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT58), .B1(new_n798), .B2(G141gat), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n807), .A2(KEYINPUT123), .A3(new_n803), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT123), .B1(new_n807), .B2(new_n803), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n805), .A2(new_n806), .B1(new_n808), .B2(new_n809), .ZN(G1344gat));
  NAND2_X1  g609(.A1(new_n802), .A2(new_n797), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n207), .A3(new_n585), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT57), .B1(new_n775), .B2(new_n627), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n768), .A2(new_n568), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n662), .B1(new_n791), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n795), .B(new_n252), .C1(new_n817), .C2(new_n774), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n815), .A2(new_n585), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n797), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n814), .B1(new_n820), .B2(G148gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n794), .A2(new_n797), .A3(new_n796), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n814), .B1(new_n822), .B2(new_n586), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n207), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n813), .B1(new_n821), .B2(new_n824), .ZN(G1345gat));
  NOR3_X1   g624(.A1(new_n822), .A2(new_n203), .A3(new_n520), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n520), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT124), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n826), .B1(new_n828), .B2(new_n203), .ZN(G1346gat));
  INV_X1    g628(.A(new_n659), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n822), .A2(KEYINPUT125), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT125), .B1(new_n822), .B2(new_n830), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(G162gat), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n812), .A2(new_n204), .A3(new_n568), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1347gat));
  NAND3_X1  g634(.A1(new_n776), .A2(new_n427), .A3(new_n435), .ZN(new_n836));
  OAI21_X1  g635(.A(G169gat), .B1(new_n836), .B2(new_n663), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT126), .B1(new_n775), .B2(new_n426), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT126), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n839), .B(new_n427), .C1(new_n773), .C2(new_n774), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n393), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n360), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n606), .A2(new_n273), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n837), .B1(new_n842), .B2(new_n843), .ZN(G1348gat));
  NOR3_X1   g643(.A1(new_n836), .A2(new_n289), .A3(new_n586), .ZN(new_n845));
  INV_X1    g644(.A(new_n842), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n585), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n847), .B2(new_n274), .ZN(G1349gat));
  OAI21_X1  g647(.A(G183gat), .B1(new_n836), .B2(new_n520), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n662), .A2(new_n253), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT60), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(new_n849), .C1(new_n842), .C2(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n836), .B2(new_n634), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT61), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n846), .A2(new_n254), .A3(new_n659), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1351gat));
  AND3_X1   g658(.A1(new_n841), .A2(new_n252), .A3(new_n636), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n599), .A3(new_n606), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n453), .A2(new_n426), .A3(new_n393), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n815), .A2(new_n818), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G197gat), .B1(new_n863), .B2(new_n663), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(G1352gat));
  NAND4_X1  g664(.A1(new_n841), .A2(new_n252), .A3(new_n636), .A4(new_n585), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n866), .A2(KEYINPUT62), .A3(G204gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n819), .A2(new_n862), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(G204gat), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT62), .B1(new_n866), .B2(G204gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(G1353gat));
  NAND4_X1  g670(.A1(new_n815), .A2(new_n662), .A3(new_n818), .A4(new_n862), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G211gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n874));
  OR2_X1    g673(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n875));
  NAND2_X1  g674(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n872), .A2(G211gat), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n662), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n874), .B(new_n877), .C1(new_n878), .C2(G211gat), .ZN(G1354gat));
  INV_X1    g678(.A(G218gat), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n863), .A2(new_n880), .A3(new_n634), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n860), .A2(new_n659), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n880), .ZN(G1355gat));
endmodule


