

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U553 ( .A1(G2105), .A2(G2104), .ZN(n877) );
  XNOR2_X2 U554 ( .A(n527), .B(KEYINPUT64), .ZN(n613) );
  INV_X1 U555 ( .A(KEYINPUT26), .ZN(n688) );
  NOR2_X1 U556 ( .A1(n915), .A2(n692), .ZN(n698) );
  AND2_X1 U557 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U558 ( .A1(n759), .A2(n745), .ZN(n746) );
  NOR2_X1 U559 ( .A1(n751), .A2(n750), .ZN(n753) );
  NOR2_X1 U560 ( .A1(n759), .A2(n683), .ZN(n764) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n766) );
  INV_X1 U562 ( .A(G2105), .ZN(n526) );
  NOR2_X1 U563 ( .A1(n637), .A2(n543), .ZN(n646) );
  NOR2_X1 U564 ( .A1(G651), .A2(n637), .ZN(n644) );
  NOR2_X2 U565 ( .A1(n530), .A2(n529), .ZN(G160) );
  AND2_X1 U566 ( .A1(n526), .A2(G2104), .ZN(n873) );
  NAND2_X1 U567 ( .A1(n873), .A2(G101), .ZN(n519) );
  XNOR2_X1 U568 ( .A(n519), .B(KEYINPUT23), .ZN(n522) );
  NAND2_X1 U569 ( .A1(G113), .A2(n877), .ZN(n520) );
  XOR2_X1 U570 ( .A(KEYINPUT66), .B(n520), .Z(n521) );
  NOR2_X1 U571 ( .A1(n522), .A2(n521), .ZN(n525) );
  NOR2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X2 U573 ( .A(KEYINPUT17), .B(n523), .Z(n872) );
  NAND2_X1 U574 ( .A1(n872), .A2(G137), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n530) );
  NOR2_X1 U576 ( .A1(n526), .A2(G2104), .ZN(n527) );
  NAND2_X1 U577 ( .A1(G125), .A2(n613), .ZN(n528) );
  XNOR2_X1 U578 ( .A(KEYINPUT65), .B(n528), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G138), .A2(n872), .ZN(n532) );
  NAND2_X1 U580 ( .A1(G102), .A2(n873), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U582 ( .A1(G114), .A2(n877), .ZN(n534) );
  NAND2_X1 U583 ( .A1(G126), .A2(n613), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U585 ( .A1(n536), .A2(n535), .ZN(G164) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U587 ( .A1(n645), .A2(G89), .ZN(n537) );
  XNOR2_X1 U588 ( .A(KEYINPUT4), .B(n537), .ZN(n541) );
  XNOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .ZN(n538) );
  XNOR2_X1 U590 ( .A(n538), .B(KEYINPUT67), .ZN(n637) );
  INV_X1 U591 ( .A(G651), .ZN(n543) );
  NAND2_X1 U592 ( .A1(n646), .A2(G76), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT75), .B(n539), .Z(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U595 ( .A(KEYINPUT5), .B(n542), .ZN(n551) );
  NAND2_X1 U596 ( .A1(n644), .A2(G51), .ZN(n547) );
  NOR2_X1 U597 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U598 ( .A(KEYINPUT68), .B(n544), .Z(n545) );
  XNOR2_X1 U599 ( .A(KEYINPUT1), .B(n545), .ZN(n649) );
  NAND2_X1 U600 ( .A1(G63), .A2(n649), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n549) );
  XOR2_X1 U602 ( .A(KEYINPUT6), .B(KEYINPUT76), .Z(n548) );
  XNOR2_X1 U603 ( .A(n549), .B(n548), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U605 ( .A(KEYINPUT7), .B(n552), .ZN(G168) );
  XNOR2_X1 U606 ( .A(G168), .B(KEYINPUT8), .ZN(n553) );
  XNOR2_X1 U607 ( .A(n553), .B(KEYINPUT77), .ZN(G286) );
  NAND2_X1 U608 ( .A1(G85), .A2(n645), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G72), .A2(n646), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U611 ( .A1(n644), .A2(G47), .ZN(n557) );
  NAND2_X1 U612 ( .A1(G60), .A2(n649), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n558) );
  OR2_X1 U614 ( .A1(n559), .A2(n558), .ZN(G290) );
  NAND2_X1 U615 ( .A1(n644), .A2(G52), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G64), .A2(n649), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n566) );
  NAND2_X1 U618 ( .A1(G90), .A2(n645), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G77), .A2(n646), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n564), .Z(n565) );
  NOR2_X1 U622 ( .A1(n566), .A2(n565), .ZN(G171) );
  AND2_X1 U623 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n819) );
  NAND2_X1 U628 ( .A1(n819), .A2(G567), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  NAND2_X1 U630 ( .A1(n645), .A2(G81), .ZN(n569) );
  XNOR2_X1 U631 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G68), .A2(n646), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U634 ( .A(KEYINPUT13), .B(n572), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n649), .A2(G56), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n573), .Z(n576) );
  NAND2_X1 U637 ( .A1(G43), .A2(n644), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT71), .B(n574), .ZN(n575) );
  NOR2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n915) );
  INV_X1 U641 ( .A(n915), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n579), .A2(G860), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT72), .B(n580), .ZN(G153) );
  INV_X1 U644 ( .A(G171), .ZN(G301) );
  NAND2_X1 U645 ( .A1(G54), .A2(n644), .ZN(n587) );
  NAND2_X1 U646 ( .A1(G92), .A2(n645), .ZN(n582) );
  NAND2_X1 U647 ( .A1(G66), .A2(n649), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G79), .A2(n646), .ZN(n583) );
  XNOR2_X1 U650 ( .A(KEYINPUT73), .B(n583), .ZN(n584) );
  NOR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X2 U653 ( .A(n588), .B(KEYINPUT15), .ZN(n920) );
  INV_X1 U654 ( .A(n920), .ZN(n605) );
  NOR2_X1 U655 ( .A1(G868), .A2(n605), .ZN(n590) );
  INV_X1 U656 ( .A(G868), .ZN(n663) );
  NOR2_X1 U657 ( .A1(n663), .A2(G301), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U659 ( .A(KEYINPUT74), .B(n591), .ZN(G284) );
  NAND2_X1 U660 ( .A1(n649), .A2(G65), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n592), .B(KEYINPUT70), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G91), .A2(n645), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G53), .A2(n644), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G78), .A2(n646), .ZN(n595) );
  XNOR2_X1 U666 ( .A(KEYINPUT69), .B(n595), .ZN(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n599), .A2(n598), .ZN(G299) );
  NOR2_X1 U669 ( .A1(G286), .A2(n663), .ZN(n601) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(G297) );
  INV_X1 U672 ( .A(G559), .ZN(n602) );
  NOR2_X1 U673 ( .A1(G860), .A2(n602), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n603), .B(KEYINPUT78), .ZN(n604) );
  NOR2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(KEYINPUT16), .ZN(n607) );
  XNOR2_X1 U677 ( .A(n607), .B(KEYINPUT79), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n915), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G868), .A2(n920), .ZN(n608) );
  NOR2_X1 U680 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G99), .A2(n873), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G111), .A2(n877), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n618) );
  NAND2_X1 U685 ( .A1(n613), .A2(G123), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n872), .A2(G135), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n970) );
  XNOR2_X1 U690 ( .A(G2096), .B(n970), .ZN(n620) );
  INV_X1 U691 ( .A(G2100), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(G156) );
  NAND2_X1 U693 ( .A1(G73), .A2(n646), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT2), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(KEYINPUT84), .ZN(n624) );
  NAND2_X1 U696 ( .A1(G86), .A2(n645), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G48), .A2(n644), .ZN(n625) );
  XNOR2_X1 U699 ( .A(KEYINPUT85), .B(n625), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n649), .A2(G61), .ZN(n628) );
  XOR2_X1 U702 ( .A(KEYINPUT83), .B(n628), .Z(n629) );
  NAND2_X1 U703 ( .A1(n630), .A2(n629), .ZN(G305) );
  NAND2_X1 U704 ( .A1(G88), .A2(n645), .ZN(n632) );
  NAND2_X1 U705 ( .A1(G75), .A2(n646), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n644), .A2(G50), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G62), .A2(n649), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U710 ( .A1(n636), .A2(n635), .ZN(G166) );
  NAND2_X1 U711 ( .A1(G87), .A2(n637), .ZN(n639) );
  NAND2_X1 U712 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U714 ( .A1(n649), .A2(n640), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n644), .A2(G49), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U717 ( .A1(G559), .A2(n920), .ZN(n643) );
  XOR2_X1 U718 ( .A(n915), .B(n643), .Z(n823) );
  NAND2_X1 U719 ( .A1(G55), .A2(n644), .ZN(n654) );
  NAND2_X1 U720 ( .A1(G93), .A2(n645), .ZN(n648) );
  NAND2_X1 U721 ( .A1(G80), .A2(n646), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U723 ( .A1(G67), .A2(n649), .ZN(n650) );
  XNOR2_X1 U724 ( .A(KEYINPUT81), .B(n650), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n655), .B(KEYINPUT82), .ZN(n826) );
  XOR2_X1 U728 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n656) );
  XNOR2_X1 U729 ( .A(G288), .B(n656), .ZN(n657) );
  XNOR2_X1 U730 ( .A(G166), .B(n657), .ZN(n659) );
  INV_X1 U731 ( .A(G299), .ZN(n923) );
  XNOR2_X1 U732 ( .A(G290), .B(n923), .ZN(n658) );
  XNOR2_X1 U733 ( .A(n659), .B(n658), .ZN(n660) );
  XOR2_X1 U734 ( .A(n826), .B(n660), .Z(n661) );
  XNOR2_X1 U735 ( .A(G305), .B(n661), .ZN(n893) );
  XNOR2_X1 U736 ( .A(n823), .B(n893), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n662), .A2(G868), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n663), .A2(n826), .ZN(n664) );
  NAND2_X1 U739 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2084), .A2(G2078), .ZN(n666) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U742 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U746 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n671) );
  NAND2_X1 U747 ( .A1(G132), .A2(G82), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U749 ( .A1(n672), .A2(G218), .ZN(n673) );
  NAND2_X1 U750 ( .A1(G96), .A2(n673), .ZN(n828) );
  NAND2_X1 U751 ( .A1(n828), .A2(G2106), .ZN(n678) );
  NAND2_X1 U752 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U753 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U754 ( .A1(G108), .A2(n675), .ZN(n827) );
  NAND2_X1 U755 ( .A1(G567), .A2(n827), .ZN(n676) );
  XNOR2_X1 U756 ( .A(KEYINPUT88), .B(n676), .ZN(n677) );
  NAND2_X1 U757 ( .A1(n678), .A2(n677), .ZN(n829) );
  NAND2_X1 U758 ( .A1(G661), .A2(G483), .ZN(n679) );
  XOR2_X1 U759 ( .A(KEYINPUT89), .B(n679), .Z(n680) );
  NOR2_X1 U760 ( .A1(n829), .A2(n680), .ZN(n822) );
  NAND2_X1 U761 ( .A1(n822), .A2(G36), .ZN(G176) );
  INV_X1 U762 ( .A(G166), .ZN(G303) );
  NAND2_X1 U763 ( .A1(G160), .A2(G40), .ZN(n765) );
  INV_X1 U764 ( .A(n765), .ZN(n681) );
  NAND2_X2 U765 ( .A1(n681), .A2(n766), .ZN(n725) );
  NAND2_X1 U766 ( .A1(G8), .A2(n725), .ZN(n759) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n682) );
  XOR2_X1 U768 ( .A(n682), .B(KEYINPUT24), .Z(n683) );
  XOR2_X1 U769 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NOR2_X1 U770 ( .A1(n948), .A2(n725), .ZN(n684) );
  XNOR2_X1 U771 ( .A(n684), .B(KEYINPUT97), .ZN(n686) );
  INV_X1 U772 ( .A(G1961), .ZN(n989) );
  NAND2_X1 U773 ( .A1(n989), .A2(n725), .ZN(n685) );
  NAND2_X1 U774 ( .A1(n686), .A2(n685), .ZN(n718) );
  NAND2_X1 U775 ( .A1(n718), .A2(G171), .ZN(n714) );
  INV_X1 U776 ( .A(G1996), .ZN(n687) );
  NOR2_X2 U777 ( .A1(n725), .A2(n687), .ZN(n689) );
  XNOR2_X1 U778 ( .A(n689), .B(n688), .ZN(n691) );
  NAND2_X1 U779 ( .A1(n725), .A2(G1341), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U781 ( .A1(n920), .A2(n698), .ZN(n697) );
  NAND2_X1 U782 ( .A1(n725), .A2(G1348), .ZN(n693) );
  XNOR2_X1 U783 ( .A(n693), .B(KEYINPUT98), .ZN(n695) );
  INV_X1 U784 ( .A(n725), .ZN(n701) );
  NAND2_X1 U785 ( .A1(n701), .A2(G2067), .ZN(n694) );
  NAND2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n700) );
  OR2_X1 U788 ( .A1(n920), .A2(n698), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n700), .A2(n699), .ZN(n706) );
  NAND2_X1 U790 ( .A1(n701), .A2(G2072), .ZN(n702) );
  XNOR2_X1 U791 ( .A(n702), .B(KEYINPUT27), .ZN(n704) );
  AND2_X1 U792 ( .A1(G1956), .A2(n725), .ZN(n703) );
  NOR2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U794 ( .A1(n923), .A2(n707), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U796 ( .A1(n923), .A2(n707), .ZN(n708) );
  XOR2_X1 U797 ( .A(n708), .B(KEYINPUT28), .Z(n709) );
  NAND2_X1 U798 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U799 ( .A(n711), .B(KEYINPUT29), .ZN(n712) );
  INV_X1 U800 ( .A(n712), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n723) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n759), .ZN(n736) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n725), .ZN(n733) );
  NOR2_X1 U804 ( .A1(n736), .A2(n733), .ZN(n715) );
  NAND2_X1 U805 ( .A1(G8), .A2(n715), .ZN(n716) );
  XNOR2_X1 U806 ( .A(KEYINPUT30), .B(n716), .ZN(n717) );
  NOR2_X1 U807 ( .A1(G168), .A2(n717), .ZN(n720) );
  NOR2_X1 U808 ( .A1(G171), .A2(n718), .ZN(n719) );
  NOR2_X1 U809 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U810 ( .A(KEYINPUT31), .B(n721), .Z(n722) );
  NAND2_X1 U811 ( .A1(n723), .A2(n722), .ZN(n734) );
  NAND2_X1 U812 ( .A1(n734), .A2(G286), .ZN(n724) );
  XNOR2_X1 U813 ( .A(n724), .B(KEYINPUT100), .ZN(n730) );
  NOR2_X1 U814 ( .A1(G1971), .A2(n759), .ZN(n727) );
  NOR2_X1 U815 ( .A1(G2090), .A2(n725), .ZN(n726) );
  NOR2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U817 ( .A1(n728), .A2(G303), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U820 ( .A(n732), .B(KEYINPUT32), .ZN(n754) );
  NAND2_X1 U821 ( .A1(G8), .A2(n733), .ZN(n738) );
  XNOR2_X1 U822 ( .A(KEYINPUT99), .B(n734), .ZN(n735) );
  NOR2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n755) );
  NAND2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n924) );
  AND2_X1 U826 ( .A1(n755), .A2(n924), .ZN(n739) );
  NAND2_X1 U827 ( .A1(n754), .A2(n739), .ZN(n744) );
  INV_X1 U828 ( .A(n924), .ZN(n742) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n748) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n748), .A2(n740), .ZN(n919) );
  XOR2_X1 U832 ( .A(n919), .B(KEYINPUT101), .Z(n741) );
  OR2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U834 ( .A1(n746), .A2(KEYINPUT33), .ZN(n747) );
  XNOR2_X1 U835 ( .A(n747), .B(KEYINPUT102), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n748), .A2(KEYINPUT33), .ZN(n749) );
  NOR2_X1 U837 ( .A1(n759), .A2(n749), .ZN(n750) );
  XNOR2_X1 U838 ( .A(G1981), .B(KEYINPUT103), .ZN(n752) );
  XNOR2_X1 U839 ( .A(n752), .B(G305), .ZN(n932) );
  NAND2_X1 U840 ( .A1(n753), .A2(n932), .ZN(n762) );
  NAND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n758) );
  NOR2_X1 U842 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U843 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n760) );
  NAND2_X1 U845 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U847 ( .A1(n764), .A2(n763), .ZN(n784) );
  NOR2_X1 U848 ( .A1(n766), .A2(n765), .ZN(n814) );
  XNOR2_X1 U849 ( .A(n814), .B(KEYINPUT96), .ZN(n783) );
  XOR2_X1 U850 ( .A(KEYINPUT95), .B(G1991), .Z(n942) );
  NAND2_X1 U851 ( .A1(G95), .A2(n873), .ZN(n768) );
  NAND2_X1 U852 ( .A1(G107), .A2(n877), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U854 ( .A1(G131), .A2(n872), .ZN(n769) );
  XOR2_X1 U855 ( .A(KEYINPUT94), .B(n769), .Z(n770) );
  NOR2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G119), .A2(n613), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n859) );
  NAND2_X1 U859 ( .A1(n942), .A2(n859), .ZN(n782) );
  NAND2_X1 U860 ( .A1(G117), .A2(n877), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G129), .A2(n613), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U863 ( .A1(n873), .A2(G105), .ZN(n776) );
  XOR2_X1 U864 ( .A(KEYINPUT38), .B(n776), .Z(n777) );
  NOR2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n872), .A2(G141), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n889) );
  NAND2_X1 U868 ( .A1(G1996), .A2(n889), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n977) );
  AND2_X1 U870 ( .A1(n783), .A2(n977), .ZN(n804) );
  NOR2_X1 U871 ( .A1(n784), .A2(n804), .ZN(n800) );
  XNOR2_X1 U872 ( .A(G1986), .B(G290), .ZN(n917) );
  NAND2_X1 U873 ( .A1(n917), .A2(n814), .ZN(n785) );
  XNOR2_X1 U874 ( .A(n785), .B(KEYINPUT90), .ZN(n798) );
  XOR2_X1 U875 ( .A(G2067), .B(KEYINPUT37), .Z(n801) );
  NAND2_X1 U876 ( .A1(G116), .A2(n877), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G128), .A2(n613), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U879 ( .A(KEYINPUT35), .B(n788), .ZN(n795) );
  XNOR2_X1 U880 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n872), .A2(G140), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n873), .A2(G104), .ZN(n789) );
  XOR2_X1 U883 ( .A(KEYINPUT91), .B(n789), .Z(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U885 ( .A(n793), .B(n792), .Z(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U887 ( .A(KEYINPUT36), .B(n796), .ZN(n883) );
  NAND2_X1 U888 ( .A1(n801), .A2(n883), .ZN(n797) );
  XNOR2_X1 U889 ( .A(n797), .B(KEYINPUT93), .ZN(n973) );
  NAND2_X1 U890 ( .A1(n814), .A2(n973), .ZN(n809) );
  AND2_X1 U891 ( .A1(n798), .A2(n809), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n817) );
  NOR2_X1 U893 ( .A1(n883), .A2(n801), .ZN(n982) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n889), .ZN(n966) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n942), .A2(n859), .ZN(n971) );
  NOR2_X1 U897 ( .A1(n802), .A2(n971), .ZN(n803) );
  NOR2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U899 ( .A(n805), .B(KEYINPUT104), .ZN(n806) );
  NOR2_X1 U900 ( .A1(n966), .A2(n806), .ZN(n808) );
  XOR2_X1 U901 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n807) );
  XNOR2_X1 U902 ( .A(n808), .B(n807), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U904 ( .A(KEYINPUT106), .B(n811), .Z(n812) );
  NOR2_X1 U905 ( .A1(n982), .A2(n812), .ZN(n813) );
  XNOR2_X1 U906 ( .A(KEYINPUT107), .B(n813), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U909 ( .A(n818), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U912 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n822), .A2(n821), .ZN(G188) );
  XOR2_X1 U916 ( .A(n823), .B(KEYINPUT80), .Z(n824) );
  NOR2_X1 U917 ( .A1(G860), .A2(n824), .ZN(n825) );
  XOR2_X1 U918 ( .A(n826), .B(n825), .Z(G145) );
  INV_X1 U919 ( .A(G132), .ZN(G219) );
  INV_X1 U920 ( .A(G120), .ZN(G236) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  INV_X1 U922 ( .A(G82), .ZN(G220) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  INV_X1 U926 ( .A(n829), .ZN(G319) );
  XOR2_X1 U927 ( .A(KEYINPUT112), .B(G1961), .Z(n831) );
  XNOR2_X1 U928 ( .A(G1991), .B(G1996), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U930 ( .A(n832), .B(KEYINPUT41), .Z(n834) );
  XNOR2_X1 U931 ( .A(G1966), .B(G1981), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U933 ( .A(G1976), .B(G1971), .Z(n836) );
  XNOR2_X1 U934 ( .A(G1986), .B(G1956), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U936 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U937 ( .A(G2474), .B(KEYINPUT111), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT110), .Z(n842) );
  XNOR2_X1 U940 ( .A(G2067), .B(KEYINPUT43), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U942 ( .A(n843), .B(KEYINPUT42), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2072), .B(G2090), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U945 ( .A(G2678), .B(G2100), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2084), .B(G2078), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(G227) );
  NAND2_X1 U949 ( .A1(G112), .A2(n877), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n850), .B(KEYINPUT114), .ZN(n853) );
  NAND2_X1 U951 ( .A1(G136), .A2(n872), .ZN(n851) );
  XOR2_X1 U952 ( .A(KEYINPUT113), .B(n851), .Z(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U954 ( .A1(n613), .A2(G124), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n873), .A2(G100), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U958 ( .A1(n858), .A2(n857), .ZN(G162) );
  XNOR2_X1 U959 ( .A(G160), .B(n970), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n859), .B(G164), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n871) );
  NAND2_X1 U962 ( .A1(G118), .A2(n877), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G130), .A2(n613), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U965 ( .A1(n873), .A2(G106), .ZN(n864) );
  XOR2_X1 U966 ( .A(KEYINPUT115), .B(n864), .Z(n866) );
  NAND2_X1 U967 ( .A1(n872), .A2(G142), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U969 ( .A(KEYINPUT45), .B(n867), .Z(n868) );
  NOR2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U971 ( .A(n871), .B(n870), .Z(n885) );
  NAND2_X1 U972 ( .A1(G139), .A2(n872), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G103), .A2(n873), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U975 ( .A(KEYINPUT116), .B(n876), .ZN(n882) );
  NAND2_X1 U976 ( .A1(G115), .A2(n877), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G127), .A2(n613), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n961) );
  XNOR2_X1 U981 ( .A(n883), .B(n961), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n891) );
  XOR2_X1 U983 ( .A(KEYINPUT117), .B(KEYINPUT46), .Z(n887) );
  XNOR2_X1 U984 ( .A(G162), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U988 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U989 ( .A(n915), .B(n893), .ZN(n895) );
  XNOR2_X1 U990 ( .A(G171), .B(n920), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n896), .B(G286), .ZN(n897) );
  NOR2_X1 U993 ( .A1(G37), .A2(n897), .ZN(G397) );
  XNOR2_X1 U994 ( .A(G2435), .B(G2443), .ZN(n907) );
  XOR2_X1 U995 ( .A(G2454), .B(G2430), .Z(n899) );
  XNOR2_X1 U996 ( .A(G2446), .B(KEYINPUT109), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U998 ( .A(G2451), .B(G2427), .Z(n901) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1001 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT108), .B(G2438), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n908), .A2(G14), .ZN(n914) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n914), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n914), .ZN(G401) );
  XNOR2_X1 U1015 ( .A(G16), .B(KEYINPUT56), .ZN(n938) );
  XNOR2_X1 U1016 ( .A(G1341), .B(n915), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n931) );
  XNOR2_X1 U1019 ( .A(n920), .B(G1348), .ZN(n929) );
  XNOR2_X1 U1020 ( .A(G171), .B(G1961), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(G1971), .A2(G303), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n923), .B(G1956), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(G1966), .B(G168), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(n934), .B(KEYINPUT57), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n1020) );
  XNOR2_X1 U1033 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n985) );
  XNOR2_X1 U1034 ( .A(G1996), .B(G32), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G33), .B(G2072), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n947) );
  XOR2_X1 U1037 ( .A(G2067), .B(G26), .Z(n941) );
  NAND2_X1 U1038 ( .A1(n941), .A2(G28), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(KEYINPUT122), .B(n942), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(G25), .B(n943), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G27), .B(n948), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT53), .B(n951), .Z(n954) );
  XOR2_X1 U1046 ( .A(KEYINPUT54), .B(G34), .Z(n952) );
  XNOR2_X1 U1047 ( .A(G2084), .B(n952), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G35), .B(G2090), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n985), .B(n957), .ZN(n959) );
  INV_X1 U1052 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n960), .A2(G11), .ZN(n1018) );
  XOR2_X1 U1055 ( .A(G2072), .B(n961), .Z(n963) );
  XOR2_X1 U1056 ( .A(G164), .B(G2078), .Z(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1058 ( .A(KEYINPUT50), .B(n964), .Z(n969) );
  XOR2_X1 U1059 ( .A(G2090), .B(G162), .Z(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT51), .B(n967), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n980) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n975) );
  XOR2_X1 U1064 ( .A(G160), .B(G2084), .Z(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(n978), .B(KEYINPUT118), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1070 ( .A1(n982), .A2(n981), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(n984), .B(n983), .ZN(n986) );
  NOR2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  NAND2_X1 U1075 ( .A1(n988), .A2(G29), .ZN(n1016) );
  XNOR2_X1 U1076 ( .A(G5), .B(n989), .ZN(n1009) );
  XOR2_X1 U1077 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n996) );
  XNOR2_X1 U1078 ( .A(G1986), .B(G24), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n994) );
  XOR2_X1 U1081 ( .A(G1976), .B(KEYINPUT124), .Z(n992) );
  XNOR2_X1 U1082 ( .A(G23), .B(n992), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n996), .B(n995), .ZN(n1007) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G20), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G1341), .B(G19), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G6), .B(G1981), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(KEYINPUT123), .B(n999), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(G4), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(G21), .B(G1966), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(KEYINPUT61), .B(n1012), .Z(n1013) );
  NOR2_X1 U1100 ( .A1(G16), .A2(n1013), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1014), .Z(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(n1021), .B(KEYINPUT127), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1022), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

