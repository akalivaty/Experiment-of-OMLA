//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n468), .B2(new_n470), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n467), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT67), .Z(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n463), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  INV_X1    g057(.A(new_n465), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n463), .A2(KEYINPUT68), .A3(G126), .A4(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n464), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n463), .A2(new_n498), .A3(G138), .A4(new_n464), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n472), .B2(new_n473), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n495), .B1(new_n500), .B2(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(G62), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n511), .B1(new_n515), .B2(G651), .ZN(G166));
  NAND3_X1  g091(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n517));
  XOR2_X1   g092(.A(new_n517), .B(KEYINPUT71), .Z(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  OAI221_X1 g097(.A(new_n520), .B1(new_n509), .B2(new_n521), .C1(new_n522), .C2(new_n507), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n518), .A2(new_n523), .ZN(G168));
  AND2_X1   g099(.A1(new_n505), .A2(new_n506), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n506), .A2(G543), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT72), .B(G52), .Z(new_n527));
  AOI22_X1  g102(.A1(G90), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT73), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  INV_X1    g110(.A(G43), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n507), .A2(new_n535), .B1(new_n509), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n531), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT74), .Z(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  XNOR2_X1  g122(.A(new_n505), .B(KEYINPUT75), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n531), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n525), .A2(G91), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n526), .A2(new_n552), .A3(G53), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n552), .B1(new_n526), .B2(G53), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(G299));
  INV_X1    g132(.A(G168), .ZN(G286));
  INV_X1    g133(.A(G166), .ZN(G303));
  OAI21_X1  g134(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n505), .A2(new_n506), .A3(G87), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n506), .A2(G49), .A3(G543), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(G288));
  NAND2_X1  g138(.A1(new_n525), .A2(G86), .ZN(new_n564));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT5), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n565), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n526), .A2(G48), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n564), .A2(new_n573), .A3(new_n574), .ZN(G305));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  INV_X1    g151(.A(G47), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n507), .A2(new_n576), .B1(new_n509), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G72), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G60), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n570), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(G651), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n582), .B(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n570), .B(KEYINPUT75), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(G79), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n507), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n591), .A2(new_n594), .B1(G54), .B2(new_n526), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n590), .A2(KEYINPUT77), .A3(new_n595), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n585), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n585), .B1(new_n600), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  AOI22_X1  g179(.A1(G299), .A2(new_n603), .B1(new_n604), .B2(KEYINPUT78), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(KEYINPUT78), .B2(new_n604), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(KEYINPUT78), .B2(new_n604), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n600), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND3_X1  g184(.A1(new_n598), .A2(new_n608), .A3(new_n599), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g188(.A1(new_n469), .A2(G2104), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT66), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n461), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT12), .Z(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT13), .Z(new_n621));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OR3_X1    g198(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n483), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n481), .A2(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n631));
  OR3_X1    g206(.A1(new_n631), .A2(new_n464), .A3(G111), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n629), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n631), .B1(new_n464), .B2(G111), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n630), .A2(new_n632), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n626), .A2(new_n627), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n622), .B2(new_n623), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n624), .A2(new_n625), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT82), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2435), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  XOR2_X1   g238(.A(new_n660), .B(KEYINPUT85), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n661), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n658), .B(KEYINPUT17), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n661), .B1(KEYINPUT86), .B2(new_n658), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(KEYINPUT86), .B2(new_n658), .ZN(new_n670));
  OAI22_X1  g245(.A1(new_n670), .A2(new_n664), .B1(new_n667), .B2(new_n666), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n663), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n682), .B(KEYINPUT87), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(KEYINPUT20), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n679), .A2(new_n680), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n678), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n678), .A2(new_n681), .A3(new_n689), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n686), .A2(new_n688), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT21), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT22), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT88), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n692), .A2(KEYINPUT21), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n692), .A2(KEYINPUT21), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n699), .A2(KEYINPUT22), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n695), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n698), .B1(new_n695), .B2(new_n701), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n676), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n701), .ZN(new_n706));
  AOI21_X1  g281(.A(KEYINPUT22), .B1(new_n699), .B2(new_n700), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n697), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n708), .A2(new_n675), .A3(new_n702), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(new_n709), .ZN(G229));
  MUX2_X1   g285(.A(G6), .B(G305), .S(G16), .Z(new_n711));
  XOR2_X1   g286(.A(KEYINPUT32), .B(G1981), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n714), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(G1971), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(G1971), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G23), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n713), .A2(new_n717), .A3(new_n718), .A4(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT34), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n582), .B(KEYINPUT76), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(new_n714), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n714), .B2(G24), .ZN(new_n728));
  INV_X1    g303(.A(G1986), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n481), .A2(G119), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n483), .A2(G131), .ZN(new_n734));
  OR2_X1    g309(.A1(G95), .A2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n732), .B1(new_n737), .B2(new_n731), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  XOR2_X1   g314(.A(new_n738), .B(new_n739), .Z(new_n740));
  NOR3_X1   g315(.A1(new_n730), .A2(KEYINPUT89), .A3(new_n740), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n725), .B(new_n741), .C1(new_n729), .C2(new_n728), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT36), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n714), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n714), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT99), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1961), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n731), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n731), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT29), .Z(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n714), .A2(G20), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT100), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT23), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n556), .B2(new_n714), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT101), .B(G1956), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n751), .A2(G2090), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n756), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n481), .A2(G129), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n483), .A2(G141), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n461), .A2(G105), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT26), .Z(new_n765));
  NAND4_X1  g340(.A1(new_n761), .A2(new_n762), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n760), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT27), .B(G1996), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT95), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n768), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n714), .A2(G19), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n540), .B2(new_n714), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G1341), .Z(new_n774));
  NOR2_X1   g349(.A1(new_n636), .A2(new_n731), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT96), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n731), .B1(new_n779), .B2(G28), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT98), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n780), .A2(new_n781), .B1(new_n779), .B2(G28), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n771), .A2(new_n774), .A3(new_n776), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n714), .A2(G21), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G168), .B2(new_n714), .ZN(new_n787));
  INV_X1    g362(.A(G1966), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n751), .B2(G2090), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n747), .A2(new_n759), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(G104), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT91), .ZN(new_n794));
  INV_X1    g369(.A(G128), .ZN(new_n795));
  INV_X1    g370(.A(G140), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n795), .A2(new_n480), .B1(new_n465), .B2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G29), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT92), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n731), .A2(G26), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT28), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G2067), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G27), .A2(G29), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G164), .B2(G29), .ZN(new_n807));
  INV_X1    g382(.A(G2078), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n791), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT24), .ZN(new_n811));
  INV_X1    g386(.A(G34), .ZN(new_n812));
  AOI21_X1  g387(.A(G29), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G160), .B2(new_n731), .ZN(new_n815));
  INV_X1    g390(.A(G2084), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G2072), .ZN(new_n818));
  OR2_X1    g393(.A1(G29), .A2(G33), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n461), .A2(G103), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT25), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G139), .B2(new_n483), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n618), .A2(G127), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n824));
  NAND2_X1  g399(.A1(G115), .A2(G2104), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G2105), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n819), .B1(new_n829), .B2(new_n731), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n817), .B1(new_n818), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n714), .A2(G4), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n600), .B2(new_n714), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT90), .Z(new_n834));
  AOI21_X1  g409(.A(new_n831), .B1(new_n834), .B2(G1348), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(new_n818), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT94), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n835), .B(new_n837), .C1(G1348), .C2(new_n834), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n743), .A2(new_n810), .A3(new_n838), .ZN(G311));
  OR3_X1    g414(.A1(new_n743), .A2(new_n838), .A3(new_n810), .ZN(G150));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n507), .A2(new_n841), .B1(new_n509), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n505), .A2(G67), .ZN(new_n844));
  NAND2_X1  g419(.A1(G80), .A2(G543), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n531), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT104), .B(G860), .Z(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n598), .A2(new_n599), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n608), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n843), .A2(new_n846), .A3(KEYINPUT102), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT102), .B1(new_n843), .B2(new_n846), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n856), .A2(new_n540), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n540), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT39), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n849), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n855), .A2(new_n861), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n851), .B1(new_n863), .B2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n487), .B(KEYINPUT105), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n829), .A2(KEYINPUT106), .A3(new_n766), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n766), .B1(new_n829), .B2(KEYINPUT106), .ZN(new_n869));
  OAI21_X1  g444(.A(G164), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n500), .A2(new_n503), .ZN(new_n872));
  INV_X1    g447(.A(new_n495), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(new_n874), .A3(new_n867), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n875), .A3(new_n798), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n620), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n481), .A2(G130), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n483), .A2(G142), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n737), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n885), .A2(new_n879), .A3(new_n880), .A4(new_n882), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n884), .B2(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n878), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n886), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT107), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n620), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n890), .A2(new_n894), .A3(KEYINPUT108), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT108), .B1(new_n890), .B2(new_n894), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n798), .B1(new_n870), .B2(new_n875), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n877), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n895), .B1(new_n900), .B2(new_n876), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n866), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n478), .B(new_n636), .Z(new_n903));
  OAI211_X1 g478(.A(new_n900), .B(new_n876), .C1(new_n895), .C2(new_n896), .ZN(new_n904));
  INV_X1    g479(.A(new_n895), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n877), .B2(new_n898), .ZN(new_n906));
  INV_X1    g481(.A(new_n866), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n903), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n903), .B1(new_n902), .B2(new_n908), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT40), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n909), .A4(new_n910), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(G395));
  NAND3_X1  g492(.A1(new_n600), .A2(new_n608), .A3(new_n860), .ZN(new_n918));
  INV_X1    g493(.A(new_n860), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n610), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n556), .A2(new_n596), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n590), .B(new_n595), .C1(new_n550), .C2(new_n555), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n924), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n922), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n921), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(G305), .B(KEYINPUT111), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n726), .ZN(new_n937));
  NAND2_X1  g512(.A1(G290), .A2(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(G166), .B(new_n720), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(KEYINPUT42), .A3(new_n943), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n921), .B(KEYINPUT110), .C1(new_n929), .C2(new_n931), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n918), .A2(new_n920), .A3(new_n925), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n934), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n948), .ZN(new_n954));
  INV_X1    g529(.A(new_n928), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT41), .B1(new_n923), .B2(new_n924), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT109), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n957), .A2(new_n930), .B1(new_n918), .B2(new_n920), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n950), .B1(new_n958), .B2(KEYINPUT110), .ZN(new_n959));
  INV_X1    g534(.A(new_n949), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n954), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n950), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n932), .B2(new_n933), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n963), .A2(KEYINPUT112), .A3(new_n949), .A4(new_n948), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n953), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G868), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n847), .A2(G868), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n965), .B2(G868), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n967), .B2(new_n970), .ZN(G295));
  OAI21_X1  g546(.A(new_n968), .B1(new_n967), .B2(new_n970), .ZN(G331));
  NAND2_X1  g547(.A1(G171), .A2(G286), .ZN(new_n973));
  NAND2_X1  g548(.A1(G301), .A2(G168), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n919), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n860), .A3(new_n974), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n957), .A2(new_n930), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n925), .A3(new_n977), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n944), .ZN(new_n982));
  AOI21_X1  g557(.A(G37), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n944), .B1(new_n978), .B2(new_n980), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT43), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n976), .A2(new_n977), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n955), .A2(new_n956), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n979), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(G37), .B1(new_n988), .B2(new_n944), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n981), .A2(new_n982), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT43), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT44), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n983), .B2(new_n984), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n992), .B1(new_n996), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g572(.A(KEYINPUT114), .B(G40), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT115), .B1(new_n477), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n464), .B1(new_n474), .B2(new_n475), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n1002));
  NOR4_X1   g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n467), .A4(new_n998), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G164), .B2(G1384), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n798), .B(G2067), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1009), .A2(KEYINPUT116), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n737), .B(new_n739), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n766), .B(G1996), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1009), .A2(KEYINPUT116), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1010), .A2(new_n1012), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(G290), .B(G1986), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1007), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  INV_X1    g595(.A(new_n467), .ZN(new_n1021));
  INV_X1    g596(.A(new_n475), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n618), .B2(G125), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1021), .B(new_n999), .C1(new_n1023), .C2(new_n464), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1002), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n476), .A2(G2105), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1026), .A2(KEYINPUT115), .A3(new_n1021), .A4(new_n999), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G164), .A2(G1384), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1020), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G86), .ZN(new_n1031));
  INV_X1    g606(.A(G48), .ZN(new_n1032));
  OAI22_X1  g607(.A1(new_n507), .A2(new_n1031), .B1(new_n509), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n505), .A2(G61), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n531), .B1(new_n1034), .B2(new_n565), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n573), .A2(new_n564), .A3(new_n574), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1038), .A3(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1019), .B1(new_n1030), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1384), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n874), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1048));
  NOR4_X1   g623(.A1(new_n1048), .A2(new_n1043), .A3(KEYINPUT121), .A4(new_n1020), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G288), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1030), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1051), .B1(new_n720), .B2(G1976), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT120), .B(new_n1051), .C1(new_n720), .C2(G1976), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1050), .A2(KEYINPUT52), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NOR4_X1   g637(.A1(new_n1048), .A2(new_n1062), .A3(new_n1020), .A4(new_n1054), .ZN(new_n1063));
  OAI22_X1  g638(.A1(new_n1045), .A2(new_n1049), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(G166), .B2(new_n1020), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1065), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n531), .B1(new_n513), .B2(new_n514), .ZN(new_n1068));
  OAI211_X1 g643(.A(G8), .B(new_n1067), .C1(new_n1068), .C2(new_n511), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G2090), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n874), .A2(new_n1072), .A3(new_n1046), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1028), .A2(new_n1071), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n874), .A2(KEYINPUT45), .A3(new_n1046), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1006), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1004), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1075), .B1(new_n1078), .B2(G1971), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1070), .B1(new_n1079), .B2(G8), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1064), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1070), .B(KEYINPUT118), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1082), .A3(G8), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1028), .A2(new_n808), .A3(new_n1006), .A4(new_n1076), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1073), .B(new_n1074), .C1(new_n1000), .C2(new_n1003), .ZN(new_n1088));
  INV_X1    g663(.A(G1961), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT45), .B1(new_n874), .B2(new_n1046), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1005), .B(G1384), .C1(new_n872), .C2(new_n873), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(KEYINPUT53), .A3(new_n808), .A4(new_n1028), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1087), .A2(G301), .A3(new_n1090), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n808), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n477), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1087), .A2(new_n1099), .A3(new_n1090), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G171), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1085), .A2(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1102), .A2(KEYINPUT125), .A3(G301), .A4(new_n1094), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1097), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT54), .ZN(new_n1105));
  AOI21_X1  g680(.A(G301), .B1(new_n1102), .B2(new_n1094), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(KEYINPUT54), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(G171), .B2(new_n1100), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1956), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1088), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1093), .A2(new_n1028), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n556), .A2(KEYINPUT57), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n550), .B2(new_n555), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1111), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1348), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1088), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1048), .A2(new_n804), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n852), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1120), .A2(new_n852), .A3(new_n1121), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT60), .B1(new_n1125), .B2(new_n1122), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1111), .A2(new_n1117), .A3(new_n1113), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1128), .B2(new_n1123), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1117), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1126), .A2(new_n1129), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1028), .A2(new_n1006), .A3(new_n1076), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT58), .B(G1341), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1135), .A2(G1996), .B1(new_n1048), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n540), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(KEYINPUT59), .A3(new_n540), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1120), .A2(new_n600), .A3(new_n1142), .A4(new_n1121), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1124), .B1(new_n1134), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G168), .A2(new_n1020), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1135), .A2(new_n788), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1028), .A2(new_n816), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1149), .B2(G8), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT51), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1146), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1153), .B(G8), .C1(new_n1149), .C2(G286), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1109), .A2(new_n1145), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(KEYINPUT62), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1151), .A2(new_n1158), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(new_n1106), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1084), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT63), .ZN(new_n1163));
  OAI21_X1  g738(.A(G168), .B1(new_n1162), .B2(KEYINPUT63), .ZN(new_n1164));
  AOI211_X1 g739(.A(new_n1020), .B(new_n1164), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1081), .A2(new_n1083), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1029), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(G8), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT121), .B1(new_n1168), .B2(new_n1043), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1030), .A2(new_n1019), .A3(new_n1044), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1167), .A2(G8), .A3(new_n1055), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1052), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1062), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1030), .A2(new_n1055), .A3(new_n1174), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1169), .A2(new_n1170), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1075), .ZN(new_n1177));
  AOI21_X1  g752(.A(G1971), .B1(new_n1093), .B2(new_n1028), .ZN(new_n1178));
  OAI21_X1  g753(.A(G8), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1070), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1176), .A2(new_n1181), .A3(new_n1083), .A4(new_n1165), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1163), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(G288), .A2(G1976), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT122), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1038), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1083), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1188), .A2(new_n1030), .B1(new_n1189), .B2(new_n1176), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1166), .A2(new_n1184), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1166), .A2(new_n1184), .A3(new_n1190), .A4(KEYINPUT124), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1018), .B1(new_n1161), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1010), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n737), .A2(new_n739), .ZN(new_n1198));
  OAI22_X1  g773(.A1(new_n1197), .A2(new_n1198), .B1(G2067), .B2(new_n798), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1007), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1016), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1007), .A2(new_n729), .A3(new_n726), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1016), .A2(new_n1201), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1007), .B1(new_n766), .B2(new_n1008), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT126), .ZN(new_n1208));
  OR3_X1    g783(.A1(new_n1004), .A2(G1996), .A3(new_n1006), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT46), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  AND2_X1   g786(.A1(new_n1211), .A2(KEYINPUT47), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1211), .A2(KEYINPUT47), .ZN(new_n1213));
  OAI221_X1 g788(.A(new_n1200), .B1(new_n1205), .B2(new_n1206), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1196), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g791(.A1(new_n911), .A2(new_n912), .ZN(new_n1218));
  NOR2_X1   g792(.A1(G227), .A2(new_n458), .ZN(new_n1219));
  AND2_X1   g793(.A1(new_n656), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g794(.A1(new_n705), .A2(new_n709), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g795(.A(new_n1221), .B1(new_n994), .B2(new_n995), .ZN(new_n1222));
  NOR2_X1   g796(.A1(new_n1218), .A2(new_n1222), .ZN(G308));
  OAI221_X1 g797(.A(new_n1221), .B1(new_n994), .B2(new_n995), .C1(new_n911), .C2(new_n912), .ZN(G225));
endmodule


