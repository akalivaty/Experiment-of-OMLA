//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n202), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(new_n208), .A2(new_n209), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n215), .B1(new_n209), .B2(new_n208), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT2), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G226), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(G50), .B(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G13), .ZN(new_n241));
  NOR2_X1   g0041(.A1(new_n241), .A2(G1), .ZN(new_n242));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n242), .A2(G20), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT12), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  AOI22_X1  g0046(.A1(new_n246), .A2(G50), .B1(G20), .B2(new_n243), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G20), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n212), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n254), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G68), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n245), .A2(new_n255), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT11), .B1(new_n252), .B2(new_n254), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G169), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT67), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT67), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n271), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n275), .A2(new_n277), .B1(G238), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G226), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(G232), .A3(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G97), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT13), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT13), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n283), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n265), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT14), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(G179), .A3(new_n297), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n298), .B2(new_n299), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n264), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n295), .A2(new_n297), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n295), .A2(new_n308), .A3(new_n297), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n264), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT78), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n253), .A2(new_n212), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n250), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT72), .ZN(new_n317));
  NAND2_X1  g0117(.A1(KEYINPUT8), .A2(G58), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT8), .A2(G58), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(KEYINPUT8), .A2(G58), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT72), .A3(new_n318), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n323), .A3(new_n246), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G20), .A2(G77), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n316), .B1(new_n326), .B2(KEYINPUT73), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT73), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n324), .A2(new_n328), .A3(new_n325), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n314), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n257), .A2(G77), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT74), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n259), .A2(G77), .A3(new_n260), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT75), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n275), .A2(new_n277), .B1(G244), .B2(new_n282), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n286), .A2(G232), .ZN(new_n338));
  INV_X1    g0138(.A(G107), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n338), .A2(G1698), .B1(new_n339), .B2(new_n286), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n287), .B1(new_n284), .B2(new_n285), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT68), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(new_n342), .B2(G238), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n337), .B1(new_n343), .B2(new_n279), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G200), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT75), .ZN(new_n346));
  INV_X1    g0146(.A(new_n335), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n324), .A2(new_n328), .A3(new_n325), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n328), .B1(new_n324), .B2(new_n325), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n348), .A2(new_n349), .A3(new_n316), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n346), .B(new_n347), .C1(new_n350), .C2(new_n314), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n336), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT76), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n336), .A2(new_n345), .A3(new_n351), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n337), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n342), .A2(G238), .ZN(new_n357));
  INV_X1    g0157(.A(new_n340), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n356), .B1(new_n359), .B2(new_n292), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G190), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n353), .A2(new_n355), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT69), .B(G58), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n320), .B1(new_n363), .B2(KEYINPUT8), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n257), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n364), .A2(new_n260), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n259), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n246), .ZN(new_n369));
  INV_X1    g0169(.A(G159), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n363), .A2(G68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n202), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n373), .B2(G20), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n284), .A2(new_n213), .A3(new_n285), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(KEYINPUT3), .A2(G33), .ZN(new_n378));
  NOR2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT7), .B1(new_n380), .B2(new_n213), .ZN(new_n381));
  OAI21_X1  g0181(.A(G68), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n374), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n201), .B1(new_n363), .B2(G68), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n385), .A2(new_n213), .B1(new_n370), .B2(new_n369), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n375), .A2(new_n376), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n380), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n243), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT16), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n368), .B1(new_n391), .B2(new_n254), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n282), .A2(G232), .ZN(new_n393));
  INV_X1    g0193(.A(new_n277), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n276), .B1(new_n271), .B2(new_n273), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n341), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n286), .A2(G223), .A3(new_n287), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n279), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n306), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n341), .A2(G226), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n292), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n275), .A2(new_n277), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(new_n393), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n400), .B1(new_n406), .B2(G190), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n392), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(G169), .B1(new_n396), .B2(new_n399), .ZN(new_n411));
  AND2_X1   g0211(.A1(KEYINPUT71), .A2(G179), .ZN(new_n412));
  NOR2_X1   g0212(.A1(KEYINPUT71), .A2(G179), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n404), .A2(new_n405), .A3(new_n414), .A4(new_n393), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n314), .B1(new_n384), .B2(new_n390), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n416), .B(new_n417), .C1(new_n418), .C2(new_n368), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n416), .B1(new_n418), .B2(new_n368), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT18), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n407), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n410), .A2(new_n419), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n336), .A2(new_n351), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n414), .B(new_n337), .C1(new_n343), .C2(new_n279), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n360), .B2(new_n265), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n362), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n313), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G223), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n286), .A2(G222), .A3(new_n287), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n251), .B2(new_n286), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n292), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n275), .A2(new_n277), .B1(G226), .B2(new_n282), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(G190), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n306), .B1(new_n437), .B2(new_n438), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT10), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n364), .A2(new_n249), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT70), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n246), .A2(G150), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n254), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G50), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n256), .B2(G20), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n259), .A2(new_n453), .B1(new_n452), .B2(new_n258), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT9), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n451), .A2(KEYINPUT9), .A3(new_n454), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n442), .A2(new_n443), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT77), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n441), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n462), .A2(new_n458), .A3(new_n439), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(KEYINPUT77), .A3(new_n443), .A4(new_n457), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n443), .B1(new_n463), .B2(new_n457), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n437), .A2(new_n438), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G169), .ZN(new_n470));
  INV_X1    g0270(.A(new_n414), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n455), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n430), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT20), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n213), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  INV_X1    g0279(.A(G97), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(G33), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n481), .B2(new_n213), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n476), .B1(new_n482), .B2(new_n314), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n248), .A2(G97), .ZN(new_n484));
  AOI21_X1  g0284(.A(G20), .B1(new_n484), .B2(new_n479), .ZN(new_n485));
  OAI211_X1 g0285(.A(KEYINPUT20), .B(new_n254), .C1(new_n485), .C2(new_n478), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n256), .A2(G33), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n314), .A2(new_n257), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n257), .A2(new_n477), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(G264), .B(G1698), .C1(new_n378), .C2(new_n379), .ZN(new_n494));
  OAI211_X1 g0294(.A(G257), .B(new_n287), .C1(new_n378), .C2(new_n379), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n284), .A2(G303), .A3(new_n285), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n292), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n266), .A2(G1), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(G274), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G41), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G270), .A3(new_n279), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT84), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT84), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n505), .A2(new_n508), .A3(G270), .A4(new_n279), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n498), .A2(new_n501), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n493), .A2(new_n510), .A3(KEYINPUT21), .A4(G169), .ZN(new_n511));
  INV_X1    g0311(.A(new_n212), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n499), .A2(new_n500), .B1(new_n512), .B2(new_n278), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n508), .B1(new_n513), .B2(G270), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n509), .A2(new_n501), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n493), .A2(G179), .A3(new_n516), .A4(new_n498), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n510), .A2(new_n306), .ZN(new_n519));
  INV_X1    g0319(.A(new_n515), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n520), .A2(new_n308), .A3(new_n498), .A4(new_n507), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n493), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n265), .B1(new_n487), .B2(new_n492), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT21), .B1(new_n523), .B2(new_n510), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n518), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G244), .B(G1698), .C1(new_n378), .C2(new_n379), .ZN(new_n526));
  OAI211_X1 g0326(.A(G238), .B(new_n287), .C1(new_n378), .C2(new_n379), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G116), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n292), .ZN(new_n530));
  OAI21_X1  g0330(.A(G250), .B1(new_n266), .B2(G1), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n273), .A2(G45), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n292), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(G190), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT83), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(new_n529), .B2(new_n292), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT83), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(G190), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n286), .A2(new_n213), .A3(G68), .ZN(new_n541));
  INV_X1    g0341(.A(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G87), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G97), .A2(G107), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n213), .B1(new_n290), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n290), .B2(G20), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n541), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n254), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n315), .A2(new_n258), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n259), .A2(G87), .A3(new_n488), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n537), .A2(new_n306), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n553), .B(new_n554), .C1(new_n315), .C2(new_n489), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n530), .A2(new_n414), .A3(new_n534), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n265), .B2(new_n537), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n540), .A2(new_n558), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n213), .A2(G107), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n242), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n564), .B(KEYINPUT25), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n489), .A2(new_n339), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT23), .B1(new_n213), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n213), .A2(G33), .A3(G116), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT85), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n339), .A2(G20), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(KEYINPUT23), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT23), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n574), .A2(new_n339), .A3(KEYINPUT85), .A4(G20), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n570), .A2(KEYINPUT86), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT86), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n568), .A3(new_n569), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT85), .B1(new_n563), .B2(new_n574), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n213), .B(G87), .C1(new_n378), .C2(new_n379), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n582), .B(KEYINPUT22), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(KEYINPUT24), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n254), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT24), .B1(new_n581), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n567), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G250), .B(new_n287), .C1(new_n378), .C2(new_n379), .ZN(new_n588));
  OAI211_X1 g0388(.A(G257), .B(G1698), .C1(new_n378), .C2(new_n379), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n292), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n513), .A2(G264), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n501), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G169), .ZN(new_n595));
  INV_X1    g0395(.A(G179), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n594), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n587), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n306), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n591), .A2(new_n292), .B1(new_n513), .B2(G264), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(new_n308), .A3(new_n501), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n602), .B(new_n567), .C1(new_n586), .C2(new_n585), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n525), .A2(new_n562), .A3(new_n598), .A4(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(G107), .B1(new_n377), .B2(new_n381), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT6), .ZN(new_n606));
  AND2_X1   g0406(.A1(G97), .A2(G107), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n546), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n339), .A2(KEYINPUT6), .A3(G97), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(G20), .B1(G77), .B2(new_n246), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n314), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n258), .A2(new_n480), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n489), .B2(new_n480), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n612), .A2(KEYINPUT81), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT81), .ZN(new_n616));
  INV_X1    g0416(.A(new_n609), .ZN(new_n617));
  XNOR2_X1  g0417(.A(G97), .B(G107), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n606), .B2(new_n618), .ZN(new_n619));
  OAI22_X1  g0419(.A1(new_n619), .A2(new_n213), .B1(new_n251), .B2(new_n369), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n339), .B1(new_n387), .B2(new_n388), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n254), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n614), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n616), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT4), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(G1698), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(G244), .C1(new_n379), .C2(new_n378), .ZN(new_n628));
  INV_X1    g0428(.A(G244), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n284), .B2(new_n285), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n628), .B(new_n479), .C1(new_n630), .C2(KEYINPUT4), .ZN(new_n631));
  OAI21_X1  g0431(.A(G250), .B1(new_n378), .B2(new_n379), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n287), .B1(new_n632), .B2(KEYINPUT4), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT79), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(KEYINPUT4), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G1698), .ZN(new_n636));
  OAI21_X1  g0436(.A(G244), .B1(new_n378), .B2(new_n379), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n626), .B1(G33), .B2(G283), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT79), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n636), .A2(new_n638), .A3(new_n639), .A4(new_n628), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n634), .A2(new_n640), .A3(new_n292), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT80), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT80), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n634), .A2(new_n640), .A3(new_n643), .A4(new_n292), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n513), .A2(G257), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n501), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n642), .A2(new_n471), .A3(new_n644), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n641), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n265), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n625), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n646), .B1(new_n641), .B2(KEYINPUT80), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n306), .B1(new_n652), .B2(new_n644), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n612), .A2(new_n614), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n649), .B2(new_n308), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n651), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n604), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n475), .A2(new_n657), .ZN(G372));
  AOI22_X1  g0458(.A1(new_n558), .A2(new_n535), .B1(new_n559), .B2(new_n561), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n603), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT87), .B1(new_n518), .B2(new_n524), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n523), .A2(new_n510), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT21), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT87), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n511), .A4(new_n517), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n660), .B1(new_n667), .B2(new_n598), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n625), .A2(new_n648), .A3(new_n650), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n653), .A2(new_n655), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n561), .A2(new_n559), .ZN(new_n673));
  INV_X1    g0473(.A(new_n654), .ZN(new_n674));
  AND4_X1   g0474(.A1(new_n674), .A2(new_n659), .A3(new_n648), .A4(new_n650), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n562), .A2(new_n648), .A3(new_n625), .A4(new_n650), .ZN(new_n676));
  XOR2_X1   g0476(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n677));
  OAI22_X1  g0477(.A1(new_n675), .A2(KEYINPUT26), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n475), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n473), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n421), .A2(new_n419), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n298), .A2(new_n299), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(new_n300), .A3(new_n302), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n428), .B1(new_n684), .B2(new_n264), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n407), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT17), .B1(new_n392), .B2(new_n407), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n311), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n682), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n681), .B1(new_n690), .B2(new_n468), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n680), .A2(new_n691), .ZN(G369));
  INV_X1    g0492(.A(new_n598), .ZN(new_n693));
  INV_X1    g0493(.A(new_n242), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .A3(G20), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT27), .B1(new_n694), .B2(G20), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n518), .A2(new_n524), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n699), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT90), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n703), .A2(KEYINPUT90), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n587), .A2(new_n699), .ZN(new_n708));
  INV_X1    g0508(.A(new_n603), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n598), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n701), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n701), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT89), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n493), .A2(new_n699), .ZN(new_n715));
  OR3_X1    g0515(.A1(new_n667), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n667), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n525), .A2(new_n715), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n711), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G330), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n713), .A2(new_n721), .ZN(G399));
  OR2_X1    g0522(.A1(new_n547), .A2(G116), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT91), .ZN(new_n724));
  INV_X1    g0524(.A(new_n207), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n724), .A2(new_n256), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n211), .B2(new_n726), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT28), .Z(new_n729));
  INV_X1    g0529(.A(KEYINPUT95), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n679), .A2(new_n700), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT93), .ZN(new_n732));
  INV_X1    g0532(.A(new_n673), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n668), .B2(new_n671), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n699), .B1(new_n734), .B2(new_n678), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n732), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n675), .A2(KEYINPUT26), .B1(new_n676), .B2(new_n677), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n660), .B1(new_n702), .B2(new_n598), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n733), .B1(new_n671), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n699), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n641), .A2(new_n647), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n600), .A2(new_n537), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n748), .A2(new_n510), .A3(new_n596), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n747), .A2(KEYINPUT30), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT30), .B1(new_n747), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n642), .A2(new_n644), .A3(new_n647), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(KEYINPUT92), .A3(new_n594), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n414), .B(new_n537), .C1(new_n516), .C2(new_n498), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(KEYINPUT92), .B1(new_n753), .B2(new_n594), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT31), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n758), .A2(new_n759), .A3(new_n699), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(new_n657), .B2(new_n700), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(new_n699), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G330), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n730), .B1(new_n746), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n746), .A2(new_n730), .A3(new_n764), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n729), .B1(new_n768), .B2(G1), .ZN(G364));
  NOR2_X1   g0569(.A1(new_n241), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n256), .B1(new_n770), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OR3_X1    g0572(.A1(new_n726), .A2(new_n772), .A3(KEYINPUT96), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT96), .B1(new_n726), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n719), .A2(G330), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n719), .A2(G330), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n719), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n306), .A2(G179), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(G20), .A3(G190), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n543), .B2(new_n545), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G179), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G190), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n380), .B(new_n787), .C1(G97), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n308), .A2(new_n306), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n414), .A2(G20), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n791), .B1(new_n452), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n213), .A2(G190), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n788), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n370), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n414), .A2(G200), .A3(new_n795), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n414), .A2(new_n306), .A3(new_n795), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n243), .B2(new_n800), .C1(new_n251), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n795), .A2(new_n785), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT100), .Z(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n471), .A2(new_n213), .A3(new_n308), .A4(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n363), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n339), .A2(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n794), .A2(new_n802), .A3(new_n809), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT101), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT101), .ZN(new_n812));
  INV_X1    g0612(.A(new_n796), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n286), .B1(new_n813), .B2(G329), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n786), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G294), .B2(new_n790), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G283), .A2(new_n804), .B1(new_n806), .B2(G322), .ZN(new_n818));
  INV_X1    g0618(.A(new_n801), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G311), .ZN(new_n820));
  INV_X1    g0620(.A(new_n793), .ZN(new_n821));
  INV_X1    g0621(.A(new_n800), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT33), .B(G317), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G326), .A2(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n817), .A2(new_n818), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n811), .A2(new_n812), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n212), .B1(G20), .B2(new_n265), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n782), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n725), .A2(new_n380), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(G355), .B1(new_n477), .B2(new_n725), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT97), .Z(new_n831));
  NAND2_X1  g0631(.A1(new_n380), .A2(new_n207), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT98), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n267), .A2(new_n269), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n236), .A2(new_n266), .B1(new_n210), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n831), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n826), .A2(new_n827), .B1(new_n828), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n775), .B1(new_n784), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n779), .A2(new_n840), .ZN(G396));
  NOR2_X1   g0641(.A1(new_n827), .A2(new_n780), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n775), .B1(new_n251), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n827), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G137), .A2(new_n821), .B1(new_n819), .B2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G150), .ZN(new_n846));
  INV_X1    g0646(.A(G143), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n845), .B1(new_n846), .B2(new_n800), .C1(new_n847), .C2(new_n807), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT34), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n380), .B1(new_n813), .B2(G132), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n452), .B2(new_n786), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n805), .A2(new_n243), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(new_n363), .C2(new_n790), .ZN(new_n853));
  INV_X1    g0653(.A(new_n790), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n380), .B1(new_n786), .B2(new_n339), .C1(new_n854), .C2(new_n480), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G283), .A2(new_n822), .B1(new_n821), .B2(G303), .ZN(new_n856));
  INV_X1    g0656(.A(G294), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n807), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n855), .B(new_n858), .C1(G116), .C2(new_n819), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n804), .A2(G87), .ZN(new_n860));
  INV_X1    g0660(.A(G311), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n861), .B2(new_n796), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT102), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n849), .A2(new_n853), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n428), .A2(new_n699), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT103), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n427), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n424), .A2(new_n699), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT103), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n865), .B1(new_n870), .B2(new_n362), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n843), .B1(new_n844), .B2(new_n864), .C1(new_n871), .C2(new_n781), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n679), .A2(new_n871), .A3(new_n700), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n732), .A2(new_n737), .ZN(new_n875));
  INV_X1    g0675(.A(new_n871), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n764), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n776), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n877), .A2(new_n878), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n872), .B1(new_n880), .B2(new_n881), .ZN(G384));
  NAND3_X1  g0682(.A1(new_n211), .A2(new_n372), .A3(G77), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n883), .A2(KEYINPUT105), .B1(G50), .B2(new_n243), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n883), .A2(KEYINPUT105), .ZN(new_n885));
  OAI211_X1 g0685(.A(G1), .B(new_n241), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(G116), .B(new_n214), .C1(new_n610), .C2(KEYINPUT35), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(KEYINPUT35), .B2(new_n610), .ZN(new_n888));
  XOR2_X1   g0688(.A(KEYINPUT104), .B(KEYINPUT36), .Z(new_n889));
  XNOR2_X1  g0689(.A(new_n888), .B(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  INV_X1    g0691(.A(new_n697), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n418), .B2(new_n368), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n682), .B2(new_n688), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n408), .A2(new_n420), .A3(new_n893), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n408), .A2(KEYINPUT37), .A3(new_n420), .A4(new_n893), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n891), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n893), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n423), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n897), .A4(new_n898), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n353), .A2(new_n355), .A3(new_n361), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n905), .A2(new_n868), .A3(new_n867), .A4(new_n869), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n264), .B(new_n699), .C1(new_n684), .C2(new_n310), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n264), .A2(new_n699), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n304), .A2(new_n311), .A3(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n865), .A2(new_n906), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n598), .A2(new_n562), .A3(new_n603), .ZN(new_n911));
  INV_X1    g0711(.A(new_n522), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n912), .A2(new_n664), .A3(new_n511), .A4(new_n517), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n671), .A2(new_n914), .A3(new_n700), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n762), .A2(new_n915), .A3(KEYINPUT31), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n758), .A2(new_n759), .A3(new_n699), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n904), .A2(new_n910), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT107), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT107), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n918), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n920), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n475), .A2(new_n763), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(G330), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n904), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n900), .A2(new_n903), .A3(KEYINPUT39), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n684), .A2(new_n264), .A3(new_n700), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n682), .A2(new_n892), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n907), .A2(new_n909), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n867), .A2(new_n869), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n700), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n939), .B1(new_n873), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n904), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n739), .A2(new_n475), .A3(new_n745), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n691), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n929), .A2(new_n947), .B1(new_n256), .B2(new_n770), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT108), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n929), .A2(new_n947), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n886), .B(new_n890), .C1(new_n950), .C2(new_n952), .ZN(G367));
  AOI22_X1  g0753(.A1(new_n806), .A2(G303), .B1(G311), .B2(new_n821), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT113), .Z(new_n955));
  NOR2_X1   g0755(.A1(new_n786), .A2(new_n477), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT46), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G107), .B2(new_n790), .ZN(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n380), .B1(new_n796), .B2(new_n959), .C1(new_n480), .C2(new_n803), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n800), .A2(new_n857), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(G283), .C2(new_n819), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n854), .A2(new_n243), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n806), .B2(G150), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n847), .B2(new_n793), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT114), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  INV_X1    g0769(.A(G137), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n286), .B1(new_n796), .B2(new_n970), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n808), .A2(new_n786), .B1(new_n803), .B2(new_n251), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(G159), .C2(new_n822), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n969), .B(new_n973), .C1(new_n452), .C2(new_n801), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n963), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT47), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n827), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n833), .A2(new_n232), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n980), .B(new_n828), .C1(new_n207), .C2(new_n315), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT112), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n776), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n982), .B2(new_n981), .ZN(new_n984));
  INV_X1    g0784(.A(new_n659), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n556), .A2(new_n699), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n673), .A2(new_n556), .A3(new_n699), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n979), .B(new_n984), .C1(new_n783), .C2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n674), .A2(new_n699), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n671), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n648), .A2(new_n674), .A3(new_n650), .A4(new_n699), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n995), .B(new_n720), .C1(new_n706), .C2(new_n705), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT42), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT42), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n669), .B1(new_n995), .B2(new_n693), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n997), .B(new_n998), .C1(new_n699), .C2(new_n999), .ZN(new_n1000));
  OR3_X1    g0800(.A1(new_n1000), .A2(KEYINPUT43), .A3(new_n990), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n989), .B(KEYINPUT43), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n1000), .A2(KEYINPUT109), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT109), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n995), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n721), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n721), .A2(new_n1006), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1001), .B(new_n1008), .C1(new_n1004), .C2(new_n1003), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n712), .A2(new_n1011), .A3(new_n1006), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT45), .B1(new_n713), .B2(new_n995), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n712), .A2(new_n1006), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1014), .B1(new_n712), .B2(new_n1006), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n721), .B1(new_n1012), .B2(new_n1013), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n721), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1017), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1019), .B1(new_n1022), .B2(new_n1015), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1013), .A2(new_n1012), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n778), .A2(new_n711), .A3(new_n707), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT111), .B1(new_n707), .B2(new_n711), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n707), .A2(new_n711), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(G330), .A3(new_n719), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1029), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n768), .B1(new_n1026), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n726), .B(KEYINPUT41), .Z(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n772), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n991), .B1(new_n1010), .B2(new_n1038), .ZN(G387));
  INV_X1    g0839(.A(new_n1034), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n767), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1040), .B1(new_n1041), .B2(new_n765), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n766), .A2(new_n767), .A3(new_n1034), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1042), .A2(new_n1043), .A3(new_n726), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n286), .B1(new_n786), .B2(new_n251), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n854), .A2(new_n315), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(G150), .C2(new_n813), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n804), .A2(G97), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G159), .A2(new_n821), .B1(new_n822), .B2(new_n364), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n806), .A2(G50), .B1(G68), .B2(new_n819), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n801), .A2(new_n815), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n807), .A2(new_n959), .B1(new_n861), .B2(new_n800), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(G322), .C2(new_n821), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT48), .ZN(new_n1055));
  INV_X1    g0855(.A(G283), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n854), .A2(new_n1056), .B1(new_n786), .B2(new_n857), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n1054), .B2(KEYINPUT48), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(KEYINPUT49), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n813), .A2(G326), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n803), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n286), .B1(new_n1061), .B2(G116), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT49), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1051), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n827), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n834), .B1(new_n229), .B2(new_n836), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n724), .B2(new_n829), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n321), .A2(new_n323), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1069), .A2(G50), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT50), .Z(new_n1071));
  OAI21_X1  g0871(.A(new_n266), .B1(new_n243), .B2(new_n251), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1071), .A2(new_n724), .A3(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1068), .A2(new_n1073), .B1(G107), .B2(new_n207), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n775), .B1(new_n1074), .B2(new_n828), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1066), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n711), .B2(new_n782), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1040), .B2(new_n772), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1044), .A2(new_n1078), .ZN(G393));
  INV_X1    g0879(.A(new_n726), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1042), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1026), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n772), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n828), .B1(new_n480), .B2(new_n207), .C1(new_n834), .C2(new_n239), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n776), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n806), .A2(G311), .B1(G317), .B2(new_n821), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT52), .Z(new_n1089));
  OAI21_X1  g0889(.A(new_n380), .B1(new_n786), .B2(new_n1056), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G322), .B2(new_n813), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(new_n339), .C2(new_n805), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n822), .A2(G303), .B1(G116), .B2(new_n790), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n857), .B2(new_n801), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT115), .Z(new_n1095));
  AOI22_X1  g0895(.A1(new_n806), .A2(G159), .B1(G150), .B2(new_n821), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n860), .B1(new_n452), .B2(new_n800), .C1(new_n1069), .C2(new_n801), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n854), .A2(new_n251), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n286), .B1(new_n796), .B2(new_n847), .C1(new_n243), .C2(new_n786), .ZN(new_n1100));
  OR3_X1    g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1092), .A2(new_n1095), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1087), .B1(new_n1102), .B2(new_n827), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n995), .B2(new_n783), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1084), .A2(new_n1085), .A3(new_n1104), .ZN(G390));
  INV_X1    g0905(.A(new_n934), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n933), .B1(new_n942), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n906), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n744), .A2(new_n1108), .B1(new_n700), .B2(new_n940), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n904), .B(new_n934), .C1(new_n1109), .C2(new_n939), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n916), .A2(G330), .A3(new_n917), .A4(new_n871), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1112), .A2(new_n939), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n904), .A2(new_n934), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n702), .A2(new_n598), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n603), .A3(new_n659), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n673), .B1(new_n1117), .B2(new_n656), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n700), .B1(new_n1118), .B2(new_n740), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n941), .B1(new_n1119), .B2(new_n906), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1115), .B1(new_n938), .B2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n735), .A2(new_n871), .B1(new_n700), .B2(new_n940), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n934), .B1(new_n1122), .B2(new_n939), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n933), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n763), .A2(G330), .A3(new_n871), .A4(new_n938), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT116), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT116), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1111), .A2(new_n1127), .A3(new_n1113), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1114), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n933), .A2(new_n780), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n842), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n776), .B1(new_n364), .B2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n806), .A2(G132), .B1(G137), .B2(new_n822), .ZN(new_n1133));
  INV_X1    g0933(.A(G125), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n286), .B1(new_n796), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G50), .B2(new_n1061), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1133), .B(new_n1136), .C1(new_n370), .C2(new_n854), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n786), .A2(new_n846), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  INV_X1    g0939(.A(G128), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n793), .C1(new_n801), .C2(new_n1141), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n380), .B1(new_n796), .B2(new_n857), .C1(new_n542), .C2(new_n786), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(new_n1099), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n339), .B2(new_n800), .C1(new_n805), .C2(new_n243), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G97), .A2(new_n819), .B1(new_n821), .B2(G283), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n477), .B2(new_n807), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1137), .A2(new_n1142), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1132), .B1(new_n1148), .B2(new_n827), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1129), .A2(new_n772), .B1(new_n1130), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1112), .A2(new_n939), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1125), .A2(new_n1109), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT117), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1112), .A2(new_n1153), .A3(new_n939), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1112), .B2(new_n939), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1125), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1122), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1152), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n475), .A2(G330), .A3(new_n763), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n945), .A2(new_n691), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT118), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1125), .A2(new_n1109), .A3(new_n1151), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1151), .A2(KEYINPUT117), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1112), .A2(new_n1153), .A3(new_n939), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1113), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1162), .B1(new_n1165), .B2(new_n1122), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT118), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n945), .A2(new_n691), .A3(new_n1159), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT119), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1161), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(new_n1129), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n726), .B1(new_n1171), .B2(new_n1129), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1150), .B1(new_n1172), .B2(new_n1173), .ZN(G378));
  NOR3_X1   g0974(.A1(new_n1158), .A2(KEYINPUT118), .A3(new_n1160), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1167), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1129), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1168), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n918), .A2(new_n919), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n918), .A2(new_n924), .A3(new_n921), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n924), .B1(new_n918), .B2(new_n921), .ZN(new_n1181));
  OAI211_X1 g0981(.A(G330), .B(new_n1179), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1183));
  INV_X1    g0983(.A(KEYINPUT121), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n468), .A2(new_n1184), .A3(new_n473), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n466), .B1(new_n461), .B2(new_n464), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT121), .B1(new_n1186), .B2(new_n681), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n455), .A2(new_n892), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1185), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1189), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1183), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1188), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1183), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1190), .A3(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1182), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n923), .A2(new_n925), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(new_n1201), .A3(G330), .A4(new_n1179), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT123), .B1(new_n937), .B2(new_n943), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1199), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT57), .B1(new_n1178), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1161), .A2(new_n1169), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1160), .B1(new_n1208), .B2(new_n1129), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n944), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1199), .A2(new_n1202), .A3(new_n944), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(KEYINPUT57), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n726), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1207), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1198), .A2(new_n780), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n776), .B1(G50), .B2(new_n1131), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n806), .A2(G107), .B1(G97), .B2(new_n822), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n477), .B2(new_n793), .C1(new_n315), .C2(new_n801), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n808), .A2(new_n803), .B1(new_n786), .B2(new_n251), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n270), .B(new_n380), .C1(new_n796), .C2(new_n1056), .ZN(new_n1222));
  OR4_X1    g1022(.A1(new_n964), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT58), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G50), .B1(new_n248), .B2(new_n270), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n286), .B2(G41), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT120), .Z(new_n1229));
  NAND2_X1  g1029(.A1(new_n790), .A2(G150), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n786), .B2(new_n1141), .C1(new_n793), .C2(new_n1134), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n807), .A2(new_n1140), .B1(new_n970), .B2(new_n801), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(G132), .C2(new_n822), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n248), .B(new_n270), .C1(new_n803), .C2(new_n370), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G124), .B2(new_n813), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT59), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1237), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1229), .B1(new_n1224), .B2(new_n1223), .C1(new_n1235), .C2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1218), .B1(new_n1240), .B2(new_n827), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1217), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT122), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1242), .B(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n772), .B2(new_n1206), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1216), .A2(new_n1245), .ZN(G375));
  OAI21_X1  g1046(.A(new_n776), .B1(G68), .B2(new_n1131), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n786), .A2(new_n370), .B1(new_n796), .B2(new_n1140), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n286), .B1(new_n808), .B2(new_n803), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(G50), .C2(new_n790), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n800), .A2(new_n1141), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n806), .B2(G137), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G132), .A2(new_n821), .B1(new_n819), .B2(G150), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n286), .B1(new_n804), .B2(G77), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT124), .Z(new_n1256));
  OAI22_X1  g1056(.A1(new_n786), .A2(new_n480), .B1(new_n796), .B2(new_n815), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1257), .B(new_n1046), .C1(G294), .C2(new_n821), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n806), .A2(G283), .B1(G116), .B2(new_n822), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(new_n339), .C2(new_n801), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1254), .B1(new_n1256), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1247), .B1(new_n1261), .B2(new_n827), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n938), .B2(new_n781), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1158), .B2(new_n771), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1161), .A2(new_n1169), .A3(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1265), .B1(new_n1267), .B2(new_n1036), .ZN(G381));
  INV_X1    g1068(.A(new_n1150), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1161), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1127), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1272));
  AOI211_X1 g1072(.A(KEYINPUT116), .B(new_n1125), .C1(new_n1107), .C2(new_n1110), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1080), .B1(new_n1270), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1171), .A2(new_n1129), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1269), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1216), .A2(new_n1277), .A3(new_n1245), .ZN(new_n1278));
  INV_X1    g1078(.A(G390), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n991), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n771), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1280), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(G384), .ZN(new_n1285));
  INV_X1    g1085(.A(G396), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1044), .A2(new_n1286), .A3(new_n1078), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1279), .A2(new_n1284), .A3(new_n1285), .A4(new_n1288), .ZN(new_n1289));
  OR3_X1    g1089(.A1(new_n1278), .A2(G381), .A3(new_n1289), .ZN(G407));
  NAND2_X1  g1090(.A1(new_n698), .A2(G213), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1291), .B(KEYINPUT125), .Z(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G407), .B(G213), .C1(new_n1278), .C2(new_n1293), .ZN(G409));
  OAI211_X1 g1094(.A(G378), .B(new_n1245), .C1(new_n1207), .C2(new_n1215), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1274), .B1(new_n1169), .B2(new_n1161), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1037), .B(new_n1206), .C1(new_n1296), .C2(new_n1160), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1199), .A2(new_n1202), .A3(new_n944), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n944), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1300), .A2(new_n772), .B1(new_n1217), .B2(new_n1241), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1277), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1295), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1267), .A2(KEYINPUT60), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n726), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1305), .A2(new_n1306), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1265), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1309), .B1(new_n1267), .B2(KEYINPUT60), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1313), .A2(new_n1306), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1285), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1264), .B1(new_n1313), .B2(new_n1306), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT126), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1316), .A2(new_n1318), .A3(G384), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1304), .A2(new_n1293), .A3(new_n1315), .A4(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT62), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1304), .A2(new_n1293), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1312), .A2(new_n1314), .A3(new_n1285), .ZN(new_n1323));
  AOI21_X1  g1123(.A(G384), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1324));
  OAI211_X1 g1124(.A(G2897), .B(new_n1292), .C1(new_n1323), .C2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1292), .A2(G2897), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1315), .A2(new_n1319), .A3(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1322), .A2(new_n1325), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1292), .B1(new_n1295), .B2(new_n1303), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT62), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1330), .A2(new_n1331), .A3(new_n1332), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1321), .A2(new_n1328), .A3(new_n1329), .A4(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1286), .B1(new_n1044), .B2(new_n1078), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  AND3_X1   g1136(.A1(G387), .A2(new_n1287), .A3(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  AOI22_X1  g1138(.A1(G387), .A2(new_n1338), .B1(new_n1336), .B2(new_n1287), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1279), .B1(new_n1337), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  OAI22_X1  g1141(.A1(new_n1284), .A2(KEYINPUT127), .B1(new_n1288), .B2(new_n1335), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(G387), .A2(new_n1287), .A3(new_n1336), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(G390), .A3(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1341), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1334), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(KEYINPUT61), .B1(new_n1340), .B2(new_n1344), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1330), .A2(KEYINPUT63), .A3(new_n1332), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT63), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1326), .B1(new_n1315), .B2(new_n1319), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1330), .A2(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1351), .B1(new_n1353), .B2(new_n1327), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1320), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1350), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1347), .A2(new_n1356), .ZN(G405));
  OAI22_X1  g1157(.A1(new_n1345), .A2(new_n1341), .B1(new_n1324), .B2(new_n1323), .ZN(new_n1358));
  XNOR2_X1  g1158(.A(G375), .B(new_n1277), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1340), .A2(new_n1332), .A3(new_n1344), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1358), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1359), .B1(new_n1358), .B2(new_n1360), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1361), .A2(new_n1362), .ZN(G402));
endmodule


