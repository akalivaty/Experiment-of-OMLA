

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  XNOR2_X1 U324 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U325 ( .A(KEYINPUT38), .B(n457), .ZN(n502) );
  XOR2_X1 U326 ( .A(n381), .B(n380), .Z(n534) );
  XOR2_X1 U327 ( .A(n401), .B(n374), .Z(n292) );
  NOR2_X1 U328 ( .A1(n480), .A2(n520), .ZN(n293) );
  INV_X1 U329 ( .A(G176GAT), .ZN(n371) );
  INV_X1 U330 ( .A(KEYINPUT103), .ZN(n394) );
  XNOR2_X1 U331 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n476) );
  INV_X1 U332 ( .A(KEYINPUT4), .ZN(n333) );
  XNOR2_X1 U333 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U334 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U335 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U336 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U337 ( .A(n336), .B(n335), .ZN(n340) );
  XNOR2_X1 U338 ( .A(n434), .B(n433), .ZN(n576) );
  NOR2_X1 U339 ( .A1(n534), .A2(n482), .ZN(n563) );
  INV_X1 U340 ( .A(n504), .ZN(n550) );
  XOR2_X1 U341 ( .A(n348), .B(n347), .Z(n520) );
  INV_X1 U342 ( .A(G43GAT), .ZN(n461) );
  XNOR2_X1 U343 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U344 ( .A(n461), .B(KEYINPUT40), .ZN(n462) );
  XNOR2_X1 U345 ( .A(n486), .B(n485), .ZN(G1349GAT) );
  XNOR2_X1 U346 ( .A(n463), .B(n462), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n295) );
  XNOR2_X1 U348 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U350 ( .A(G169GAT), .B(n296), .Z(n381) );
  XOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .Z(n402) );
  XOR2_X1 U352 ( .A(n402), .B(KEYINPUT98), .Z(n298) );
  NAND2_X1 U353 ( .A1(G226GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U355 ( .A(G92GAT), .B(G64GAT), .Z(n300) );
  XNOR2_X1 U356 ( .A(G204GAT), .B(KEYINPUT78), .ZN(n299) );
  XNOR2_X1 U357 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U358 ( .A(G176GAT), .B(n301), .Z(n429) );
  XOR2_X1 U359 ( .A(n302), .B(n429), .Z(n307) );
  XOR2_X1 U360 ( .A(KEYINPUT21), .B(G218GAT), .Z(n304) );
  XNOR2_X1 U361 ( .A(KEYINPUT92), .B(G211GAT), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U363 ( .A(G197GAT), .B(n305), .Z(n363) );
  XNOR2_X1 U364 ( .A(G8GAT), .B(n363), .ZN(n306) );
  XNOR2_X1 U365 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U366 ( .A(n381), .B(n308), .Z(n522) );
  INV_X1 U367 ( .A(n522), .ZN(n508) );
  XOR2_X1 U368 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n456) );
  XOR2_X1 U369 ( .A(KEYINPUT87), .B(KEYINPUT12), .Z(n310) );
  XNOR2_X1 U370 ( .A(KEYINPUT83), .B(KEYINPUT14), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n310), .B(n309), .ZN(n328) );
  XOR2_X1 U372 ( .A(G22GAT), .B(G155GAT), .Z(n360) );
  XOR2_X1 U373 ( .A(n360), .B(G78GAT), .Z(n312) );
  XOR2_X1 U374 ( .A(G15GAT), .B(G127GAT), .Z(n367) );
  XNOR2_X1 U375 ( .A(n367), .B(G211GAT), .ZN(n311) );
  XNOR2_X1 U376 ( .A(n312), .B(n311), .ZN(n324) );
  XOR2_X1 U377 ( .A(KEYINPUT84), .B(G64GAT), .Z(n314) );
  XNOR2_X1 U378 ( .A(G183GAT), .B(G71GAT), .ZN(n313) );
  XNOR2_X1 U379 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U380 ( .A(KEYINPUT15), .B(KEYINPUT86), .Z(n316) );
  XNOR2_X1 U381 ( .A(KEYINPUT82), .B(KEYINPUT85), .ZN(n315) );
  XNOR2_X1 U382 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U383 ( .A(n318), .B(n317), .Z(n322) );
  XNOR2_X1 U384 ( .A(G1GAT), .B(KEYINPUT72), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n319), .B(G8GAT), .ZN(n446) );
  XNOR2_X1 U386 ( .A(G57GAT), .B(KEYINPUT75), .ZN(n320) );
  XNOR2_X1 U387 ( .A(n320), .B(KEYINPUT13), .ZN(n431) );
  XNOR2_X1 U388 ( .A(n446), .B(n431), .ZN(n321) );
  XNOR2_X1 U389 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U390 ( .A(n324), .B(n323), .Z(n326) );
  NAND2_X1 U391 ( .A1(G231GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U392 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U393 ( .A(n328), .B(n327), .Z(n580) );
  XOR2_X1 U394 ( .A(G134GAT), .B(KEYINPUT81), .Z(n401) );
  XNOR2_X1 U395 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n329) );
  XNOR2_X1 U396 ( .A(n329), .B(KEYINPUT88), .ZN(n374) );
  NAND2_X1 U397 ( .A1(G225GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U398 ( .A(n292), .B(n330), .ZN(n336) );
  XOR2_X1 U399 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n332) );
  XNOR2_X1 U400 ( .A(G141GAT), .B(KEYINPUT93), .ZN(n331) );
  XNOR2_X1 U401 ( .A(n332), .B(n331), .ZN(n353) );
  XNOR2_X1 U402 ( .A(n353), .B(KEYINPUT5), .ZN(n334) );
  XOR2_X1 U403 ( .A(G85GAT), .B(G155GAT), .Z(n338) );
  XNOR2_X1 U404 ( .A(G29GAT), .B(G162GAT), .ZN(n337) );
  XOR2_X1 U405 ( .A(n338), .B(n337), .Z(n339) );
  XNOR2_X1 U406 ( .A(n340), .B(n339), .ZN(n348) );
  XOR2_X1 U407 ( .A(KEYINPUT97), .B(KEYINPUT1), .Z(n342) );
  XNOR2_X1 U408 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U410 ( .A(G57GAT), .B(G148GAT), .Z(n344) );
  XNOR2_X1 U411 ( .A(G127GAT), .B(G120GAT), .ZN(n343) );
  XNOR2_X1 U412 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U414 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n350) );
  NAND2_X1 U415 ( .A1(G228GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U417 ( .A(n351), .B(KEYINPUT96), .Z(n355) );
  XNOR2_X1 U418 ( .A(G106GAT), .B(G78GAT), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n352), .B(G148GAT), .ZN(n430) );
  XNOR2_X1 U420 ( .A(n353), .B(n430), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U422 ( .A(G204GAT), .B(KEYINPUT22), .Z(n357) );
  XNOR2_X1 U423 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n356) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U425 ( .A(n359), .B(n358), .Z(n362) );
  XOR2_X1 U426 ( .A(G50GAT), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U427 ( .A(n409), .B(n360), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U429 ( .A(n364), .B(n363), .Z(n480) );
  XOR2_X1 U430 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n366) );
  XNOR2_X1 U431 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n379) );
  XOR2_X1 U433 ( .A(G190GAT), .B(G134GAT), .Z(n369) );
  XOR2_X1 U434 ( .A(G120GAT), .B(G71GAT), .Z(n422) );
  XNOR2_X1 U435 ( .A(n367), .B(n422), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U437 ( .A(n370), .B(G99GAT), .Z(n377) );
  NAND2_X1 U438 ( .A1(G227GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U439 ( .A(G43GAT), .B(n375), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U441 ( .A(n379), .B(n378), .Z(n380) );
  NOR2_X1 U442 ( .A1(n534), .A2(n508), .ZN(n382) );
  NOR2_X1 U443 ( .A1(n480), .A2(n382), .ZN(n383) );
  XOR2_X1 U444 ( .A(KEYINPUT25), .B(n383), .Z(n386) );
  XOR2_X1 U445 ( .A(KEYINPUT27), .B(n522), .Z(n388) );
  NAND2_X1 U446 ( .A1(n480), .A2(n534), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n384), .B(KEYINPUT26), .ZN(n568) );
  NOR2_X1 U448 ( .A1(n388), .A2(n568), .ZN(n385) );
  NOR2_X1 U449 ( .A1(n386), .A2(n385), .ZN(n387) );
  NOR2_X1 U450 ( .A1(n520), .A2(n387), .ZN(n393) );
  INV_X1 U451 ( .A(n520), .ZN(n569) );
  NOR2_X1 U452 ( .A1(n569), .A2(n388), .ZN(n532) );
  XNOR2_X1 U453 ( .A(n480), .B(KEYINPUT28), .ZN(n537) );
  INV_X1 U454 ( .A(n537), .ZN(n513) );
  NAND2_X1 U455 ( .A1(n532), .A2(n513), .ZN(n389) );
  XNOR2_X1 U456 ( .A(KEYINPUT99), .B(n389), .ZN(n390) );
  NAND2_X1 U457 ( .A1(n390), .A2(n534), .ZN(n391) );
  XOR2_X1 U458 ( .A(KEYINPUT100), .B(n391), .Z(n392) );
  NOR2_X1 U459 ( .A1(n393), .A2(n392), .ZN(n490) );
  NOR2_X1 U460 ( .A1(n580), .A2(n490), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n417) );
  XOR2_X1 U462 ( .A(KEYINPUT8), .B(KEYINPUT71), .Z(n397) );
  XNOR2_X1 U463 ( .A(G43GAT), .B(G29GAT), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U465 ( .A(KEYINPUT7), .B(n398), .ZN(n451) );
  INV_X1 U466 ( .A(n451), .ZN(n415) );
  XOR2_X1 U467 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n400) );
  XNOR2_X1 U468 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n413) );
  XOR2_X1 U470 ( .A(n402), .B(n401), .Z(n404) );
  XNOR2_X1 U471 ( .A(G218GAT), .B(G106GAT), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U473 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n406) );
  NAND2_X1 U474 ( .A1(G232GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U476 ( .A(n408), .B(n407), .Z(n411) );
  XOR2_X1 U477 ( .A(G99GAT), .B(G85GAT), .Z(n421) );
  XNOR2_X1 U478 ( .A(n409), .B(n421), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U480 ( .A(n413), .B(n412), .Z(n414) );
  XOR2_X1 U481 ( .A(n415), .B(n414), .Z(n487) );
  INV_X1 U482 ( .A(n487), .ZN(n562) );
  XOR2_X1 U483 ( .A(KEYINPUT36), .B(KEYINPUT102), .Z(n416) );
  XOR2_X1 U484 ( .A(n562), .B(n416), .Z(n583) );
  NAND2_X1 U485 ( .A1(n417), .A2(n583), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n418), .B(KEYINPUT37), .ZN(n517) );
  XOR2_X1 U487 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n420) );
  XNOR2_X1 U488 ( .A(KEYINPUT32), .B(KEYINPUT79), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n420), .B(n419), .ZN(n426) );
  XOR2_X1 U490 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n424) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U492 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U493 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n430), .B(n429), .ZN(n432) );
  INV_X1 U497 ( .A(n576), .ZN(n471) );
  XOR2_X1 U498 ( .A(G15GAT), .B(G113GAT), .Z(n436) );
  XNOR2_X1 U499 ( .A(G169GAT), .B(G197GAT), .ZN(n435) );
  XNOR2_X1 U500 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U501 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n438) );
  XNOR2_X1 U502 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n437) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U504 ( .A(n440), .B(n439), .Z(n445) );
  XOR2_X1 U505 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n442) );
  NAND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U508 ( .A(KEYINPUT68), .B(n443), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n450) );
  XOR2_X1 U510 ( .A(G36GAT), .B(G50GAT), .Z(n448) );
  XNOR2_X1 U511 ( .A(G22GAT), .B(n446), .ZN(n447) );
  XNOR2_X1 U512 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U513 ( .A(n450), .B(n449), .Z(n453) );
  XOR2_X1 U514 ( .A(n451), .B(G141GAT), .Z(n452) );
  XNOR2_X1 U515 ( .A(n453), .B(n452), .ZN(n571) );
  NAND2_X1 U516 ( .A1(n471), .A2(n571), .ZN(n454) );
  XOR2_X1 U517 ( .A(KEYINPUT80), .B(n454), .Z(n491) );
  NAND2_X1 U518 ( .A1(n517), .A2(n491), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U520 ( .A1(n508), .A2(n502), .ZN(n460) );
  INV_X1 U521 ( .A(G36GAT), .ZN(n458) );
  XNOR2_X1 U522 ( .A(n458), .B(KEYINPUT106), .ZN(n459) );
  XNOR2_X1 U523 ( .A(n460), .B(n459), .ZN(G1329GAT) );
  NOR2_X1 U524 ( .A1(n534), .A2(n502), .ZN(n463) );
  XOR2_X1 U525 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n465) );
  XNOR2_X1 U526 ( .A(n576), .B(KEYINPUT41), .ZN(n504) );
  NAND2_X1 U527 ( .A1(n571), .A2(n550), .ZN(n464) );
  XOR2_X1 U528 ( .A(n465), .B(n464), .Z(n466) );
  NOR2_X1 U529 ( .A1(n580), .A2(n466), .ZN(n467) );
  NAND2_X1 U530 ( .A1(n467), .A2(n487), .ZN(n468) );
  XNOR2_X1 U531 ( .A(n468), .B(KEYINPUT47), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n580), .A2(n583), .ZN(n470) );
  XNOR2_X1 U533 ( .A(KEYINPUT67), .B(KEYINPUT45), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n473), .A2(n571), .ZN(n474) );
  NOR2_X1 U537 ( .A1(n475), .A2(n474), .ZN(n477) );
  XOR2_X1 U538 ( .A(n478), .B(KEYINPUT114), .Z(n533) );
  AND2_X1 U539 ( .A1(n522), .A2(n533), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT54), .ZN(n570) );
  AND2_X1 U541 ( .A1(n570), .A2(n293), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(KEYINPUT55), .ZN(n482) );
  NAND2_X1 U543 ( .A1(n563), .A2(n550), .ZN(n486) );
  XOR2_X1 U544 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n484) );
  XOR2_X1 U545 ( .A(G176GAT), .B(KEYINPUT119), .Z(n483) );
  NAND2_X1 U546 ( .A1(n487), .A2(n580), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT16), .B(n488), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n505) );
  NAND2_X1 U549 ( .A1(n505), .A2(n491), .ZN(n498) );
  NOR2_X1 U550 ( .A1(n569), .A2(n498), .ZN(n493) );
  XNOR2_X1 U551 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NOR2_X1 U554 ( .A1(n508), .A2(n498), .ZN(n495) );
  XOR2_X1 U555 ( .A(G8GAT), .B(n495), .Z(G1325GAT) );
  NOR2_X1 U556 ( .A1(n534), .A2(n498), .ZN(n497) );
  XNOR2_X1 U557 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(G1326GAT) );
  NOR2_X1 U559 ( .A1(n513), .A2(n498), .ZN(n499) );
  XOR2_X1 U560 ( .A(G22GAT), .B(n499), .Z(G1327GAT) );
  NOR2_X1 U561 ( .A1(n569), .A2(n502), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n513), .A2(n502), .ZN(n503) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  NOR2_X1 U566 ( .A1(n571), .A2(n504), .ZN(n518) );
  NAND2_X1 U567 ( .A1(n518), .A2(n505), .ZN(n512) );
  NOR2_X1 U568 ( .A1(n569), .A2(n512), .ZN(n506) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n506), .Z(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT42), .B(n507), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n508), .A2(n512), .ZN(n510) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n534), .A2(n512), .ZN(n511) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n511), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n515) );
  XNOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n519), .B(KEYINPUT109), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n528), .A2(n520), .ZN(n521) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT110), .ZN(n524) );
  NAND2_X1 U585 ( .A1(n522), .A2(n528), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n524), .B(n523), .ZN(G1337GAT) );
  XOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT111), .Z(n527) );
  INV_X1 U588 ( .A(n534), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n528), .A2(n525), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n527), .B(n526), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n530) );
  NAND2_X1 U592 ( .A1(n528), .A2(n537), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n531), .Z(G1339GAT) );
  NAND2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n548) );
  NOR2_X1 U596 ( .A1(n534), .A2(n548), .ZN(n535) );
  XNOR2_X1 U597 ( .A(n535), .B(KEYINPUT115), .ZN(n536) );
  NOR2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n544), .A2(n571), .ZN(n538) );
  XNOR2_X1 U600 ( .A(n538), .B(KEYINPUT116), .ZN(n539) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U603 ( .A1(n544), .A2(n550), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U605 ( .A1(n544), .A2(n580), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n546) );
  NAND2_X1 U609 ( .A1(n544), .A2(n562), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n568), .A2(n548), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n571), .A2(n556), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U616 ( .A1(n556), .A2(n550), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n556), .A2(n580), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n562), .A2(n556), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n563), .A2(n571), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n563), .A2(n580), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n560), .B(KEYINPUT120), .ZN(n561) );
  XOR2_X1 U630 ( .A(KEYINPUT58), .B(n561), .Z(n565) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT122), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(n567), .Z(n573) );
  INV_X1 U636 ( .A(n568), .ZN(n584) );
  AND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n585) );
  AND2_X1 U638 ( .A1(n584), .A2(n585), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n581), .A2(n571), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n575) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n575), .B(n574), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n576), .A2(n581), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(KEYINPUT123), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n588) );
  AND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(G218GAT), .B(n589), .Z(G1355GAT) );
endmodule

