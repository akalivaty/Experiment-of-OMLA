

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790;

  NAND2_X1 U370 ( .A1(n422), .A2(n419), .ZN(n367) );
  BUF_X1 U371 ( .A(n686), .Z(n347) );
  XNOR2_X1 U372 ( .A(n460), .B(n459), .ZN(n491) );
  XNOR2_X2 U373 ( .A(n606), .B(KEYINPUT1), .ZN(n563) );
  INV_X1 U374 ( .A(n367), .ZN(n363) );
  XNOR2_X2 U375 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n498) );
  NOR2_X2 U376 ( .A1(n712), .A2(G953), .ZN(n714) );
  XOR2_X2 U377 ( .A(KEYINPUT85), .B(KEYINPUT35), .Z(n356) );
  INV_X1 U378 ( .A(G953), .ZN(n781) );
  INV_X2 U379 ( .A(n688), .ZN(n569) );
  XNOR2_X2 U380 ( .A(KEYINPUT41), .B(n594), .ZN(n706) );
  AND2_X2 U381 ( .A1(n674), .A2(n374), .ZN(n594) );
  NOR2_X1 U382 ( .A1(n789), .A2(n788), .ZN(n614) );
  NAND2_X1 U383 ( .A1(n370), .A2(n432), .ZN(n369) );
  AND2_X1 U384 ( .A1(n441), .A2(n354), .ZN(n440) );
  XNOR2_X1 U385 ( .A(n614), .B(n613), .ZN(n426) );
  NOR2_X1 U386 ( .A1(n677), .A2(n615), .ZN(n374) );
  OR2_X1 U387 ( .A1(n731), .A2(n449), .ZN(n593) );
  XNOR2_X1 U388 ( .A(n731), .B(n733), .ZN(n734) );
  XNOR2_X1 U389 ( .A(n720), .B(KEYINPUT59), .ZN(n721) );
  XNOR2_X1 U390 ( .A(n464), .B(n463), .ZN(n764) );
  XNOR2_X1 U391 ( .A(n491), .B(KEYINPUT16), .ZN(n464) );
  INV_X1 U392 ( .A(n730), .ZN(n348) );
  INV_X1 U393 ( .A(n348), .ZN(n349) );
  AND2_X2 U394 ( .A1(n404), .A2(n434), .ZN(n730) );
  BUF_X1 U395 ( .A(n726), .Z(n350) );
  XNOR2_X2 U396 ( .A(n517), .B(n487), .ZN(n495) );
  XNOR2_X1 U397 ( .A(G137), .B(G140), .ZN(n506) );
  XNOR2_X1 U398 ( .A(G146), .B(G125), .ZN(n505) );
  XNOR2_X1 U399 ( .A(KEYINPUT66), .B(G101), .ZN(n472) );
  NOR2_X1 U400 ( .A1(n409), .A2(n408), .ZN(n407) );
  NAND2_X1 U401 ( .A1(n416), .A2(n414), .ZN(n408) );
  AND2_X1 U402 ( .A1(n731), .A2(n592), .ZN(n409) );
  INV_X1 U403 ( .A(KEYINPUT19), .ZN(n414) );
  AND2_X1 U404 ( .A1(n412), .A2(KEYINPUT19), .ZN(n411) );
  XNOR2_X1 U405 ( .A(n508), .B(n383), .ZN(n513) );
  XNOR2_X1 U406 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n383) );
  AND2_X1 U407 ( .A1(n423), .A2(n424), .ZN(n365) );
  NAND2_X1 U408 ( .A1(n426), .A2(n425), .ZN(n368) );
  INV_X1 U409 ( .A(n666), .ZN(n424) );
  INV_X1 U410 ( .A(G134), .ZN(n486) );
  NAND2_X1 U411 ( .A1(n477), .A2(n590), .ZN(n418) );
  NAND2_X1 U412 ( .A1(n384), .A2(n439), .ZN(n691) );
  NOR2_X1 U413 ( .A1(G953), .A2(G237), .ZN(n537) );
  XNOR2_X1 U414 ( .A(G122), .B(KEYINPUT100), .ZN(n531) );
  XOR2_X1 U415 ( .A(G140), .B(G104), .Z(n541) );
  INV_X1 U416 ( .A(G104), .ZN(n459) );
  XNOR2_X1 U417 ( .A(G107), .B(KEYINPUT77), .ZN(n489) );
  XNOR2_X1 U418 ( .A(n600), .B(n430), .ZN(n616) );
  INV_X1 U419 ( .A(KEYINPUT71), .ZN(n430) );
  NAND2_X1 U420 ( .A1(G902), .A2(G469), .ZN(n456) );
  INV_X1 U421 ( .A(KEYINPUT0), .ZN(n394) );
  NAND2_X1 U422 ( .A1(n750), .A2(n484), .ZN(n485) );
  XNOR2_X1 U423 ( .A(n764), .B(n471), .ZN(n450) );
  NAND2_X1 U424 ( .A1(n634), .A2(n636), .ZN(n420) );
  AND2_X1 U425 ( .A1(n667), .A2(n665), .ZN(n446) );
  NAND2_X1 U426 ( .A1(n674), .A2(n479), .ZN(n375) );
  INV_X1 U427 ( .A(KEYINPUT108), .ZN(n438) );
  INV_X1 U428 ( .A(G237), .ZN(n475) );
  XNOR2_X1 U429 ( .A(G116), .B(G137), .ZN(n518) );
  INV_X1 U430 ( .A(KEYINPUT101), .ZN(n386) );
  XOR2_X1 U431 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n532) );
  NAND2_X1 U432 ( .A1(n646), .A2(n403), .ZN(n402) );
  NAND2_X1 U433 ( .A1(n439), .A2(n435), .ZN(n605) );
  XNOR2_X1 U434 ( .A(n436), .B(KEYINPUT79), .ZN(n435) );
  NOR2_X1 U435 ( .A1(n437), .A2(n598), .ZN(n436) );
  XNOR2_X1 U436 ( .A(n597), .B(n438), .ZN(n437) );
  NOR2_X1 U437 ( .A1(n417), .A2(n615), .ZN(n416) );
  NOR2_X1 U438 ( .A1(n477), .A2(n590), .ZN(n417) );
  NAND2_X1 U439 ( .A1(n454), .A2(n453), .ZN(n452) );
  INV_X1 U440 ( .A(G469), .ZN(n454) );
  XNOR2_X1 U441 ( .A(n512), .B(n511), .ZN(n564) );
  AND2_X2 U442 ( .A1(n644), .A2(n761), .ZN(n780) );
  NAND2_X1 U443 ( .A1(n359), .A2(n358), .ZN(n357) );
  AND2_X1 U444 ( .A1(n362), .A2(n361), .ZN(n360) );
  INV_X1 U445 ( .A(G107), .ZN(n461) );
  XNOR2_X1 U446 ( .A(G122), .B(G116), .ZN(n462) );
  AND2_X1 U447 ( .A1(n780), .A2(KEYINPUT64), .ZN(n396) );
  XNOR2_X1 U448 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n467) );
  XNOR2_X1 U449 ( .A(KEYINPUT89), .B(KEYINPUT91), .ZN(n468) );
  NOR2_X1 U450 ( .A1(n670), .A2(n672), .ZN(n432) );
  NAND2_X1 U451 ( .A1(n433), .A2(n351), .ZN(n372) );
  INV_X1 U452 ( .A(n626), .ZN(n378) );
  BUF_X1 U453 ( .A(n688), .Z(n389) );
  XNOR2_X1 U454 ( .A(n562), .B(n561), .ZN(n587) );
  XNOR2_X1 U455 ( .A(n388), .B(KEYINPUT62), .ZN(n650) );
  BUF_X1 U456 ( .A(n649), .Z(n388) );
  XNOR2_X1 U457 ( .A(n539), .B(n387), .ZN(n720) );
  XNOR2_X1 U458 ( .A(n542), .B(n538), .ZN(n387) );
  NOR2_X1 U459 ( .A1(n781), .A2(G952), .ZN(n736) );
  NOR2_X1 U460 ( .A1(n616), .A2(n569), .ZN(n429) );
  NAND2_X1 U461 ( .A1(n353), .A2(n413), .ZN(n750) );
  NAND2_X1 U462 ( .A1(n410), .A2(n407), .ZN(n413) );
  AND2_X1 U463 ( .A1(n710), .A2(n709), .ZN(n351) );
  BUF_X1 U464 ( .A(n564), .Z(n686) );
  XNOR2_X1 U465 ( .A(n515), .B(n514), .ZN(n685) );
  INV_X1 U466 ( .A(n564), .ZN(n384) );
  AND2_X1 U467 ( .A1(n560), .A2(n439), .ZN(n352) );
  AND2_X1 U468 ( .A1(n415), .A2(n406), .ZN(n353) );
  AND2_X1 U469 ( .A1(n588), .A2(n739), .ZN(n354) );
  INV_X1 U470 ( .A(G902), .ZN(n453) );
  AND2_X1 U471 ( .A1(n592), .A2(KEYINPUT19), .ZN(n355) );
  INV_X1 U472 ( .A(KEYINPUT86), .ZN(n366) );
  BUF_X1 U473 ( .A(n563), .Z(n584) );
  BUF_X1 U474 ( .A(n682), .Z(n707) );
  OR2_X2 U475 ( .A1(n455), .A2(n451), .ZN(n606) );
  XNOR2_X1 U476 ( .A(n377), .B(n356), .ZN(n572) );
  NOR2_X1 U477 ( .A1(n629), .A2(n679), .ZN(n631) );
  NOR2_X1 U478 ( .A1(n648), .A2(n767), .ZN(n673) );
  NAND2_X1 U479 ( .A1(n360), .A2(n357), .ZN(n644) );
  AND2_X1 U480 ( .A1(n367), .A2(KEYINPUT86), .ZN(n358) );
  INV_X1 U481 ( .A(n364), .ZN(n359) );
  NAND2_X1 U482 ( .A1(n364), .A2(n366), .ZN(n361) );
  NAND2_X1 U483 ( .A1(n363), .A2(n366), .ZN(n362) );
  NAND2_X1 U484 ( .A1(n365), .A2(n368), .ZN(n364) );
  NAND2_X1 U485 ( .A1(n371), .A2(n369), .ZN(n382) );
  INV_X1 U486 ( .A(n671), .ZN(n370) );
  NOR2_X1 U487 ( .A1(n373), .A2(n372), .ZN(n371) );
  AND2_X1 U488 ( .A1(n671), .A2(n672), .ZN(n373) );
  NOR2_X1 U489 ( .A1(n679), .A2(n375), .ZN(n680) );
  XNOR2_X2 U490 ( .A(n548), .B(n376), .ZN(n775) );
  XNOR2_X2 U491 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n376) );
  XNOR2_X2 U492 ( .A(G143), .B(G128), .ZN(n548) );
  NOR2_X2 U493 ( .A1(n572), .A2(KEYINPUT44), .ZN(n559) );
  NAND2_X1 U494 ( .A1(n379), .A2(n378), .ZN(n377) );
  XNOR2_X1 U495 ( .A(n391), .B(n380), .ZN(n379) );
  INV_X1 U496 ( .A(KEYINPUT34), .ZN(n380) );
  XNOR2_X1 U497 ( .A(n381), .B(n589), .ZN(n647) );
  XNOR2_X1 U498 ( .A(n530), .B(n529), .ZN(n682) );
  INV_X1 U499 ( .A(n673), .ZN(n434) );
  NAND2_X1 U500 ( .A1(n444), .A2(n440), .ZN(n381) );
  NAND2_X1 U501 ( .A1(n457), .A2(n456), .ZN(n455) );
  NOR2_X2 U502 ( .A1(n658), .A2(n736), .ZN(n660) );
  NAND2_X1 U503 ( .A1(n382), .A2(n431), .ZN(n711) );
  XNOR2_X1 U504 ( .A(n429), .B(KEYINPUT28), .ZN(n428) );
  NAND2_X1 U505 ( .A1(n563), .A2(n576), .ZN(n390) );
  XNOR2_X2 U506 ( .A(n775), .B(n472), .ZN(n487) );
  XNOR2_X1 U507 ( .A(n534), .B(n385), .ZN(n535) );
  XNOR2_X1 U508 ( .A(n533), .B(n386), .ZN(n385) );
  NAND2_X1 U509 ( .A1(n443), .A2(n446), .ZN(n442) );
  XNOR2_X1 U510 ( .A(n445), .B(KEYINPUT74), .ZN(n444) );
  XNOR2_X1 U511 ( .A(n390), .B(n516), .ZN(n528) );
  NAND2_X1 U512 ( .A1(n682), .A2(n579), .ZN(n391) );
  NAND2_X1 U513 ( .A1(n442), .A2(KEYINPUT44), .ZN(n441) );
  XNOR2_X1 U514 ( .A(n392), .B(n504), .ZN(n507) );
  XNOR2_X1 U515 ( .A(n393), .B(n502), .ZN(n392) );
  INV_X1 U516 ( .A(n501), .ZN(n393) );
  NOR2_X2 U517 ( .A1(n652), .A2(n736), .ZN(n654) );
  NOR2_X2 U518 ( .A1(n723), .A2(n736), .ZN(n724) );
  NOR2_X2 U519 ( .A1(n737), .A2(n736), .ZN(n738) );
  INV_X1 U520 ( .A(n715), .ZN(n443) );
  NAND2_X1 U521 ( .A1(n400), .A2(n399), .ZN(n398) );
  INV_X1 U522 ( .A(n579), .ZN(n574) );
  NAND2_X1 U523 ( .A1(n579), .A2(n352), .ZN(n562) );
  XNOR2_X2 U524 ( .A(n485), .B(n394), .ZN(n579) );
  NAND2_X1 U525 ( .A1(n397), .A2(n395), .ZN(n404) );
  NAND2_X1 U526 ( .A1(n645), .A2(n396), .ZN(n395) );
  NOR2_X1 U527 ( .A1(n401), .A2(n398), .ZN(n397) );
  OR2_X1 U528 ( .A1(n646), .A2(n403), .ZN(n399) );
  OR2_X1 U529 ( .A1(n780), .A2(n402), .ZN(n400) );
  NOR2_X1 U530 ( .A1(n645), .A2(n402), .ZN(n401) );
  INV_X1 U531 ( .A(KEYINPUT64), .ZN(n403) );
  NAND2_X1 U532 ( .A1(n405), .A2(n411), .ZN(n406) );
  NAND2_X1 U533 ( .A1(n731), .A2(n416), .ZN(n405) );
  NAND2_X1 U534 ( .A1(n731), .A2(n355), .ZN(n415) );
  OR2_X1 U535 ( .A1(n731), .A2(n418), .ZN(n410) );
  NAND2_X1 U536 ( .A1(n416), .A2(n418), .ZN(n412) );
  NAND2_X1 U537 ( .A1(n633), .A2(n634), .ZN(n427) );
  NOR2_X1 U538 ( .A1(n421), .A2(n420), .ZN(n419) );
  INV_X1 U539 ( .A(n633), .ZN(n421) );
  INV_X1 U540 ( .A(n426), .ZN(n422) );
  NAND2_X1 U541 ( .A1(n427), .A2(n425), .ZN(n423) );
  INV_X1 U542 ( .A(n636), .ZN(n425) );
  NAND2_X1 U543 ( .A1(n428), .A2(n606), .ZN(n629) );
  NAND2_X1 U544 ( .A1(n673), .A2(n351), .ZN(n431) );
  NAND2_X1 U545 ( .A1(n670), .A2(n672), .ZN(n433) );
  INV_X1 U546 ( .A(n685), .ZN(n439) );
  NAND2_X1 U547 ( .A1(n447), .A2(n446), .ZN(n445) );
  XNOR2_X1 U548 ( .A(n559), .B(n448), .ZN(n447) );
  INV_X1 U549 ( .A(KEYINPUT67), .ZN(n448) );
  XNOR2_X2 U550 ( .A(n776), .B(G146), .ZN(n517) );
  XNOR2_X2 U551 ( .A(n533), .B(n486), .ZN(n776) );
  XNOR2_X2 U552 ( .A(KEYINPUT69), .B(G131), .ZN(n533) );
  INV_X1 U553 ( .A(n590), .ZN(n449) );
  XNOR2_X2 U554 ( .A(n450), .B(n524), .ZN(n731) );
  NOR2_X1 U555 ( .A1(n726), .A2(n452), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n726), .A2(G469), .ZN(n457) );
  XNOR2_X2 U557 ( .A(n495), .B(n494), .ZN(n726) );
  NAND2_X1 U558 ( .A1(n730), .A2(G478), .ZN(n657) );
  XOR2_X1 U559 ( .A(n526), .B(G472), .Z(n458) );
  INV_X1 U560 ( .A(n615), .ZN(n479) );
  INV_X1 U561 ( .A(KEYINPUT46), .ZN(n613) );
  XNOR2_X1 U562 ( .A(n635), .B(KEYINPUT70), .ZN(n636) );
  BUF_X1 U563 ( .A(n775), .Z(n777) );
  INV_X1 U564 ( .A(n592), .ZN(n477) );
  INV_X1 U565 ( .A(KEYINPUT63), .ZN(n653) );
  BUF_X1 U566 ( .A(n572), .Z(n715) );
  XNOR2_X2 U567 ( .A(KEYINPUT90), .B(G110), .ZN(n460) );
  XNOR2_X1 U568 ( .A(n462), .B(n461), .ZN(n553) );
  INV_X1 U569 ( .A(n553), .ZN(n463) );
  NAND2_X1 U570 ( .A1(n781), .A2(G224), .ZN(n465) );
  XNOR2_X1 U571 ( .A(n465), .B(KEYINPUT78), .ZN(n466) );
  XNOR2_X1 U572 ( .A(n466), .B(n505), .ZN(n470) );
  XNOR2_X1 U573 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U574 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U575 ( .A(G119), .B(G113), .ZN(n474) );
  XNOR2_X1 U576 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n473) );
  XNOR2_X1 U577 ( .A(n474), .B(n473), .ZN(n762) );
  XNOR2_X1 U578 ( .A(n487), .B(n762), .ZN(n524) );
  XNOR2_X1 U579 ( .A(G902), .B(KEYINPUT15), .ZN(n590) );
  NAND2_X1 U580 ( .A1(n453), .A2(n475), .ZN(n478) );
  NAND2_X1 U581 ( .A1(n478), .A2(G210), .ZN(n476) );
  XNOR2_X1 U582 ( .A(n476), .B(KEYINPUT92), .ZN(n592) );
  AND2_X1 U583 ( .A1(n478), .A2(G214), .ZN(n615) );
  NAND2_X1 U584 ( .A1(G237), .A2(G234), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n480), .B(KEYINPUT14), .ZN(n481) );
  NAND2_X1 U586 ( .A1(G902), .A2(n481), .ZN(n595) );
  XNOR2_X1 U587 ( .A(G898), .B(KEYINPUT93), .ZN(n770) );
  NAND2_X1 U588 ( .A1(G953), .A2(n770), .ZN(n765) );
  NOR2_X1 U589 ( .A1(n595), .A2(n765), .ZN(n482) );
  NAND2_X1 U590 ( .A1(G952), .A2(n481), .ZN(n703) );
  NOR2_X1 U591 ( .A1(G953), .A2(n703), .ZN(n598) );
  OR2_X1 U592 ( .A1(n482), .A2(n598), .ZN(n483) );
  XNOR2_X1 U593 ( .A(n483), .B(KEYINPUT94), .ZN(n484) );
  NAND2_X1 U594 ( .A1(n781), .A2(G227), .ZN(n488) );
  XNOR2_X1 U595 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U596 ( .A(n490), .B(n506), .ZN(n493) );
  INV_X1 U597 ( .A(n491), .ZN(n492) );
  XNOR2_X1 U598 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U599 ( .A(KEYINPUT76), .B(G110), .Z(n497) );
  XNOR2_X1 U600 ( .A(G128), .B(G119), .ZN(n496) );
  XNOR2_X1 U601 ( .A(n497), .B(n496), .ZN(n502) );
  INV_X1 U602 ( .A(n498), .ZN(n500) );
  XNOR2_X1 U603 ( .A(KEYINPUT95), .B(KEYINPUT81), .ZN(n499) );
  XNOR2_X1 U604 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U605 ( .A1(G234), .A2(n781), .ZN(n503) );
  XOR2_X1 U606 ( .A(KEYINPUT8), .B(n503), .Z(n545) );
  NAND2_X1 U607 ( .A1(G221), .A2(n545), .ZN(n504) );
  XNOR2_X1 U608 ( .A(n505), .B(KEYINPUT10), .ZN(n536) );
  XNOR2_X1 U609 ( .A(n536), .B(n506), .ZN(n779) );
  XNOR2_X1 U610 ( .A(n507), .B(n779), .ZN(n716) );
  NAND2_X1 U611 ( .A1(n716), .A2(n453), .ZN(n512) );
  XOR2_X1 U612 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n510) );
  NAND2_X1 U613 ( .A1(n590), .A2(G234), .ZN(n508) );
  NAND2_X1 U614 ( .A1(G217), .A2(n513), .ZN(n509) );
  XNOR2_X1 U615 ( .A(n510), .B(n509), .ZN(n511) );
  AND2_X1 U616 ( .A1(n513), .A2(G221), .ZN(n515) );
  INV_X1 U617 ( .A(KEYINPUT21), .ZN(n514) );
  INV_X1 U618 ( .A(n691), .ZN(n576) );
  INV_X1 U619 ( .A(KEYINPUT106), .ZN(n516) );
  INV_X1 U620 ( .A(n517), .ZN(n523) );
  NAND2_X1 U621 ( .A1(n537), .A2(G210), .ZN(n519) );
  XNOR2_X1 U622 ( .A(n519), .B(n518), .ZN(n521) );
  XNOR2_X1 U623 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n520) );
  XNOR2_X1 U624 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U625 ( .A(n523), .B(n522), .ZN(n525) );
  XNOR2_X1 U626 ( .A(n524), .B(n525), .ZN(n649) );
  NOR2_X2 U627 ( .A1(n649), .A2(G902), .ZN(n527) );
  INV_X1 U628 ( .A(KEYINPUT99), .ZN(n526) );
  XNOR2_X2 U629 ( .A(n527), .B(n458), .ZN(n688) );
  XNOR2_X2 U630 ( .A(n569), .B(KEYINPUT6), .ZN(n619) );
  NAND2_X1 U631 ( .A1(n528), .A2(n619), .ZN(n530) );
  XNOR2_X1 U632 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n529) );
  XNOR2_X1 U633 ( .A(n532), .B(n531), .ZN(n534) );
  XOR2_X1 U634 ( .A(n536), .B(n535), .Z(n539) );
  NAND2_X1 U635 ( .A1(G214), .A2(n537), .ZN(n538) );
  XNOR2_X1 U636 ( .A(G143), .B(G113), .ZN(n540) );
  XNOR2_X1 U637 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U638 ( .A1(n720), .A2(n453), .ZN(n544) );
  XOR2_X1 U639 ( .A(KEYINPUT13), .B(G475), .Z(n543) );
  XNOR2_X1 U640 ( .A(n544), .B(n543), .ZN(n582) );
  NAND2_X1 U641 ( .A1(G217), .A2(n545), .ZN(n547) );
  XOR2_X1 U642 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n546) );
  XNOR2_X1 U643 ( .A(n547), .B(n546), .ZN(n550) );
  XNOR2_X1 U644 ( .A(n548), .B(KEYINPUT7), .ZN(n549) );
  XNOR2_X1 U645 ( .A(n550), .B(n549), .ZN(n556) );
  XOR2_X1 U646 ( .A(KEYINPUT103), .B(KEYINPUT105), .Z(n552) );
  XNOR2_X1 U647 ( .A(G134), .B(KEYINPUT104), .ZN(n551) );
  XNOR2_X1 U648 ( .A(n552), .B(n551), .ZN(n554) );
  XNOR2_X1 U649 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U650 ( .A(n556), .B(n555), .ZN(n655) );
  NAND2_X1 U651 ( .A1(n655), .A2(n453), .ZN(n557) );
  XNOR2_X1 U652 ( .A(n557), .B(G478), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n582), .A2(n580), .ZN(n558) );
  XOR2_X1 U654 ( .A(KEYINPUT107), .B(n558), .Z(n626) );
  OR2_X1 U655 ( .A1(n582), .A2(n580), .ZN(n677) );
  INV_X1 U656 ( .A(n677), .ZN(n560) );
  XNOR2_X1 U657 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n561) );
  NAND2_X1 U658 ( .A1(n584), .A2(n347), .ZN(n565) );
  NOR2_X1 U659 ( .A1(n619), .A2(n565), .ZN(n566) );
  NAND2_X1 U660 ( .A1(n587), .A2(n566), .ZN(n568) );
  XOR2_X1 U661 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n567) );
  XNOR2_X1 U662 ( .A(n568), .B(n567), .ZN(n667) );
  NAND2_X1 U663 ( .A1(n569), .A2(n347), .ZN(n570) );
  NOR2_X1 U664 ( .A1(n584), .A2(n570), .ZN(n571) );
  NAND2_X1 U665 ( .A1(n587), .A2(n571), .ZN(n665) );
  AND2_X1 U666 ( .A1(n576), .A2(n584), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n573), .A2(n389), .ZN(n696) );
  NOR2_X1 U668 ( .A1(n574), .A2(n696), .ZN(n575) );
  XNOR2_X1 U669 ( .A(n575), .B(KEYINPUT31), .ZN(n757) );
  NAND2_X1 U670 ( .A1(n576), .A2(n606), .ZN(n577) );
  NOR2_X1 U671 ( .A1(n577), .A2(n389), .ZN(n578) );
  NAND2_X1 U672 ( .A1(n579), .A2(n578), .ZN(n742) );
  NAND2_X1 U673 ( .A1(n757), .A2(n742), .ZN(n583) );
  INV_X1 U674 ( .A(n580), .ZN(n581) );
  OR2_X1 U675 ( .A1(n582), .A2(n581), .ZN(n758) );
  AND2_X1 U676 ( .A1(n582), .A2(n581), .ZN(n617) );
  INV_X1 U677 ( .A(n617), .ZN(n754) );
  NAND2_X1 U678 ( .A1(n758), .A2(n754), .ZN(n630) );
  NAND2_X1 U679 ( .A1(n583), .A2(n630), .ZN(n588) );
  INV_X1 U680 ( .A(n584), .ZN(n692) );
  NAND2_X1 U681 ( .A1(n692), .A2(n384), .ZN(n585) );
  NOR2_X1 U682 ( .A1(n585), .A2(n619), .ZN(n586) );
  NAND2_X1 U683 ( .A1(n587), .A2(n586), .ZN(n739) );
  XNOR2_X1 U684 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n589) );
  NAND2_X1 U685 ( .A1(n647), .A2(n449), .ZN(n591) );
  XNOR2_X1 U686 ( .A(n591), .B(KEYINPUT83), .ZN(n645) );
  XNOR2_X2 U687 ( .A(n593), .B(n592), .ZN(n640) );
  XNOR2_X2 U688 ( .A(n640), .B(KEYINPUT38), .ZN(n674) );
  NOR2_X1 U689 ( .A1(G900), .A2(n595), .ZN(n596) );
  NAND2_X1 U690 ( .A1(G953), .A2(n596), .ZN(n597) );
  XOR2_X1 U691 ( .A(n605), .B(KEYINPUT72), .Z(n599) );
  NAND2_X1 U692 ( .A1(n599), .A2(n686), .ZN(n600) );
  NOR2_X1 U693 ( .A1(n706), .A2(n629), .ZN(n601) );
  XNOR2_X1 U694 ( .A(n601), .B(KEYINPUT42), .ZN(n789) );
  NAND2_X1 U695 ( .A1(n688), .A2(n479), .ZN(n604) );
  XNOR2_X1 U696 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n602) );
  XNOR2_X1 U697 ( .A(n602), .B(KEYINPUT110), .ZN(n603) );
  XNOR2_X1 U698 ( .A(n604), .B(n603), .ZN(n609) );
  NOR2_X1 U699 ( .A1(n686), .A2(n605), .ZN(n607) );
  AND2_X1 U700 ( .A1(n606), .A2(n607), .ZN(n608) );
  AND2_X1 U701 ( .A1(n609), .A2(n608), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n627), .A2(n674), .ZN(n610) );
  XNOR2_X1 U703 ( .A(n610), .B(KEYINPUT39), .ZN(n643) );
  AND2_X1 U704 ( .A1(n643), .A2(n617), .ZN(n612) );
  XNOR2_X1 U705 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n611) );
  XNOR2_X1 U706 ( .A(n612), .B(n611), .ZN(n788) );
  NOR2_X1 U707 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U708 ( .A1(n618), .A2(n617), .ZN(n621) );
  INV_X1 U709 ( .A(n619), .ZN(n620) );
  NOR2_X1 U710 ( .A1(n621), .A2(n620), .ZN(n637) );
  INV_X1 U711 ( .A(n640), .ZN(n622) );
  NAND2_X1 U712 ( .A1(n637), .A2(n622), .ZN(n624) );
  XOR2_X1 U713 ( .A(KEYINPUT113), .B(KEYINPUT36), .Z(n623) );
  XNOR2_X1 U714 ( .A(n624), .B(n623), .ZN(n625) );
  NOR2_X1 U715 ( .A1(n625), .A2(n692), .ZN(n662) );
  NOR2_X1 U716 ( .A1(n626), .A2(n640), .ZN(n628) );
  AND2_X1 U717 ( .A1(n628), .A2(n627), .ZN(n661) );
  NOR2_X1 U718 ( .A1(n662), .A2(n661), .ZN(n634) );
  INV_X1 U719 ( .A(n630), .ZN(n679) );
  NAND2_X1 U720 ( .A1(n631), .A2(n750), .ZN(n632) );
  XOR2_X1 U721 ( .A(KEYINPUT47), .B(n632), .Z(n633) );
  INV_X1 U722 ( .A(KEYINPUT48), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n637), .A2(n692), .ZN(n639) );
  XOR2_X1 U724 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n638) );
  XNOR2_X1 U725 ( .A(n639), .B(n638), .ZN(n641) );
  AND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n666) );
  INV_X1 U727 ( .A(n758), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n761) );
  NAND2_X1 U729 ( .A1(n449), .A2(KEYINPUT2), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n780), .A2(KEYINPUT2), .ZN(n648) );
  BUF_X1 U731 ( .A(n647), .Z(n669) );
  INV_X1 U732 ( .A(n669), .ZN(n767) );
  NAND2_X1 U733 ( .A1(n730), .A2(G472), .ZN(n651) );
  XNOR2_X1 U734 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U735 ( .A(n654), .B(n653), .ZN(G57) );
  INV_X1 U736 ( .A(n655), .ZN(n656) );
  XNOR2_X1 U737 ( .A(n657), .B(n656), .ZN(n658) );
  INV_X1 U738 ( .A(KEYINPUT125), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n660), .B(n659), .ZN(G63) );
  XOR2_X1 U740 ( .A(G143), .B(n661), .Z(G45) );
  XOR2_X1 U741 ( .A(G125), .B(KEYINPUT37), .Z(n663) );
  XOR2_X1 U742 ( .A(n663), .B(n662), .Z(G27) );
  XNOR2_X1 U743 ( .A(G110), .B(KEYINPUT116), .ZN(n664) );
  XNOR2_X1 U744 ( .A(n665), .B(n664), .ZN(G12) );
  XOR2_X1 U745 ( .A(G140), .B(n666), .Z(G42) );
  XNOR2_X1 U746 ( .A(n667), .B(G119), .ZN(G21) );
  NOR2_X2 U747 ( .A1(n780), .A2(KEYINPUT2), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(KEYINPUT82), .ZN(n671) );
  NOR2_X1 U749 ( .A1(n669), .A2(KEYINPUT2), .ZN(n670) );
  INV_X1 U750 ( .A(KEYINPUT80), .ZN(n672) );
  NOR2_X1 U751 ( .A1(n674), .A2(n479), .ZN(n675) );
  XOR2_X1 U752 ( .A(KEYINPUT121), .B(n675), .Z(n676) );
  NOR2_X1 U753 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U754 ( .A(n678), .B(KEYINPUT122), .ZN(n681) );
  NOR2_X1 U755 ( .A1(n681), .A2(n680), .ZN(n684) );
  INV_X1 U756 ( .A(n707), .ZN(n683) );
  OR2_X1 U757 ( .A1(n684), .A2(n683), .ZN(n701) );
  AND2_X1 U758 ( .A1(n347), .A2(n685), .ZN(n687) );
  XOR2_X1 U759 ( .A(KEYINPUT49), .B(n687), .Z(n689) );
  NOR2_X1 U760 ( .A1(n689), .A2(n389), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n690), .B(KEYINPUT120), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n693), .B(KEYINPUT50), .ZN(n694) );
  NAND2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U766 ( .A(KEYINPUT51), .B(n698), .ZN(n699) );
  OR2_X1 U767 ( .A1(n706), .A2(n699), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U769 ( .A(n702), .B(KEYINPUT52), .ZN(n705) );
  INV_X1 U770 ( .A(n703), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n710) );
  INV_X1 U772 ( .A(n706), .ZN(n708) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U774 ( .A(n711), .B(KEYINPUT123), .ZN(n712) );
  XNOR2_X1 U775 ( .A(KEYINPUT124), .B(KEYINPUT53), .ZN(n713) );
  XNOR2_X1 U776 ( .A(n714), .B(n713), .ZN(G75) );
  XOR2_X1 U777 ( .A(n715), .B(G122), .Z(G24) );
  NAND2_X1 U778 ( .A1(n349), .A2(G217), .ZN(n718) );
  XOR2_X1 U779 ( .A(n716), .B(KEYINPUT126), .Z(n717) );
  XNOR2_X1 U780 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U781 ( .A1(n719), .A2(n736), .ZN(G66) );
  NAND2_X1 U782 ( .A1(n730), .A2(G475), .ZN(n722) );
  XNOR2_X1 U783 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U784 ( .A(n724), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U785 ( .A1(n349), .A2(G469), .ZN(n728) );
  XOR2_X1 U786 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n725) );
  XNOR2_X1 U787 ( .A(n350), .B(n725), .ZN(n727) );
  XNOR2_X1 U788 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U789 ( .A1(n729), .A2(n736), .ZN(G54) );
  NAND2_X1 U790 ( .A1(n730), .A2(G210), .ZN(n735) );
  XNOR2_X1 U791 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n732) );
  XNOR2_X1 U792 ( .A(n732), .B(KEYINPUT55), .ZN(n733) );
  XNOR2_X1 U793 ( .A(n735), .B(n734), .ZN(n737) );
  XNOR2_X1 U794 ( .A(n738), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U795 ( .A(G101), .B(n739), .ZN(G3) );
  NOR2_X1 U796 ( .A1(n742), .A2(n754), .ZN(n740) );
  XOR2_X1 U797 ( .A(KEYINPUT114), .B(n740), .Z(n741) );
  XNOR2_X1 U798 ( .A(G104), .B(n741), .ZN(G6) );
  NOR2_X1 U799 ( .A1(n742), .A2(n758), .ZN(n746) );
  XOR2_X1 U800 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n744) );
  XNOR2_X1 U801 ( .A(G107), .B(KEYINPUT115), .ZN(n743) );
  XNOR2_X1 U802 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U803 ( .A(n746), .B(n745), .ZN(G9) );
  NOR2_X1 U804 ( .A1(n629), .A2(n758), .ZN(n747) );
  AND2_X1 U805 ( .A1(n747), .A2(n750), .ZN(n749) );
  XNOR2_X1 U806 ( .A(G128), .B(KEYINPUT29), .ZN(n748) );
  XNOR2_X1 U807 ( .A(n749), .B(n748), .ZN(G30) );
  NOR2_X1 U808 ( .A1(n629), .A2(n754), .ZN(n751) );
  AND2_X1 U809 ( .A1(n751), .A2(n750), .ZN(n753) );
  XNOR2_X1 U810 ( .A(G146), .B(KEYINPUT117), .ZN(n752) );
  XNOR2_X1 U811 ( .A(n753), .B(n752), .ZN(G48) );
  NOR2_X1 U812 ( .A1(n754), .A2(n757), .ZN(n755) );
  XOR2_X1 U813 ( .A(KEYINPUT118), .B(n755), .Z(n756) );
  XNOR2_X1 U814 ( .A(G113), .B(n756), .ZN(G15) );
  NOR2_X1 U815 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U816 ( .A(G116), .B(KEYINPUT119), .ZN(n759) );
  XNOR2_X1 U817 ( .A(n760), .B(n759), .ZN(G18) );
  XNOR2_X1 U818 ( .A(G134), .B(n761), .ZN(G36) );
  XOR2_X1 U819 ( .A(G101), .B(n762), .Z(n763) );
  XNOR2_X1 U820 ( .A(n764), .B(n763), .ZN(n766) );
  NAND2_X1 U821 ( .A1(n766), .A2(n765), .ZN(n774) );
  NOR2_X1 U822 ( .A1(n767), .A2(G953), .ZN(n772) );
  NAND2_X1 U823 ( .A1(G953), .A2(G224), .ZN(n768) );
  XOR2_X1 U824 ( .A(KEYINPUT61), .B(n768), .Z(n769) );
  NOR2_X1 U825 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U826 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U827 ( .A(n774), .B(n773), .ZN(G69) );
  XNOR2_X1 U828 ( .A(n776), .B(n777), .ZN(n778) );
  XNOR2_X1 U829 ( .A(n779), .B(n778), .ZN(n783) );
  XNOR2_X1 U830 ( .A(n780), .B(n783), .ZN(n782) );
  NAND2_X1 U831 ( .A1(n782), .A2(n781), .ZN(n787) );
  XOR2_X1 U832 ( .A(G227), .B(n783), .Z(n784) );
  NAND2_X1 U833 ( .A1(n784), .A2(G900), .ZN(n785) );
  NAND2_X1 U834 ( .A1(G953), .A2(n785), .ZN(n786) );
  NAND2_X1 U835 ( .A1(n787), .A2(n786), .ZN(G72) );
  XOR2_X1 U836 ( .A(G131), .B(n788), .Z(G33) );
  XNOR2_X1 U837 ( .A(G137), .B(KEYINPUT127), .ZN(n790) );
  XNOR2_X1 U838 ( .A(n790), .B(n789), .ZN(G39) );
endmodule

