//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT40), .ZN(new_n202));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n203), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G141gat), .B(G148gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n207), .B(new_n206), .C1(new_n211), .C2(KEYINPUT2), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G113gat), .ZN(new_n214));
  INV_X1    g013(.A(G120gat), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT1), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(new_n214), .B2(new_n215), .ZN(new_n217));
  XNOR2_X1  g016(.A(G127gat), .B(G134gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G113gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n216), .B(new_n218), .C1(new_n221), .C2(new_n215), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n213), .A2(KEYINPUT76), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT76), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(new_n222), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n212), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G225gat), .A2(G233gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n226), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n223), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT80), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n225), .A2(new_n226), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(KEYINPUT4), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n223), .A2(new_n227), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(KEYINPUT4), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n226), .A2(KEYINPUT3), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n210), .A2(new_n212), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n238), .A3(new_n225), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT75), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n226), .A2(KEYINPUT3), .B1(new_n220), .B2(new_n222), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT75), .A3(new_n238), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n228), .B1(new_n235), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT39), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n231), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n246), .ZN(new_n248));
  XNOR2_X1  g047(.A(G1gat), .B(G29gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT0), .ZN(new_n250));
  XNOR2_X1  g049(.A(G57gat), .B(G85gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n250), .B(new_n251), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n202), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(G197gat), .A2(G204gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(G197gat), .A2(G204gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(G211gat), .A2(G218gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(KEYINPUT22), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G211gat), .B(G218gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(KEYINPUT71), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  OAI221_X1 g061(.A(new_n257), .B1(KEYINPUT22), .B2(new_n258), .C1(new_n260), .C2(KEYINPUT71), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT72), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT27), .B(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n272), .A2(KEYINPUT66), .A3(new_n277), .A4(new_n273), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(G169gat), .B2(G176gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n281), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n276), .A2(new_n278), .A3(new_n280), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n281), .A2(KEYINPUT23), .ZN(new_n291));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT25), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n294), .A4(new_n292), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n287), .A2(new_n288), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT24), .B1(new_n284), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n300), .B2(new_n284), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n283), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n271), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n302), .A2(new_n299), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n289), .A2(new_n295), .ZN(new_n308));
  OAI22_X1  g107(.A1(new_n307), .A2(new_n298), .B1(new_n308), .B2(KEYINPUT25), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n270), .B1(new_n309), .B2(new_n283), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n269), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(new_n271), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT29), .B1(new_n309), .B2(new_n283), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n312), .B(new_n268), .C1(new_n313), .C2(new_n271), .ZN(new_n314));
  XOR2_X1   g113(.A(G8gat), .B(G36gat), .Z(new_n315));
  XOR2_X1   g114(.A(G64gat), .B(G92gat), .Z(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT73), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n311), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT30), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n311), .A2(new_n314), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n317), .ZN(new_n325));
  INV_X1    g124(.A(new_n317), .ZN(new_n326));
  AOI211_X1 g125(.A(KEYINPUT30), .B(new_n326), .C1(new_n311), .C2(new_n314), .ZN(new_n327));
  OAI22_X1  g126(.A1(new_n321), .A2(new_n322), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n245), .A2(new_n246), .ZN(new_n329));
  INV_X1    g128(.A(new_n231), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n252), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n332), .B1(new_n245), .B2(new_n246), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(KEYINPUT40), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT5), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n223), .A2(new_n227), .A3(new_n229), .ZN(new_n336));
  INV_X1    g135(.A(new_n228), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n239), .A2(new_n240), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT75), .B1(new_n242), .B2(new_n238), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n228), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n223), .A2(new_n227), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n232), .A2(KEYINPUT4), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n338), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n342), .B1(new_n223), .B2(new_n227), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n347), .A2(KEYINPUT5), .A3(new_n233), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n337), .B1(new_n241), .B2(new_n243), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n252), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n254), .A2(new_n328), .A3(new_n334), .A4(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n331), .A2(new_n333), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n351), .B1(new_n356), .B2(new_n202), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n357), .A2(KEYINPUT81), .A3(new_n328), .A4(new_n334), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n238), .A2(new_n305), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n268), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G228gat), .A2(G233gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n259), .A2(new_n260), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n305), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n259), .A2(new_n260), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n237), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n226), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n361), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT29), .B1(new_n262), .B2(new_n263), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n226), .B1(new_n370), .B2(KEYINPUT3), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n362), .B1(new_n361), .B2(new_n371), .ZN(new_n372));
  OR3_X1    g171(.A1(new_n369), .A2(G22gat), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(G22gat), .B1(new_n369), .B2(new_n372), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G78gat), .B(G106gat), .Z(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT31), .B(G50gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n378), .B(new_n379), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n373), .A2(new_n374), .A3(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n351), .A2(KEYINPUT6), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n346), .A2(new_n252), .A3(new_n350), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n388), .B2(new_n351), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT37), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n324), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n311), .A2(new_n314), .A3(KEYINPUT37), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n326), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT38), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n324), .A2(new_n317), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n311), .A2(new_n314), .A3(KEYINPUT82), .A4(KEYINPUT37), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT38), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n318), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n399), .A2(new_n391), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT83), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n384), .B1(new_n397), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT84), .B1(new_n359), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n244), .A2(new_n228), .A3(new_n343), .A4(new_n344), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n408), .A2(new_n338), .B1(new_n348), .B2(new_n349), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT77), .B1(new_n409), .B2(new_n252), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT6), .B1(new_n409), .B2(new_n252), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n346), .A2(new_n350), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT77), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n332), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n385), .ZN(new_n416));
  INV_X1    g215(.A(new_n328), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT78), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n419));
  AOI211_X1 g218(.A(new_n419), .B(new_n328), .C1(new_n415), .C2(new_n385), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n384), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G15gat), .B(G43gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G71gat), .B(G99gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n304), .B(new_n225), .ZN(new_n425));
  NAND2_X1  g224(.A1(G227gat), .A2(G233gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n426), .B(KEYINPUT64), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(KEYINPUT32), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n425), .A2(KEYINPUT34), .A3(new_n427), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n433), .A2(KEYINPUT70), .ZN(new_n434));
  XOR2_X1   g233(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n435));
  INV_X1    g234(.A(new_n426), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n425), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT69), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n438), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(KEYINPUT70), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n434), .A2(new_n439), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n432), .A2(new_n442), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT36), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT36), .ZN(new_n447));
  INV_X1    g246(.A(new_n445), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(new_n443), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n359), .A2(new_n405), .A3(KEYINPUT84), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n407), .A2(new_n421), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  XOR2_X1   g251(.A(KEYINPUT85), .B(KEYINPUT35), .Z(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n381), .B2(new_n383), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n444), .A2(new_n417), .A3(new_n445), .A4(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n389), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n416), .A2(new_n417), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n419), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n448), .A2(new_n443), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n416), .A2(KEYINPUT78), .A3(new_n417), .ZN(new_n461));
  INV_X1    g260(.A(new_n384), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n457), .B1(new_n463), .B2(KEYINPUT35), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n452), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n467), .A2(G1gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT16), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n469), .B2(G1gat), .ZN(new_n470));
  INV_X1    g269(.A(G8gat), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(KEYINPUT86), .A3(new_n471), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n468), .A2(new_n470), .A3(new_n475), .A4(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n478));
  INV_X1    g277(.A(G29gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n481));
  AOI21_X1  g280(.A(G36gat), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G36gat), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n478), .A2(new_n483), .A3(G29gat), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT15), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n484), .ZN(new_n486));
  INV_X1    g285(.A(new_n481), .ZN(new_n487));
  NOR2_X1   g286(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT15), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G43gat), .B(G50gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n485), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  INV_X1    g293(.A(new_n492), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(KEYINPUT15), .C1(new_n482), .C2(new_n484), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n494), .B1(new_n493), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n477), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G229gat), .A2(G233gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n493), .A2(new_n496), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n474), .A3(new_n476), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT87), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n499), .A2(new_n502), .A3(new_n505), .A4(new_n500), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n499), .A2(new_n502), .A3(KEYINPUT18), .A4(new_n500), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n500), .B(KEYINPUT13), .Z(new_n510));
  INV_X1    g309(.A(new_n502), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n501), .B1(new_n474), .B2(new_n476), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G113gat), .B(G141gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G197gat), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT11), .B(G169gat), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT12), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n508), .A2(new_n520), .A3(new_n514), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g323(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(G85gat), .A3(G92gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT93), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G85gat), .A2(G92gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g330(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n532));
  INV_X1    g331(.A(new_n530), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n526), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G99gat), .B(G106gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(G85gat), .A2(G92gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(KEYINPUT8), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n536), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n525), .B1(new_n543), .B2(new_n501), .ZN(new_n544));
  OAI22_X1  g343(.A1(new_n497), .A2(new_n498), .B1(new_n541), .B2(new_n542), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G190gat), .B(G218gat), .Z(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n546), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n549), .A2(new_n552), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n556));
  INV_X1    g355(.A(G64gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G57gat), .ZN(new_n558));
  INV_X1    g357(.A(G57gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(G64gat), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n556), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G71gat), .B(G78gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n566), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT90), .B(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G127gat), .B(G155gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G183gat), .B(G211gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT21), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n477), .B1(new_n579), .B2(new_n569), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n582), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n555), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n569), .B1(new_n541), .B2(new_n542), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n535), .A2(new_n531), .ZN(new_n587));
  AND2_X1   g386(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(new_n530), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n534), .B1(new_n589), .B2(new_n532), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n540), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n537), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n566), .A2(new_n568), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n567), .B1(new_n561), .B2(new_n565), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n586), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n543), .A2(KEYINPUT10), .A3(new_n596), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n603), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n600), .B2(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT94), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n586), .A2(new_n598), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n607), .ZN(new_n611));
  XNOR2_X1  g410(.A(G120gat), .B(G148gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n606), .A2(new_n609), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT95), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT94), .B1(new_n602), .B2(new_n603), .ZN(new_n619));
  AOI211_X1 g418(.A(new_n605), .B(new_n607), .C1(new_n600), .C2(new_n601), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n622), .A3(new_n616), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n614), .ZN(new_n625));
  INV_X1    g424(.A(new_n611), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n625), .B1(new_n608), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n466), .A2(new_n524), .A3(new_n585), .A4(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n415), .A2(KEYINPUT96), .A3(new_n385), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT96), .B1(new_n415), .B2(new_n385), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT97), .B(G1gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(G1324gat));
  NOR2_X1   g436(.A1(new_n630), .A2(new_n417), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n471), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT16), .B(G8gat), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n630), .A2(new_n417), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT42), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(KEYINPUT42), .B2(new_n641), .ZN(G1325gat));
  OAI21_X1  g442(.A(G15gat), .B1(new_n630), .B2(new_n450), .ZN(new_n644));
  INV_X1    g443(.A(new_n460), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n645), .A2(G15gat), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n630), .B2(new_n646), .ZN(G1326gat));
  NOR2_X1   g446(.A1(new_n630), .A2(new_n462), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT43), .B(G22gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(G1327gat));
  NAND2_X1  g449(.A1(new_n583), .A2(new_n584), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n628), .ZN(new_n652));
  AND4_X1   g451(.A1(new_n524), .A2(new_n466), .A3(new_n555), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(new_n479), .A3(new_n633), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(KEYINPUT98), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(KEYINPUT98), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT45), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n359), .A2(new_n405), .A3(KEYINPUT84), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n406), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n421), .A2(new_n450), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n464), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n555), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n660), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n466), .A2(KEYINPUT44), .A3(new_n555), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n524), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n651), .A2(new_n670), .A3(new_n628), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(G29gat), .B1(new_n672), .B2(new_n634), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n655), .A2(KEYINPUT45), .A3(new_n656), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n673), .A3(new_n674), .ZN(G1328gat));
  AOI21_X1  g474(.A(G36gat), .B1(KEYINPUT99), .B2(KEYINPUT46), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n653), .A2(new_n328), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(KEYINPUT99), .A2(KEYINPUT46), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G36gat), .B1(new_n672), .B2(new_n417), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(G1329gat));
  INV_X1    g480(.A(G43gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n450), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n667), .A2(new_n668), .A3(new_n683), .A4(new_n671), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n685), .B2(new_n684), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n653), .A2(new_n682), .A3(new_n460), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(KEYINPUT47), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(G43gat), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n690), .A2(new_n688), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(KEYINPUT47), .B2(new_n691), .ZN(G1330gat));
  NOR2_X1   g491(.A1(new_n462), .A2(G50gat), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT103), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n653), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n667), .A2(new_n668), .A3(new_n384), .A4(new_n671), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT104), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G50gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n696), .A2(KEYINPUT104), .ZN(new_n699));
  OAI211_X1 g498(.A(KEYINPUT48), .B(new_n695), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n696), .A2(new_n701), .A3(G50gat), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n696), .B2(G50gat), .ZN(new_n703));
  INV_X1    g502(.A(new_n695), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT101), .B(KEYINPUT48), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n700), .B1(new_n705), .B2(new_n706), .ZN(G1331gat));
  AND3_X1   g506(.A1(new_n585), .A2(new_n670), .A3(new_n628), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n466), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n634), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n559), .ZN(G1332gat));
  NOR2_X1   g510(.A1(new_n709), .A2(new_n417), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  AND2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n712), .B2(new_n713), .ZN(G1333gat));
  XNOR2_X1  g515(.A(new_n460), .B(KEYINPUT105), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n563), .B1(new_n709), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n466), .A2(G71gat), .A3(new_n683), .A4(new_n708), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g520(.A1(new_n709), .A2(new_n462), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(new_n564), .ZN(G1335gat));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n663), .A2(new_n661), .A3(new_n406), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT107), .B(new_n555), .C1(new_n725), .C2(new_n464), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n651), .A2(new_n524), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT106), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT107), .B1(new_n466), .B2(new_n555), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n724), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n665), .B2(new_n666), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n728), .A4(new_n726), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n734), .A3(KEYINPUT108), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n736), .B(new_n724), .C1(new_n729), .C2(new_n730), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT109), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n735), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n634), .A2(G85gat), .A3(new_n629), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n728), .A2(new_n628), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n669), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n634), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1336gat));
  NAND4_X1  g546(.A1(new_n667), .A2(new_n668), .A3(new_n328), .A4(new_n744), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(G92gat), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(KEYINPUT52), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n629), .A2(G92gat), .A3(new_n417), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n738), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n731), .B2(new_n734), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT52), .B1(new_n753), .B2(new_n749), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1337gat));
  NOR3_X1   g554(.A1(new_n645), .A2(G99gat), .A3(new_n629), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n741), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G99gat), .B1(new_n745), .B2(new_n450), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1338gat));
  NAND4_X1  g558(.A1(new_n667), .A2(new_n668), .A3(new_n384), .A4(new_n744), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT110), .B(G106gat), .Z(new_n761));
  AND2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(KEYINPUT53), .ZN(new_n763));
  OR3_X1    g562(.A1(new_n462), .A2(new_n629), .A3(G106gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n738), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n731), .B2(new_n734), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT53), .B1(new_n766), .B2(new_n762), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1339gat));
  INV_X1    g567(.A(new_n651), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n600), .A2(new_n607), .A3(new_n601), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(KEYINPUT54), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n606), .A2(new_n771), .A3(new_n609), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n614), .B1(new_n608), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(KEYINPUT55), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n622), .B1(new_n621), .B2(new_n616), .ZN(new_n776));
  NOR4_X1   g575(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT95), .A4(new_n615), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n625), .B1(new_n604), .B2(KEYINPUT54), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n621), .B2(new_n771), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(KEYINPUT55), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT111), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n772), .A2(new_n774), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n624), .A2(new_n785), .A3(new_n786), .A4(new_n775), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n782), .A2(new_n524), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n500), .B1(new_n499), .B2(new_n502), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n511), .A2(new_n512), .A3(new_n510), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n519), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n523), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n628), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n555), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n666), .A2(new_n792), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n796), .A2(new_n782), .A3(new_n787), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n769), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n585), .A2(new_n670), .A3(new_n629), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n384), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n634), .A2(new_n328), .A3(new_n645), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n524), .A3(new_n221), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n800), .B(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(new_n801), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n524), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n804), .B1(new_n809), .B2(new_n214), .ZN(G1340gat));
  NAND3_X1  g609(.A1(new_n803), .A2(new_n215), .A3(new_n628), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n807), .A2(new_n628), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(G120gat), .ZN(new_n814));
  AOI211_X1 g613(.A(KEYINPUT113), .B(new_n215), .C1(new_n807), .C2(new_n628), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(G1341gat));
  INV_X1    g615(.A(G127gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n803), .A2(new_n817), .A3(new_n651), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n807), .A2(new_n651), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n817), .ZN(G1342gat));
  NAND2_X1  g620(.A1(new_n807), .A2(new_n555), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G134gat), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n802), .A2(G134gat), .A3(new_n666), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT56), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1343gat));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n798), .A2(new_n799), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n384), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n799), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n792), .B1(new_n624), .B2(new_n627), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n524), .A2(new_n624), .A3(new_n775), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n783), .B2(new_n784), .ZN(new_n836));
  AOI211_X1 g635(.A(KEYINPUT115), .B(KEYINPUT55), .C1(new_n772), .C2(new_n774), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT116), .B1(new_n839), .B2(new_n555), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n796), .A2(new_n782), .A3(new_n787), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n524), .A2(new_n624), .A3(new_n775), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT115), .B1(new_n780), .B2(KEYINPUT55), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n783), .A2(new_n835), .A3(new_n784), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n794), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n666), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n840), .A2(new_n841), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n832), .B1(new_n849), .B2(new_n769), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n462), .A2(new_n830), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n846), .A2(new_n666), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n797), .B1(new_n855), .B2(KEYINPUT116), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n651), .B1(new_n856), .B2(new_n848), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n854), .B(new_n851), .C1(new_n857), .C2(new_n832), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n831), .A2(new_n853), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n450), .A2(new_n417), .A3(new_n633), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT114), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n524), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n827), .B1(new_n862), .B2(G141gat), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n829), .A2(G141gat), .A3(new_n670), .A4(new_n860), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n862), .B2(G141gat), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n863), .A2(new_n865), .A3(KEYINPUT58), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  AOI221_X4 g666(.A(new_n864), .B1(new_n827), .B2(new_n867), .C1(new_n862), .C2(G141gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n868), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n829), .A2(new_n860), .ZN(new_n870));
  INV_X1    g669(.A(G148gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n628), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n859), .A2(new_n861), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n629), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(KEYINPUT59), .A3(new_n871), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n829), .A2(KEYINPUT57), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n796), .A2(new_n624), .A3(new_n775), .A4(new_n785), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n651), .B1(new_n855), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n830), .B(new_n384), .C1(new_n879), .C2(new_n832), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n877), .A2(new_n628), .A3(new_n861), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n872), .B1(new_n875), .B2(new_n882), .ZN(G1345gat));
  OAI21_X1  g682(.A(G155gat), .B1(new_n873), .B2(new_n769), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n870), .A2(new_n204), .A3(new_n651), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1346gat));
  OAI21_X1  g685(.A(G162gat), .B1(new_n873), .B2(new_n666), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n205), .A3(new_n555), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1347gat));
  NOR3_X1   g688(.A1(new_n645), .A2(new_n417), .A3(new_n384), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n828), .A2(new_n634), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT119), .ZN(new_n892));
  AOI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n524), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n717), .A2(new_n417), .A3(new_n633), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n806), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n524), .A2(G169gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(G1348gat));
  AOI21_X1  g696(.A(G176gat), .B1(new_n892), .B2(new_n628), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT120), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(G176gat), .A3(new_n628), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(G1349gat));
  AND2_X1   g701(.A1(new_n800), .A2(new_n805), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n800), .A2(new_n805), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n651), .B(new_n894), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT122), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n806), .A2(new_n907), .A3(new_n651), .A4(new_n894), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n908), .A3(G183gat), .ZN(new_n909));
  INV_X1    g708(.A(new_n272), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n891), .A2(new_n910), .A3(new_n769), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT60), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n909), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n892), .A2(new_n273), .A3(new_n555), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n895), .A2(new_n555), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(G190gat), .ZN(new_n921));
  AOI211_X1 g720(.A(KEYINPUT61), .B(new_n273), .C1(new_n895), .C2(new_n555), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(G1351gat));
  NAND3_X1  g722(.A1(new_n877), .A2(KEYINPUT123), .A3(new_n880), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n683), .A2(new_n633), .A3(new_n417), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n462), .B1(new_n798), .B2(new_n799), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n880), .B1(new_n926), .B2(new_n830), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n924), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n670), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n926), .A2(new_n925), .ZN(new_n932));
  INV_X1    g731(.A(G197gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n933), .A3(new_n524), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT124), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1352gat));
  OAI21_X1  g738(.A(G204gat), .B1(new_n930), .B2(new_n629), .ZN(new_n940));
  AOI21_X1  g739(.A(G204gat), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n932), .A2(new_n628), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n940), .A2(new_n944), .ZN(G1353gat));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n651), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n829), .A2(G211gat), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n927), .A2(new_n946), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT126), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n953), .B(new_n947), .C1(new_n949), .C2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1354gat));
  INV_X1    g754(.A(G218gat), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n930), .A2(new_n956), .A3(new_n666), .ZN(new_n957));
  AOI21_X1  g756(.A(G218gat), .B1(new_n932), .B2(new_n555), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


