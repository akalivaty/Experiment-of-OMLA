

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  NOR2_X2 U323 ( .A1(n542), .A2(n418), .ZN(n567) );
  XNOR2_X1 U324 ( .A(G36GAT), .B(G190GAT), .ZN(n315) );
  XNOR2_X1 U325 ( .A(n415), .B(KEYINPUT54), .ZN(n416) );
  XNOR2_X1 U326 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U327 ( .A(n435), .B(KEYINPUT55), .ZN(n452) );
  XNOR2_X1 U328 ( .A(n453), .B(KEYINPUT121), .ZN(n564) );
  XNOR2_X1 U329 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U330 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT97), .B(KEYINPUT4), .Z(n292) );
  XNOR2_X1 U332 ( .A(KEYINPUT95), .B(G57GAT), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U334 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n294) );
  XNOR2_X1 U335 ( .A(KEYINPUT5), .B(KEYINPUT94), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U337 ( .A(n296), .B(n295), .Z(n306) );
  XNOR2_X1 U338 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n297) );
  XNOR2_X1 U339 ( .A(n297), .B(G155GAT), .ZN(n298) );
  XOR2_X1 U340 ( .A(n298), .B(KEYINPUT2), .Z(n300) );
  XNOR2_X1 U341 ( .A(KEYINPUT91), .B(KEYINPUT3), .ZN(n299) );
  XNOR2_X1 U342 ( .A(n300), .B(n299), .ZN(n432) );
  XNOR2_X1 U343 ( .A(G134GAT), .B(G127GAT), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n301), .B(KEYINPUT0), .ZN(n442) );
  XOR2_X1 U345 ( .A(G113GAT), .B(G1GAT), .Z(n360) );
  XOR2_X1 U346 ( .A(n442), .B(n360), .Z(n303) );
  NAND2_X1 U347 ( .A1(G225GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n432), .B(n304), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n314) );
  XOR2_X1 U351 ( .A(KEYINPUT96), .B(KEYINPUT1), .Z(n308) );
  XNOR2_X1 U352 ( .A(G120GAT), .B(G148GAT), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U354 ( .A(G85GAT), .B(G162GAT), .Z(n310) );
  XNOR2_X1 U355 ( .A(G29GAT), .B(G141GAT), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U357 ( .A(n312), .B(n311), .Z(n313) );
  XNOR2_X1 U358 ( .A(n314), .B(n313), .ZN(n542) );
  XOR2_X1 U359 ( .A(G169GAT), .B(G8GAT), .Z(n359) );
  XNOR2_X1 U360 ( .A(n315), .B(KEYINPUT76), .ZN(n386) );
  XNOR2_X1 U361 ( .A(n386), .B(KEYINPUT98), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n316), .B(KEYINPUT78), .ZN(n317) );
  XOR2_X1 U363 ( .A(n359), .B(n317), .Z(n319) );
  NAND2_X1 U364 ( .A1(G226GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n322) );
  XOR2_X1 U366 ( .A(G64GAT), .B(G92GAT), .Z(n321) );
  XNOR2_X1 U367 ( .A(G176GAT), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n321), .B(n320), .ZN(n375) );
  XOR2_X1 U369 ( .A(n322), .B(n375), .Z(n330) );
  XOR2_X1 U370 ( .A(G183GAT), .B(KEYINPUT17), .Z(n324) );
  XNOR2_X1 U371 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n447) );
  XNOR2_X1 U373 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n325), .B(KEYINPUT21), .ZN(n326) );
  XOR2_X1 U375 ( .A(n326), .B(KEYINPUT88), .Z(n328) );
  XNOR2_X1 U376 ( .A(G197GAT), .B(G218GAT), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n431) );
  XNOR2_X1 U378 ( .A(n447), .B(n431), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n462) );
  XOR2_X1 U380 ( .A(G127GAT), .B(G71GAT), .Z(n332) );
  XNOR2_X1 U381 ( .A(G15GAT), .B(G183GAT), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U383 ( .A(KEYINPUT78), .B(G64GAT), .Z(n334) );
  XNOR2_X1 U384 ( .A(G1GAT), .B(G8GAT), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U386 ( .A(n336), .B(n335), .Z(n341) );
  XOR2_X1 U387 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n338) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U390 ( .A(KEYINPUT15), .B(n339), .ZN(n340) );
  XOR2_X1 U391 ( .A(n341), .B(n340), .Z(n346) );
  XNOR2_X1 U392 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n342), .B(KEYINPUT13), .ZN(n372) );
  XOR2_X1 U394 ( .A(n372), .B(G211GAT), .Z(n344) );
  XNOR2_X1 U395 ( .A(G22GAT), .B(G78GAT), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n351) );
  XOR2_X1 U398 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n348) );
  XNOR2_X1 U399 ( .A(KEYINPUT12), .B(KEYINPUT80), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U401 ( .A(G155GAT), .B(n349), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n563) );
  XNOR2_X1 U403 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n352), .B(G29GAT), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n353), .B(KEYINPUT7), .ZN(n355) );
  XOR2_X1 U406 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n390) );
  XOR2_X1 U408 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n357) );
  XNOR2_X1 U409 ( .A(G197GAT), .B(G15GAT), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n390), .B(n358), .ZN(n370) );
  XOR2_X1 U412 ( .A(G50GAT), .B(G36GAT), .Z(n362) );
  XNOR2_X1 U413 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U415 ( .A(G141GAT), .B(G22GAT), .Z(n419) );
  XOR2_X1 U416 ( .A(n363), .B(n419), .Z(n368) );
  XOR2_X1 U417 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n365) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U420 ( .A(KEYINPUT30), .B(n366), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U422 ( .A(n370), .B(n369), .ZN(n555) );
  XNOR2_X1 U423 ( .A(G99GAT), .B(G85GAT), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n371), .B(KEYINPUT73), .ZN(n398) );
  XOR2_X1 U425 ( .A(n372), .B(n398), .Z(n377) );
  XOR2_X1 U426 ( .A(G78GAT), .B(G148GAT), .Z(n374) );
  XNOR2_X1 U427 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n420) );
  XNOR2_X1 U429 ( .A(n420), .B(n375), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n384) );
  XOR2_X1 U431 ( .A(G120GAT), .B(G71GAT), .Z(n443) );
  XOR2_X1 U432 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n379) );
  XNOR2_X1 U433 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U435 ( .A(n443), .B(n380), .Z(n382) );
  NAND2_X1 U436 ( .A1(G230GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U438 ( .A(n384), .B(n383), .Z(n574) );
  XNOR2_X1 U439 ( .A(KEYINPUT41), .B(n574), .ZN(n558) );
  NAND2_X1 U440 ( .A1(n555), .A2(n558), .ZN(n385) );
  XNOR2_X1 U441 ( .A(KEYINPUT46), .B(n385), .ZN(n403) );
  XOR2_X1 U442 ( .A(n386), .B(G92GAT), .Z(n388) );
  NAND2_X1 U443 ( .A1(G232GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n402) );
  XOR2_X1 U446 ( .A(KEYINPUT9), .B(G218GAT), .Z(n392) );
  XNOR2_X1 U447 ( .A(G134GAT), .B(G106GAT), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U449 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n394) );
  XNOR2_X1 U450 ( .A(KEYINPUT10), .B(KEYINPUT77), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U452 ( .A(n396), .B(n395), .Z(n400) );
  XNOR2_X1 U453 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n397), .B(G162GAT), .ZN(n424) );
  XNOR2_X1 U455 ( .A(n424), .B(n398), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n484) );
  NAND2_X1 U458 ( .A1(n403), .A2(n484), .ZN(n404) );
  NOR2_X1 U459 ( .A1(n563), .A2(n404), .ZN(n405) );
  XOR2_X1 U460 ( .A(KEYINPUT47), .B(n405), .Z(n413) );
  INV_X1 U461 ( .A(n574), .ZN(n408) );
  INV_X1 U462 ( .A(n563), .ZN(n577) );
  XNOR2_X1 U463 ( .A(n484), .B(KEYINPUT36), .ZN(n580) );
  NOR2_X1 U464 ( .A1(n577), .A2(n580), .ZN(n406) );
  XOR2_X1 U465 ( .A(KEYINPUT45), .B(n406), .Z(n407) );
  NOR2_X1 U466 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n409), .B(KEYINPUT113), .ZN(n410) );
  NOR2_X1 U468 ( .A1(n410), .A2(n555), .ZN(n411) );
  XNOR2_X1 U469 ( .A(KEYINPUT114), .B(n411), .ZN(n412) );
  NOR2_X1 U470 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U471 ( .A(KEYINPUT48), .B(n414), .ZN(n540) );
  NOR2_X1 U472 ( .A1(n462), .A2(n540), .ZN(n417) );
  INV_X1 U473 ( .A(KEYINPUT120), .ZN(n415) );
  XOR2_X1 U474 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U477 ( .A(n423), .B(G204GAT), .Z(n426) );
  XNOR2_X1 U478 ( .A(n424), .B(KEYINPUT92), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U480 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n428) );
  XNOR2_X1 U481 ( .A(KEYINPUT23), .B(KEYINPUT86), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U483 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n470) );
  NAND2_X1 U486 ( .A1(n567), .A2(n470), .ZN(n435) );
  XOR2_X1 U487 ( .A(G99GAT), .B(G190GAT), .Z(n437) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(G113GAT), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U490 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n439) );
  XNOR2_X1 U491 ( .A(G15GAT), .B(KEYINPUT84), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n451) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U497 ( .A(n446), .B(G176GAT), .Z(n449) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U500 ( .A(n451), .B(n450), .ZN(n528) );
  NAND2_X1 U501 ( .A1(n452), .A2(n528), .ZN(n453) );
  INV_X1 U502 ( .A(n484), .ZN(n552) );
  NAND2_X1 U503 ( .A1(n564), .A2(n552), .ZN(n457) );
  XOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n455) );
  INV_X1 U505 ( .A(G190GAT), .ZN(n454) );
  INV_X1 U506 ( .A(G43GAT), .ZN(n483) );
  XNOR2_X1 U507 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n481) );
  NAND2_X1 U508 ( .A1(n555), .A2(n574), .ZN(n489) );
  XNOR2_X1 U509 ( .A(KEYINPUT25), .B(KEYINPUT102), .ZN(n461) );
  INV_X1 U510 ( .A(n462), .ZN(n519) );
  NAND2_X1 U511 ( .A1(n519), .A2(n528), .ZN(n458) );
  NAND2_X1 U512 ( .A1(n458), .A2(n470), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT103), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n461), .B(n460), .ZN(n467) );
  XNOR2_X1 U515 ( .A(n462), .B(KEYINPUT99), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(KEYINPUT27), .ZN(n472) );
  INV_X1 U517 ( .A(KEYINPUT26), .ZN(n466) );
  NOR2_X1 U518 ( .A1(n528), .A2(n470), .ZN(n464) );
  XNOR2_X1 U519 ( .A(KEYINPUT101), .B(n464), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n466), .B(n465), .ZN(n566) );
  NAND2_X1 U521 ( .A1(n472), .A2(n566), .ZN(n539) );
  NAND2_X1 U522 ( .A1(n467), .A2(n539), .ZN(n468) );
  XOR2_X1 U523 ( .A(KEYINPUT104), .B(n468), .Z(n469) );
  NOR2_X1 U524 ( .A1(n542), .A2(n469), .ZN(n476) );
  XOR2_X1 U525 ( .A(n470), .B(KEYINPUT64), .Z(n471) );
  XNOR2_X1 U526 ( .A(KEYINPUT28), .B(n471), .ZN(n524) );
  NAND2_X1 U527 ( .A1(n472), .A2(n542), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n524), .A2(n473), .ZN(n527) );
  XOR2_X1 U529 ( .A(n527), .B(KEYINPUT100), .Z(n474) );
  NOR2_X1 U530 ( .A1(n528), .A2(n474), .ZN(n475) );
  NOR2_X1 U531 ( .A1(n476), .A2(n475), .ZN(n488) );
  NOR2_X1 U532 ( .A1(n488), .A2(n580), .ZN(n477) );
  NAND2_X1 U533 ( .A1(n577), .A2(n477), .ZN(n478) );
  XOR2_X1 U534 ( .A(KEYINPUT37), .B(n478), .Z(n517) );
  NOR2_X1 U535 ( .A1(n489), .A2(n517), .ZN(n479) );
  XNOR2_X1 U536 ( .A(n479), .B(KEYINPUT38), .ZN(n503) );
  AND2_X1 U537 ( .A1(n528), .A2(n503), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n483), .B(n482), .ZN(G1330GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT83), .B(KEYINPUT16), .Z(n486) );
  NAND2_X1 U541 ( .A1(n563), .A2(n484), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n486), .B(n485), .ZN(n487) );
  OR2_X1 U543 ( .A1(n488), .A2(n487), .ZN(n505) );
  NOR2_X1 U544 ( .A1(n489), .A2(n505), .ZN(n497) );
  NAND2_X1 U545 ( .A1(n542), .A2(n497), .ZN(n493) );
  XOR2_X1 U546 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n491) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U549 ( .A(n493), .B(n492), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n519), .A2(n497), .ZN(n494) );
  XNOR2_X1 U551 ( .A(n494), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U553 ( .A1(n497), .A2(n528), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NAND2_X1 U555 ( .A1(n524), .A2(n497), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n498), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U557 ( .A1(n503), .A2(n542), .ZN(n501) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n499), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n503), .A2(n519), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n503), .A2(n524), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n508) );
  INV_X1 U566 ( .A(n555), .ZN(n568) );
  NAND2_X1 U567 ( .A1(n568), .A2(n558), .ZN(n516) );
  OR2_X1 U568 ( .A1(n505), .A2(n516), .ZN(n506) );
  XOR2_X1 U569 ( .A(KEYINPUT110), .B(n506), .Z(n513) );
  NAND2_X1 U570 ( .A1(n513), .A2(n542), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n509), .ZN(G1332GAT) );
  XOR2_X1 U573 ( .A(G64GAT), .B(KEYINPUT111), .Z(n511) );
  NAND2_X1 U574 ( .A1(n513), .A2(n519), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n528), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U579 ( .A1(n513), .A2(n524), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n523), .A2(n542), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n519), .A2(n523), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n523), .A2(n528), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(KEYINPUT112), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT115), .Z(n531) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n540), .A2(n529), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n536), .A2(n555), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U598 ( .A1(n536), .A2(n558), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NAND2_X1 U600 ( .A1(n536), .A2(n563), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U604 ( .A1(n536), .A2(n552), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT116), .B(n543), .Z(n553) );
  NAND2_X1 U609 ( .A1(n553), .A2(n555), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n546) );
  NAND2_X1 U612 ( .A1(n553), .A2(n558), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT117), .Z(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U617 ( .A1(n563), .A2(n553), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n557) );
  NAND2_X1 U623 ( .A1(n555), .A2(n564), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n560) );
  NAND2_X1 U626 ( .A1(n564), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT56), .Z(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n579) );
  NOR2_X1 U633 ( .A1(n568), .A2(n579), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT59), .B(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n579), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

