//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n629, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n462), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n465), .A2(KEYINPUT67), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n477), .B2(G2105), .ZN(G160));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n472), .A2(new_n462), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n472), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n484), .A2(new_n485), .A3(G136), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n484), .B2(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n470), .B2(new_n471), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(new_n493), .C1(new_n470), .C2(new_n471), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n462), .C1(new_n470), .C2(new_n471), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n465), .A2(new_n501), .A3(G138), .A4(new_n462), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n510), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n515), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n514), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n521), .B(KEYINPUT70), .C1(new_n514), .C2(new_n522), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n509), .A2(G51), .B1(new_n512), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n525), .A2(KEYINPUT71), .A3(new_n526), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(new_n509), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n514), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  AND2_X1   g115(.A1(KEYINPUT5), .A2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(KEYINPUT5), .A2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n517), .B1(new_n545), .B2(KEYINPUT72), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(KEYINPUT72), .B2(new_n545), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n512), .A2(new_n513), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G81), .B1(G43), .B2(new_n509), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n513), .A2(G53), .A3(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n509), .A2(KEYINPUT74), .A3(new_n559), .A4(G53), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n557), .B2(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n562), .A3(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n561), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n548), .A2(KEYINPUT75), .A3(G91), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n514), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n543), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n567), .A2(new_n570), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n566), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n509), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n514), .ZN(G288));
  OAI21_X1  g157(.A(G61), .B1(new_n541), .B2(new_n542), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(KEYINPUT76), .A3(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n548), .A2(G86), .B1(G48), .B2(new_n509), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT76), .B1(new_n585), .B2(G651), .ZN(new_n594));
  AOI211_X1 g169(.A(new_n587), .B(new_n517), .C1(new_n583), .C2(new_n584), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT77), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n517), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n509), .A2(G47), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n512), .A2(new_n513), .A3(G85), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n602), .A2(KEYINPUT78), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT78), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(KEYINPUT79), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n608), .B(new_n601), .C1(new_n604), .C2(new_n605), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n609), .ZN(G290));
  NAND3_X1  g185(.A1(new_n548), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n514), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G79), .ZN(new_n616));
  OR3_X1    g191(.A1(new_n616), .A2(new_n506), .A3(KEYINPUT80), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT80), .B1(new_n616), .B2(new_n506), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n543), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(G171), .ZN(G284));
  OAI21_X1  g200(.A(new_n624), .B1(new_n623), .B2(G171), .ZN(G321));
  AND3_X1   g201(.A1(G286), .A2(KEYINPUT81), .A3(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  AOI21_X1  g203(.A(KEYINPUT81), .B1(G299), .B2(new_n623), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(G297));
  AOI21_X1  g205(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(G280));
  AND2_X1   g206(.A1(new_n615), .A2(new_n621), .ZN(new_n632));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n547), .A2(new_n549), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(new_n623), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n622), .A2(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(new_n623), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n484), .A2(G135), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n462), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n482), .A2(new_n643), .A3(G123), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n482), .B2(G123), .ZN(new_n645));
  OAI221_X1 g220(.A(new_n640), .B1(new_n641), .B2(new_n642), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT84), .B(G2096), .Z(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n465), .A2(new_n463), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT13), .B(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n648), .A2(new_n649), .A3(new_n654), .ZN(G156));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(G401));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2096), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n684), .B2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  NOR2_X1   g274(.A1(G16), .A2(G21), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G168), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1966), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n550), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G16), .B2(G19), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT88), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT88), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G1341), .ZN(new_n708));
  INV_X1    g283(.A(G1341), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n705), .A2(new_n709), .A3(new_n706), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n702), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NOR2_X1   g287(.A1(G171), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G5), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G1961), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT31), .B(G11), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT94), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G28), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n720), .B2(G28), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n719), .B1(new_n721), .B2(new_n723), .C1(new_n646), .C2(new_n722), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n716), .A2(new_n717), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(G162), .A2(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G29), .B2(G35), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT29), .B(G2090), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(G164), .A2(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G27), .B2(G29), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n727), .A2(new_n729), .B1(new_n733), .B2(new_n732), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n722), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT25), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n484), .A2(KEYINPUT90), .A3(G139), .ZN(new_n742));
  AOI21_X1  g317(.A(KEYINPUT90), .B1(new_n484), .B2(G139), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n740), .B1(new_n462), .B2(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2072), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n725), .A2(new_n735), .A3(new_n736), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n722), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT28), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n484), .A2(G140), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n482), .A2(G128), .ZN(new_n751));
  OR2_X1    g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G29), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(KEYINPUT89), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(KEYINPUT89), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n749), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G34), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n763), .A2(KEYINPUT92), .B1(G34), .B2(new_n761), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT92), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(G160), .A2(G29), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2084), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n760), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n747), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n712), .A2(G20), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT23), .Z(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G299), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n722), .A2(G32), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n463), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n482), .A2(G129), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT93), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n775), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G4), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n632), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n785), .A2(new_n786), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n787), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n711), .A2(new_n770), .A3(new_n774), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n712), .A2(G22), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT85), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n712), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1971), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n712), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G288), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n803), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n805), .A2(G1976), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(G1976), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n799), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT34), .ZN(new_n810));
  NOR2_X1   g385(.A1(G6), .A2(G16), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n598), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT32), .B(G1981), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n814), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n809), .B(new_n810), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n722), .A2(G25), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n484), .A2(G131), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n482), .A2(G119), .ZN(new_n820));
  OR2_X1    g395(.A1(G95), .A2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n821), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n818), .B1(new_n824), .B2(new_n722), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G1991), .Z(new_n826));
  XOR2_X1   g401(.A(new_n825), .B(new_n826), .Z(new_n827));
  AOI21_X1  g402(.A(new_n712), .B1(new_n607), .B2(new_n609), .ZN(new_n828));
  INV_X1    g403(.A(G1986), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n712), .A2(G24), .ZN(new_n830));
  OR3_X1    g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n817), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT86), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT86), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n817), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n809), .B1(new_n816), .B2(new_n815), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT87), .B(KEYINPUT36), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n795), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT36), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(KEYINPUT87), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n835), .A2(new_n844), .A3(new_n837), .A4(new_n839), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(G311));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n842), .A2(new_n847), .A3(new_n845), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n847), .B1(new_n842), .B2(new_n845), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(G150));
  NAND2_X1  g425(.A1(new_n509), .A2(G55), .ZN(new_n851));
  INV_X1    g426(.A(G93), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(new_n514), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n517), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G860), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n632), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  INV_X1    g436(.A(new_n856), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n547), .A2(new_n856), .A3(new_n549), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n861), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT96), .Z(new_n869));
  OAI21_X1  g444(.A(new_n857), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n859), .B1(new_n869), .B2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(new_n784), .B(new_n754), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n652), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n744), .B(new_n504), .ZN(new_n874));
  AOI22_X1  g449(.A1(G130), .A2(new_n482), .B1(new_n484), .B2(G142), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  INV_X1    g451(.A(G118), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n876), .A2(KEYINPUT97), .B1(new_n877), .B2(G2105), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(KEYINPUT97), .B2(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n824), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n874), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n873), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n873), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n646), .B(G160), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G162), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  INV_X1    g465(.A(new_n888), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n885), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(KEYINPUT98), .B(KEYINPUT40), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(G395));
  NAND2_X1  g470(.A1(new_n598), .A2(G303), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n593), .A2(new_n597), .A3(G166), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT101), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NOR2_X1   g476(.A1(G290), .A2(G288), .ZN(new_n902));
  INV_X1    g477(.A(G288), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n607), .B2(new_n609), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n898), .B(KEYINPUT101), .C1(new_n902), .C2(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n566), .A2(new_n622), .A3(new_n574), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT100), .ZN(new_n911));
  NAND2_X1  g486(.A1(G299), .A2(new_n632), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n566), .A2(new_n622), .A3(new_n913), .A4(new_n574), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n622), .B1(new_n566), .B2(new_n574), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(new_n916), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n915), .A2(new_n916), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n865), .A2(KEYINPUT99), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n863), .A2(new_n921), .A3(new_n864), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n920), .A2(new_n922), .A3(new_n637), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n637), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n922), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n632), .A2(new_n633), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n912), .A2(new_n910), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n920), .A2(new_n922), .A3(new_n637), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n925), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n925), .B2(new_n932), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n909), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n925), .A2(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT42), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n925), .A2(new_n932), .A3(new_n933), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n908), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G868), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n856), .A2(G868), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(G295));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n942), .B2(new_n944), .ZN(new_n947));
  AOI211_X1 g522(.A(KEYINPUT102), .B(new_n943), .C1(new_n941), .C2(G868), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(G331));
  XNOR2_X1  g524(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n531), .A2(new_n532), .A3(G301), .ZN(new_n952));
  AOI21_X1  g527(.A(G301), .B1(new_n531), .B2(new_n532), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n865), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(G168), .A2(G171), .ZN(new_n955));
  INV_X1    g530(.A(new_n864), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n856), .B1(new_n547), .B2(new_n549), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n531), .A2(new_n532), .A3(G301), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n954), .A2(new_n960), .A3(new_n929), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n954), .A2(new_n960), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n919), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n890), .B1(new_n963), .B2(new_n908), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n915), .A2(new_n916), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n918), .A2(new_n910), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n954), .A2(new_n960), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n969), .A2(new_n961), .B1(new_n906), .B2(new_n907), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n951), .B1(new_n964), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n910), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n916), .B1(new_n972), .B2(new_n917), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n918), .A2(new_n911), .A3(new_n976), .A4(new_n914), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n929), .A2(KEYINPUT104), .A3(new_n916), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n918), .A2(new_n911), .A3(new_n914), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT105), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n962), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n961), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n954), .A2(new_n960), .A3(KEYINPUT106), .A4(new_n929), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n908), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n965), .A2(new_n966), .B1(new_n954), .B2(new_n960), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n954), .A2(new_n960), .A3(new_n929), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G37), .B1(new_n909), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n971), .B1(new_n992), .B2(new_n951), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n994), .B1(new_n992), .B2(KEYINPUT43), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n964), .A2(new_n951), .A3(new_n970), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n987), .B2(new_n991), .ZN(new_n1002));
  NOR4_X1   g577(.A1(new_n1002), .A2(new_n998), .A3(KEYINPUT107), .A4(new_n994), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n995), .B1(new_n1000), .B2(new_n1003), .ZN(G397));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n498), .B2(new_n503), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n477), .A2(G2105), .ZN(new_n1009));
  INV_X1    g584(.A(new_n468), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(G40), .A3(new_n1010), .ZN(new_n1011));
  AOI211_X1 g586(.A(KEYINPUT108), .B(G1384), .C1(new_n498), .C2(new_n503), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n784), .B(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n823), .B(new_n826), .Z(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT109), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n754), .B(new_n759), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(G290), .B(G1986), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1013), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1384), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n504), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT50), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1009), .A2(G40), .A3(new_n1010), .ZN(new_n1025));
  INV_X1    g600(.A(G2084), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1006), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(G40), .B(G160), .C1(new_n1006), .C2(KEYINPUT45), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(G168), .B(new_n1029), .C1(new_n1032), .C2(G1966), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(KEYINPUT123), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(KEYINPUT51), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1029), .B1(new_n1032), .B2(G1966), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(G8), .A3(G286), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1044));
  OAI211_X1 g619(.A(G40), .B(G160), .C1(new_n1006), .C2(new_n1027), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1006), .A2(new_n1027), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1045), .A2(new_n1046), .A3(G2090), .ZN(new_n1047));
  INV_X1    g622(.A(G1971), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT45), .B1(new_n504), .B2(new_n1022), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(new_n1011), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT110), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1006), .A2(new_n1053), .A3(KEYINPUT45), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1047), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(new_n1034), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G303), .A2(G8), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT55), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G288), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT112), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1006), .A2(G160), .A3(G40), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1066), .A2(KEYINPUT111), .A3(G8), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT111), .B1(new_n1066), .B2(G8), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1064), .B(new_n1065), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n596), .A2(G1981), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT49), .ZN(new_n1072));
  INV_X1    g647(.A(G1981), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n592), .B(new_n1073), .C1(new_n594), .C2(new_n595), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1067), .A2(new_n1068), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1073), .B1(new_n590), .B2(new_n592), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1074), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT49), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1084), .B(KEYINPUT114), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1070), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1059), .B1(new_n1056), .B2(new_n1034), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT113), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1064), .B(new_n1090), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(KEYINPUT52), .A3(new_n1091), .ZN(new_n1092));
  AND4_X1   g667(.A1(new_n1061), .A2(new_n1086), .A3(new_n1087), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1055), .B2(G2078), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT119), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1024), .A2(new_n1025), .A3(new_n1097), .A4(new_n1028), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n715), .A3(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1032), .A2(new_n733), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT124), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1032), .A2(new_n1103), .A3(new_n733), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(KEYINPUT53), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(G301), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1040), .A2(new_n1107), .A3(new_n1042), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1044), .A2(new_n1093), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1110));
  AOI211_X1 g685(.A(G1976), .B(G288), .C1(new_n1079), .C2(new_n1085), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1110), .B1(new_n1111), .B2(new_n1081), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1086), .A2(new_n1060), .A3(new_n1057), .A4(new_n1092), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1096), .A2(new_n790), .A3(new_n1098), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1066), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n759), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n632), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .A4(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT116), .B(G1956), .Z(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n563), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1127), .A2(new_n564), .B1(new_n558), .B2(new_n560), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n567), .A2(new_n570), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n573), .A2(G651), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1126), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n566), .A2(new_n574), .A3(new_n1125), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1121), .A2(new_n1134), .A3(new_n1123), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT118), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1121), .A2(new_n1139), .A3(new_n1134), .A4(new_n1123), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1119), .A2(new_n1136), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1136), .A2(KEYINPUT61), .A3(new_n1137), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n632), .B2(KEYINPUT122), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n632), .A2(KEYINPUT122), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1115), .A2(new_n1117), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1115), .A2(new_n1117), .A3(new_n1144), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1145), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1142), .B(new_n1146), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT61), .B1(new_n1152), .B2(new_n1136), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1155), .A2(KEYINPUT120), .A3(new_n1014), .A4(new_n1050), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1055), .B2(G1996), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(new_n709), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1156), .B(new_n1158), .C1(new_n1116), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n550), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT59), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1164), .A3(new_n550), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1141), .B1(new_n1154), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT54), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1025), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT125), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1094), .A2(G2078), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1052), .A2(new_n1054), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1173), .B(new_n1025), .C1(new_n1008), .C2(new_n1012), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1170), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1175), .A2(new_n1095), .A3(new_n1099), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1168), .B1(new_n1176), .B2(G171), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1100), .A2(G301), .A3(new_n1105), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1177), .A2(new_n1178), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1176), .A2(G171), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1168), .B1(new_n1106), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1179), .A2(new_n1093), .A3(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1109), .B(new_n1114), .C1(new_n1167), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1041), .A2(G8), .A3(G168), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1093), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1061), .A2(KEYINPUT63), .A3(new_n1185), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1086), .A2(new_n1087), .A3(new_n1092), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT115), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1184), .A2(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1021), .B1(new_n1183), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n824), .A2(new_n826), .ZN(new_n1195));
  OAI22_X1  g770(.A1(new_n1194), .A2(new_n1195), .B1(G2067), .B2(new_n754), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1013), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1019), .A2(new_n1013), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT48), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1013), .A2(new_n829), .A3(new_n607), .A4(new_n609), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1200), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1202), .A2(KEYINPUT48), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1197), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT46), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT126), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1018), .A2(new_n783), .A3(new_n782), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1013), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT127), .Z(new_n1212));
  NAND3_X1  g787(.A1(new_n1208), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  OR2_X1    g788(.A1(new_n1213), .A2(KEYINPUT47), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(KEYINPUT47), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1204), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1193), .A2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g792(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1219));
  NAND3_X1  g793(.A1(new_n1219), .A2(new_n893), .A3(new_n993), .ZN(G225));
  INV_X1    g794(.A(G225), .ZN(G308));
endmodule


