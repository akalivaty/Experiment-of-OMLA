//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NOR4_X1   g0022(.A1(new_n215), .A2(new_n218), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G50), .ZN(new_n224));
  INV_X1    g0024(.A(G226), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n206), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(G20), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n203), .A2(G50), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n210), .B(new_n233), .C1(new_n236), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n230), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n217), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n224), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n229), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  INV_X1    g0051(.A(G107), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(new_n216), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n250), .B(new_n254), .ZN(G351));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI211_X1 g0057(.A(G232), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  OAI211_X1 g0059(.A(G226), .B(new_n259), .C1(new_n256), .C2(new_n257), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G97), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n234), .B1(G33), .B2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT66), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G41), .A2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n263), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G238), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n265), .A3(G274), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n264), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n264), .A2(new_n273), .A3(new_n278), .A4(new_n274), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(KEYINPUT68), .A3(KEYINPUT13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G190), .ZN(new_n283));
  INV_X1    g0083(.A(G200), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n276), .B2(new_n279), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G20), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n288), .A2(G77), .B1(G20), .B2(new_n219), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n289), .B1(new_n224), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n234), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT11), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n294), .B1(new_n269), .B2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G68), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  AOI211_X1 g0099(.A(new_n299), .B(new_n235), .C1(new_n266), .C2(new_n268), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n219), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n283), .A2(new_n286), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT69), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n303), .B1(new_n282), .B2(G190), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT69), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(new_n286), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n282), .A2(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n276), .A2(new_n279), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT14), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n315), .A3(G169), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n311), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n303), .ZN(new_n318));
  XOR2_X1   g0118(.A(KEYINPUT8), .B(G58), .Z(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(new_n288), .B1(G150), .B2(new_n290), .ZN(new_n320));
  OAI21_X1  g0120(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n294), .B1(new_n224), .B2(new_n300), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n297), .A2(G50), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(KEYINPUT9), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT9), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n323), .B2(new_n324), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT67), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n287), .ZN(new_n332));
  NAND2_X1  g0132(.A1(KEYINPUT3), .A2(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n259), .ZN(new_n335));
  INV_X1    g0135(.A(G222), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n330), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n334), .A2(KEYINPUT67), .A3(G222), .A4(new_n259), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n256), .A2(new_n257), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G77), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(G223), .A3(G1698), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n337), .A2(new_n338), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n263), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n272), .A2(G226), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n343), .A2(new_n274), .A3(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n345), .A2(new_n284), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n343), .A2(G190), .A3(new_n274), .A4(new_n344), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n329), .A2(new_n346), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n326), .B2(new_n328), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n345), .A2(new_n284), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT10), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G179), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n345), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n355), .B(new_n325), .C1(G169), .C2(new_n345), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n310), .A2(new_n318), .A3(new_n353), .A4(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n288), .ZN(new_n360));
  INV_X1    g0160(.A(new_n319), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n360), .B1(new_n235), .B2(new_n226), .C1(new_n291), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n294), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n297), .A2(G77), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n300), .A2(new_n226), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n334), .A2(G238), .A3(G1698), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n368), .B1(new_n252), .B2(new_n334), .C1(new_n335), .C2(new_n230), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n263), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n272), .A2(G244), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n274), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n372), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(new_n284), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n229), .A2(new_n219), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n378), .B2(new_n202), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n290), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n332), .A2(KEYINPUT7), .A3(new_n235), .A4(new_n333), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n332), .A2(new_n235), .A3(new_n333), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT70), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT70), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n384), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT16), .B(new_n382), .C1(new_n391), .C2(new_n219), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n219), .B1(new_n387), .B2(new_n383), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n381), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT71), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT71), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(new_n393), .C1(new_n394), .C2(new_n381), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n392), .A2(new_n396), .A3(new_n294), .A4(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G41), .ZN(new_n400));
  OAI211_X1 g0200(.A(G1), .B(G13), .C1(new_n287), .C2(new_n400), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT66), .B(G1), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(new_n270), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n274), .B1(new_n403), .B2(new_n230), .ZN(new_n404));
  OR2_X1    g0204(.A1(G223), .A2(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n225), .A2(G1698), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(new_n406), .C1(new_n256), .C2(new_n257), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n401), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n284), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n404), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(KEYINPUT72), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT72), .ZN(new_n413));
  AOI211_X1 g0213(.A(new_n413), .B(new_n401), .C1(new_n407), .C2(new_n408), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n411), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n410), .B1(new_n415), .B2(G190), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n361), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n297), .B2(new_n361), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n399), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n399), .A2(KEYINPUT17), .A3(new_n416), .A4(new_n419), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  INV_X1    g0226(.A(new_n419), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n396), .A2(new_n398), .ZN(new_n428));
  INV_X1    g0228(.A(new_n294), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n385), .A2(new_n389), .A3(new_n386), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n389), .B1(new_n385), .B2(new_n386), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n383), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n381), .B1(new_n432), .B2(G68), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n429), .B1(new_n433), .B2(KEYINPUT16), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n427), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n411), .B(new_n354), .C1(new_n412), .C2(new_n414), .ZN(new_n436));
  INV_X1    g0236(.A(G169), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n404), .B2(new_n409), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n426), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n399), .A2(new_n419), .ZN(new_n441));
  INV_X1    g0241(.A(new_n439), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(KEYINPUT18), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n375), .A2(new_n354), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n372), .A2(new_n437), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n366), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n425), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n357), .A2(new_n377), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n269), .A2(new_n451), .A3(G45), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(G270), .A3(new_n401), .ZN(new_n453));
  INV_X1    g0253(.A(G45), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n266), .B2(new_n268), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(G274), .A3(new_n401), .A4(new_n451), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G264), .A2(G1698), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n334), .B(new_n458), .C1(new_n214), .C2(G1698), .ZN(new_n459));
  INV_X1    g0259(.A(G303), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n339), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n263), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n437), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n293), .A2(new_n234), .B1(G20), .B2(new_n216), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n235), .C1(G33), .C2(new_n213), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n464), .A2(KEYINPUT20), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT20), .B1(new_n464), .B2(new_n466), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n467), .A2(new_n468), .B1(G116), .B2(new_n417), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n294), .B1(new_n269), .B2(G33), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n470), .A2(G116), .A3(new_n417), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT78), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n216), .A2(G20), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n466), .A2(new_n294), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n464), .A2(KEYINPUT20), .A3(new_n466), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n477), .A2(new_n478), .B1(new_n216), .B2(new_n300), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n470), .A2(G116), .A3(new_n417), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT78), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n463), .B1(new_n473), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT21), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n462), .A2(G179), .A3(new_n453), .A4(new_n456), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n472), .B1(new_n469), .B2(new_n471), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n479), .A2(KEYINPUT78), .A3(new_n480), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n487), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(KEYINPUT21), .A3(new_n463), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n462), .A2(new_n453), .A3(new_n456), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G190), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(G200), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(new_n486), .A3(new_n495), .A4(new_n487), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n484), .A2(new_n489), .A3(new_n491), .A4(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n235), .B1(new_n261), .B2(new_n498), .ZN(new_n499));
  NOR4_X1   g0299(.A1(KEYINPUT76), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT76), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G87), .A2(G97), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n252), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n499), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT77), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT19), .B1(new_n288), .B2(G97), .ZN(new_n507));
  AOI21_X1  g0307(.A(G20), .B1(new_n332), .B2(new_n333), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(G68), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(KEYINPUT77), .B(new_n499), .C1(new_n500), .C2(new_n503), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n294), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n300), .A2(new_n358), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n470), .A2(new_n417), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT74), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT74), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n470), .A2(new_n516), .A3(new_n417), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n359), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n512), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(G250), .B1(new_n402), .B2(new_n454), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n269), .A2(G45), .A3(G274), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n401), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n220), .A2(new_n259), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n227), .A2(G1698), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n525), .C1(new_n256), .C2(new_n257), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n401), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n437), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n263), .B1(new_n520), .B2(new_n521), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n531), .A2(new_n354), .A3(new_n528), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n519), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n511), .A2(new_n294), .B1(new_n300), .B2(new_n358), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n523), .A2(new_n529), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n531), .A2(new_n528), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G190), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n515), .A2(G87), .A3(new_n517), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n534), .A2(new_n536), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n497), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT85), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n452), .A2(G264), .A3(new_n401), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT84), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n263), .B1(new_n455), .B2(new_n451), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(KEYINPUT84), .A3(G264), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n214), .A2(G1698), .ZN(new_n550));
  OAI221_X1 g0350(.A(new_n550), .B1(G250), .B2(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G294), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n401), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n543), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  AOI211_X1 g0355(.A(KEYINPUT85), .B(new_n553), .C1(new_n546), .C2(new_n548), .ZN(new_n556));
  OAI211_X1 g0356(.A(G179), .B(new_n456), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n544), .A2(new_n545), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT84), .B1(new_n547), .B2(G264), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(KEYINPUT83), .B2(new_n554), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT83), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n456), .B1(new_n553), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(G169), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT25), .ZN(new_n565));
  AOI211_X1 g0365(.A(KEYINPUT82), .B(new_n565), .C1(new_n300), .C2(new_n252), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(KEYINPUT82), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n565), .A2(KEYINPUT82), .ZN(new_n568));
  NOR4_X1   g0368(.A1(new_n417), .A2(G107), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n515), .A2(new_n517), .ZN(new_n570));
  AOI211_X1 g0370(.A(new_n566), .B(new_n569), .C1(new_n570), .C2(G107), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n235), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n334), .A2(KEYINPUT22), .A3(new_n235), .A4(G87), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g0376(.A(KEYINPUT79), .B(KEYINPUT24), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n288), .A2(G116), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT80), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n580), .A2(new_n252), .A3(KEYINPUT23), .A4(G20), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n580), .A2(KEYINPUT23), .B1(new_n235), .B2(G107), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n580), .A2(KEYINPUT23), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n576), .A2(new_n578), .A3(new_n579), .A4(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n574), .A2(new_n575), .A3(new_n579), .A4(new_n584), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n577), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT81), .B1(new_n588), .B2(new_n294), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT81), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n590), .B(new_n429), .C1(new_n585), .C2(new_n587), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n571), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n564), .A2(new_n592), .ZN(new_n593));
  OR3_X1    g0393(.A1(new_n560), .A2(G190), .A3(new_n562), .ZN(new_n594));
  INV_X1    g0394(.A(new_n456), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT85), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n549), .A2(new_n543), .A3(new_n554), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n594), .B1(new_n599), .B2(G200), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n570), .A2(G107), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n566), .A2(new_n569), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n588), .A2(new_n294), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n590), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n588), .A2(KEYINPUT81), .A3(new_n294), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT75), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n212), .B1(new_n332), .B2(new_n333), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT4), .ZN(new_n611));
  OAI21_X1  g0411(.A(G1698), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(G244), .B1(new_n256), .B2(new_n257), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n613), .A2(new_n611), .B1(G33), .B2(G283), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n334), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n595), .B1(new_n616), .B2(new_n263), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n547), .A2(G257), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n609), .B1(new_n619), .B2(G200), .ZN(new_n620));
  AOI211_X1 g0420(.A(KEYINPUT75), .B(new_n284), .C1(new_n617), .C2(new_n618), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n619), .A2(new_n373), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT6), .ZN(new_n624));
  AND2_X1   g0424(.A1(G97), .A2(G107), .ZN(new_n625));
  NOR2_X1   g0425(.A1(G97), .A2(G107), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n252), .A2(KEYINPUT6), .A3(G97), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n235), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n291), .A2(new_n226), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT73), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n387), .A2(new_n383), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G107), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT73), .ZN(new_n634));
  INV_X1    g0434(.A(new_n630), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n252), .A2(KEYINPUT6), .A3(G97), .ZN(new_n636));
  XNOR2_X1  g0436(.A(G97), .B(G107), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n624), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n634), .B(new_n635), .C1(new_n638), .C2(new_n235), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n631), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n294), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n300), .A2(new_n213), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n515), .A2(G97), .A3(new_n517), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n623), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n617), .A2(new_n354), .A3(new_n618), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(G169), .B1(new_n617), .B2(new_n618), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n622), .A2(new_n645), .B1(new_n649), .B2(new_n644), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n542), .A2(new_n593), .A3(new_n608), .A4(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n450), .A2(new_n651), .ZN(G372));
  NAND4_X1  g0452(.A1(new_n649), .A2(new_n533), .A3(new_n540), .A4(new_n644), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT26), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT86), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n530), .B2(new_n532), .ZN(new_n656));
  OAI21_X1  g0456(.A(G169), .B1(new_n531), .B2(new_n528), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n657), .B(KEYINPUT86), .C1(new_n535), .C2(new_n354), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n656), .A2(new_n658), .B1(new_n534), .B2(new_n518), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n649), .A2(new_n644), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n490), .A2(KEYINPUT21), .A3(new_n463), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT21), .B1(new_n490), .B2(new_n463), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n663), .A2(new_n664), .A3(new_n488), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n593), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n662), .B1(new_n666), .B2(new_n608), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n668));
  AOI221_X4 g0468(.A(new_n595), .B1(G257), .B2(new_n547), .C1(new_n616), .C2(new_n263), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT75), .B1(new_n669), .B2(new_n284), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(G190), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n619), .A2(new_n609), .A3(G200), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n668), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(new_n540), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n654), .B(new_n660), .C1(new_n667), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n449), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n447), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n310), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n424), .B1(new_n679), .B2(new_n318), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT18), .B1(new_n441), .B2(new_n442), .ZN(new_n681));
  AOI211_X1 g0481(.A(new_n426), .B(new_n439), .C1(new_n399), .C2(new_n419), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n353), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n677), .A2(new_n684), .A3(new_n356), .ZN(G369));
  AND2_X1   g0485(.A1(new_n608), .A2(new_n593), .ZN(new_n686));
  INV_X1    g0486(.A(G213), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n299), .A2(G20), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n269), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n689), .B2(KEYINPUT27), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n269), .A2(new_n691), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT87), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT87), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n269), .A2(new_n694), .A3(new_n691), .A4(new_n688), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n690), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT88), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT88), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  OR3_X1    g0500(.A1(new_n699), .A2(KEYINPUT89), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT89), .B1(new_n699), .B2(new_n700), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n686), .B1(new_n607), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n564), .A3(new_n592), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n704), .B(new_n706), .C1(new_n665), .C2(new_n705), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(new_n490), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n665), .A3(new_n496), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n484), .A2(new_n489), .A3(new_n491), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n490), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n708), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n686), .A2(new_n711), .A3(new_n703), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n707), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n593), .A2(new_n665), .B1(new_n607), .B2(new_n600), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n703), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(G399));
  NAND2_X1  g0518(.A1(new_n208), .A2(new_n400), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(KEYINPUT90), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(KEYINPUT90), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n500), .A2(new_n503), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n216), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n722), .A2(new_n265), .A3(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT91), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(KEYINPUT91), .ZN(new_n727));
  INV_X1    g0527(.A(new_n722), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n726), .B(new_n727), .C1(new_n237), .C2(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT94), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n619), .A2(new_n437), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n540), .A2(new_n644), .A3(new_n732), .A4(new_n646), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT26), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n734), .B(new_n660), .C1(new_n653), .C2(KEYINPUT26), .ZN(new_n735));
  AND4_X1   g0535(.A1(new_n534), .A2(new_n536), .A3(new_n538), .A4(new_n539), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n659), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n673), .A3(new_n661), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n735), .B1(new_n716), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n731), .B1(new_n740), .B2(new_n705), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n711), .B1(new_n564), .B2(new_n592), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n456), .B1(new_n555), .B2(new_n556), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n284), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n592), .B1(new_n594), .B2(new_n744), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n742), .A2(new_n745), .A3(new_n738), .ZN(new_n746));
  OAI211_X1 g0546(.A(KEYINPUT94), .B(new_n703), .C1(new_n746), .C2(new_n735), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n741), .A2(new_n747), .A3(KEYINPUT29), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n676), .A2(new_n749), .A3(new_n703), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT30), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n537), .B(new_n669), .C1(new_n555), .C2(new_n556), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n485), .B(KEYINPUT92), .Z(new_n754));
  OAI21_X1  g0554(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n535), .B1(new_n597), .B2(new_n598), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n485), .B(KEYINPUT92), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(KEYINPUT30), .A3(new_n669), .A4(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n669), .A2(G179), .A3(new_n493), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n743), .A2(new_n759), .A3(new_n535), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n755), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n705), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT31), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT93), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n686), .A2(new_n542), .A3(new_n650), .A4(new_n703), .ZN(new_n768));
  AOI21_X1  g0568(.A(KEYINPUT31), .B1(new_n761), .B2(new_n705), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n751), .B1(G330), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n730), .B1(new_n772), .B2(G1), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT95), .ZN(G364));
  AOI21_X1  g0574(.A(new_n265), .B1(new_n688), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n722), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n373), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n235), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G97), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n235), .A2(new_n354), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(G190), .A3(new_n284), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n782), .B1(new_n229), .B2(new_n784), .C1(new_n226), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n235), .A2(G179), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n785), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G159), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n339), .B(new_n787), .C1(KEYINPUT32), .C2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(KEYINPUT97), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n793), .A2(KEYINPUT97), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n788), .A2(new_n373), .A3(G200), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n224), .B1(new_n252), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n783), .A2(new_n373), .A3(G200), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n799), .B1(G68), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n792), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n788), .A2(G190), .A3(G200), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(KEYINPUT32), .B2(new_n791), .C1(new_n211), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n798), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n339), .B1(new_n786), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(G329), .C2(new_n790), .ZN(new_n810));
  INV_X1    g0610(.A(new_n804), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G303), .ZN(new_n812));
  INV_X1    g0612(.A(G317), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(KEYINPUT33), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(KEYINPUT33), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n800), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G294), .B2(new_n781), .ZN(new_n817));
  AND3_X1   g0617(.A1(new_n810), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G322), .ZN(new_n819));
  INV_X1    g0619(.A(G326), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n819), .B2(new_n784), .C1(new_n820), .C2(new_n797), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n805), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT98), .Z(new_n823));
  AOI21_X1  g0623(.A(new_n234), .B1(G20), .B2(new_n437), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n778), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(G13), .A2(G33), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G20), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n824), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n208), .A2(new_n334), .ZN(new_n830));
  INV_X1    g0630(.A(G355), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n830), .A2(new_n831), .B1(G116), .B2(new_n208), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT96), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n208), .A2(new_n339), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(G45), .B2(new_n237), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n250), .B2(G45), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n829), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n710), .A2(new_n712), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n828), .B(KEYINPUT99), .Z(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n825), .B(new_n838), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n713), .A2(new_n777), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(G330), .B2(new_n839), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(G396));
  INV_X1    g0645(.A(KEYINPUT101), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n447), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n445), .A2(KEYINPUT101), .A3(new_n366), .A4(new_n446), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n705), .A2(new_n366), .ZN(new_n850));
  INV_X1    g0650(.A(new_n377), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n676), .A2(new_n703), .A3(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n676), .A2(new_n703), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n705), .A2(new_n678), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n771), .A2(G330), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n778), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT102), .Z(new_n861));
  NAND2_X1  g0661(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n782), .B1(new_n252), .B2(new_n804), .C1(new_n808), .C2(new_n789), .ZN(new_n864));
  INV_X1    g0664(.A(new_n797), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n865), .A2(G303), .B1(G283), .B2(new_n801), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n216), .B2(new_n786), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT100), .ZN(new_n868));
  INV_X1    g0668(.A(G294), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n868), .B(new_n339), .C1(new_n869), .C2(new_n784), .ZN(new_n870));
  INV_X1    g0670(.A(new_n798), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n864), .B(new_n870), .C1(G87), .C2(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n865), .A2(G137), .B1(G150), .B2(new_n801), .ZN(new_n873));
  INV_X1    g0673(.A(new_n784), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(G143), .ZN(new_n875));
  INV_X1    g0675(.A(G159), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n873), .B(new_n875), .C1(new_n876), .C2(new_n786), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT34), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n877), .A2(new_n878), .B1(G50), .B2(new_n811), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n871), .A2(G68), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n879), .B(new_n880), .C1(new_n229), .C2(new_n780), .ZN(new_n881));
  INV_X1    g0681(.A(G132), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n877), .A2(new_n878), .B1(new_n882), .B2(new_n789), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n881), .A2(new_n339), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n824), .B1(new_n872), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n824), .A2(new_n826), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n226), .ZN(new_n887));
  INV_X1    g0687(.A(new_n857), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n826), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n885), .A2(new_n777), .A3(new_n887), .A4(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n863), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(G384));
  INV_X1    g0692(.A(KEYINPUT108), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n764), .B(new_n767), .C1(new_n651), .C2(new_n705), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n857), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n308), .B1(new_n307), .B2(new_n286), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n373), .B1(new_n280), .B2(new_n281), .ZN(new_n897));
  NOR4_X1   g0697(.A1(new_n897), .A2(new_n303), .A3(KEYINPUT69), .A4(new_n285), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n318), .B(KEYINPUT104), .C1(new_n896), .C2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n304), .B1(new_n701), .B2(new_n702), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n317), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n310), .A2(KEYINPUT104), .A3(new_n903), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n893), .B1(new_n895), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  INV_X1    g0708(.A(new_n699), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n441), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT106), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n435), .A2(new_n439), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n699), .B1(new_n399), .B2(new_n419), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n416), .B2(new_n435), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n912), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n915), .B2(KEYINPUT106), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n910), .A2(new_n420), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(new_n913), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n910), .B1(new_n425), .B2(new_n444), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n907), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n434), .B1(KEYINPUT16), .B2(new_n433), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n419), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n909), .B(new_n925), .C1(new_n683), .C2(new_n424), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n908), .B1(new_n919), .B2(new_n913), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n442), .B2(new_n909), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(KEYINPUT37), .A3(new_n420), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n926), .A2(KEYINPUT38), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n923), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n900), .B(KEYINPUT104), .C1(new_n896), .C2(new_n898), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n933), .A2(new_n903), .B1(new_n899), .B2(new_n901), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n893), .A2(KEYINPUT40), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n934), .A2(new_n894), .A3(new_n857), .A4(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n906), .A2(new_n931), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT40), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n939));
  AND4_X1   g0739(.A1(new_n542), .A2(new_n593), .A3(new_n608), .A4(new_n650), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(new_n703), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n888), .B1(new_n941), .B2(new_n764), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n907), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n930), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n942), .A2(new_n945), .A3(new_n934), .A4(new_n935), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n449), .A2(new_n894), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n947), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(G330), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT109), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT107), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n684), .A2(new_n356), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n751), .B2(new_n449), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT39), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n931), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n944), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n703), .A2(new_n303), .A3(new_n317), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT105), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n683), .A2(new_n699), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n849), .A2(new_n705), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n854), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n968), .A2(new_n945), .A3(new_n934), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n957), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n954), .A2(new_n956), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n954), .A2(new_n956), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n973), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n972), .B(new_n975), .C1(new_n269), .C2(new_n688), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n237), .A2(new_n226), .A3(new_n378), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n201), .A2(new_n219), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n299), .B(new_n402), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n638), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n216), .B1(new_n980), .B2(KEYINPUT35), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n981), .B(new_n236), .C1(KEYINPUT35), .C2(new_n980), .ZN(new_n982));
  XOR2_X1   g0782(.A(KEYINPUT103), .B(KEYINPUT36), .Z(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n976), .A2(new_n979), .A3(new_n984), .ZN(G367));
  XOR2_X1   g0785(.A(new_n722), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n707), .A2(new_n714), .ZN(new_n988));
  INV_X1    g0788(.A(new_n713), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n715), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n772), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n650), .B1(new_n703), .B2(new_n668), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n661), .B2(new_n703), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n995), .A2(KEYINPUT45), .A3(new_n717), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT45), .B1(new_n995), .B2(new_n717), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n673), .A2(new_n661), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n716), .A2(new_n999), .A3(new_n703), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT44), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n715), .ZN(new_n1003));
  AND3_X1   g0803(.A1(new_n1002), .A2(KEYINPUT110), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1003), .B1(new_n1002), .B2(KEYINPUT110), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n993), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n772), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n987), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n775), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n714), .A2(new_n999), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT42), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n661), .B1(new_n994), .B2(new_n593), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n703), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n534), .A2(new_n539), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n705), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(new_n660), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n737), .B2(new_n1016), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1003), .A2(new_n995), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT43), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1014), .A2(new_n1022), .A3(new_n1020), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1018), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(KEYINPUT43), .B2(new_n1019), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1009), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G150), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n334), .B1(new_n784), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n780), .A2(new_n219), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G159), .B2(new_n801), .ZN(new_n1034));
  INV_X1    g0834(.A(G137), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n789), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1032), .B(new_n1036), .C1(G143), .C2(new_n865), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n871), .A2(G77), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n229), .C2(new_n804), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n786), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(new_n201), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n804), .A2(new_n216), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1042), .A2(KEYINPUT46), .B1(new_n874), .B2(G303), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(KEYINPUT46), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n781), .A2(G107), .B1(new_n1040), .B2(G283), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n801), .A2(G294), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n339), .B1(new_n789), .B2(new_n813), .C1(new_n213), .C2(new_n798), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT111), .Z(new_n1049));
  AOI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(G311), .C2(new_n865), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1041), .A2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT47), .Z(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n824), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n829), .B1(new_n208), .B2(new_n358), .C1(new_n246), .C2(new_n834), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n1053), .A2(new_n777), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1018), .A2(new_n840), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1030), .A2(KEYINPUT112), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT112), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1029), .A2(new_n1027), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n775), .B2(new_n1008), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1057), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1058), .A2(new_n1063), .ZN(G387));
  NAND2_X1  g0864(.A1(new_n865), .A2(G159), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n784), .A2(new_n224), .B1(new_n798), .B2(new_n213), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n339), .B(new_n1066), .C1(G68), .C2(new_n1040), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n811), .A2(G77), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n789), .A2(new_n1031), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n780), .A2(new_n358), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n319), .C2(new_n801), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n865), .A2(G322), .B1(G311), .B2(new_n801), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n460), .B2(new_n786), .C1(new_n813), .C2(new_n784), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT48), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n806), .B2(new_n780), .C1(new_n869), .C2(new_n804), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT49), .Z(new_n1077));
  OAI221_X1 g0877(.A(new_n339), .B1(new_n789), .B2(new_n820), .C1(new_n216), .C2(new_n798), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1072), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n824), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n724), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1081), .A2(KEYINPUT114), .B1(G68), .B2(G77), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1082), .B(new_n454), .C1(KEYINPUT114), .C2(new_n1081), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n319), .A2(new_n224), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT50), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n835), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT115), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n243), .A2(G45), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT113), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(G107), .B2(new_n208), .C1(new_n1081), .C2(new_n830), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n829), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n704), .A2(new_n706), .A3(new_n840), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1080), .A2(new_n777), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n993), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n722), .B1(new_n772), .B2(new_n992), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1094), .B1(new_n775), .B2(new_n991), .C1(new_n1095), .C2(new_n1096), .ZN(G393));
  INV_X1    g0897(.A(new_n1002), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(new_n715), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1006), .B1(new_n993), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n722), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1099), .A2(new_n775), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n254), .A2(new_n835), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n829), .C1(new_n213), .C2(new_n208), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n995), .A2(G20), .A3(new_n827), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n797), .A2(new_n813), .B1(new_n808), .B2(new_n784), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT52), .Z(new_n1107));
  AOI211_X1 g0907(.A(new_n334), .B(new_n1107), .C1(G116), .C2(new_n781), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n460), .B2(new_n800), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n789), .A2(new_n819), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n786), .A2(new_n869), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n252), .A2(new_n798), .B1(new_n804), .B2(new_n806), .ZN(new_n1112));
  NOR4_X1   g0912(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n804), .A2(new_n219), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n797), .A2(new_n1031), .B1(new_n876), .B2(new_n784), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT51), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n790), .A2(G143), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n339), .B1(new_n781), .B2(G77), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G87), .A2(new_n871), .B1(new_n1040), .B2(new_n319), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1114), .B(new_n1120), .C1(new_n201), .C2(new_n801), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n778), .B(new_n1105), .C1(new_n1122), .C2(new_n824), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1102), .B1(new_n1104), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1101), .A2(new_n1124), .ZN(G390));
  NAND3_X1  g0925(.A1(new_n771), .A2(G330), .A3(new_n857), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n905), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT117), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n942), .A2(new_n1128), .A3(G330), .A4(new_n934), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n767), .B1(new_n651), .B2(new_n705), .ZN(new_n1130));
  OAI211_X1 g0930(.A(G330), .B(new_n857), .C1(new_n1130), .C2(new_n769), .ZN(new_n1131));
  OAI21_X1  g0931(.A(KEYINPUT117), .B1(new_n1131), .B2(new_n905), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1127), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT116), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n902), .A2(new_n1134), .A3(new_n904), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n902), .B2(new_n904), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1131), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n771), .A2(G330), .A3(new_n857), .A4(new_n934), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n741), .A2(new_n747), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n966), .B1(new_n1140), .B2(new_n857), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1133), .A2(new_n968), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n449), .A2(G330), .A3(new_n894), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT118), .B1(new_n956), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n450), .B1(new_n748), .B2(new_n750), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT118), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1146), .A2(new_n955), .A3(new_n1143), .A4(new_n1147), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1142), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n962), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1136), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n934), .A2(new_n1134), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1150), .B(new_n931), .C1(new_n1141), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n959), .A2(new_n960), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n905), .B1(new_n854), .B2(new_n967), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n962), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1138), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1154), .A2(new_n1157), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n728), .B1(new_n1149), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1164), .B2(new_n1149), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n776), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1155), .A2(new_n826), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n886), .A2(new_n361), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n880), .B1(new_n211), .B2(new_n804), .C1(new_n216), .C2(new_n784), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n334), .B1(new_n865), .B2(G283), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G77), .A2(new_n781), .B1(new_n801), .B2(G107), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n213), .C2(new_n786), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1170), .B(new_n1173), .C1(G294), .C2(new_n790), .ZN(new_n1174));
  INV_X1    g0974(.A(G128), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n797), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n811), .A2(G150), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT53), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n339), .B1(new_n790), .B2(G125), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n882), .B2(new_n784), .C1(new_n1035), .C2(new_n800), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT54), .B(G143), .Z(new_n1181));
  AOI22_X1  g0981(.A1(new_n201), .A2(new_n871), .B1(new_n1040), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n876), .B2(new_n780), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1176), .A2(new_n1178), .A3(new_n1180), .A4(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n824), .B1(new_n1174), .B2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1168), .A2(new_n777), .A3(new_n1169), .A4(new_n1185), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1166), .A2(new_n1167), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(G378));
  NAND2_X1  g0988(.A1(new_n947), .A2(G330), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n353), .A2(new_n356), .ZN(new_n1190));
  XOR2_X1   g0990(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1191));
  XOR2_X1   g0991(.A(new_n1190), .B(new_n1191), .Z(new_n1192));
  AOI21_X1  g0992(.A(new_n699), .B1(new_n324), .B2(new_n323), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1192), .B(new_n1193), .Z(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n965), .B2(new_n969), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1192), .B(new_n1193), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1156), .A2(new_n945), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1196), .A2(new_n1197), .A3(new_n964), .A4(new_n963), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1189), .A2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n947), .A2(new_n1195), .A3(G330), .A4(new_n1198), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1159), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1158), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1205), .B2(new_n1162), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1203), .B1(new_n1206), .B2(new_n1142), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  OAI21_X1  g1009(.A(KEYINPUT120), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n728), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n956), .A2(new_n1144), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1147), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n956), .A2(KEYINPUT118), .A3(new_n1144), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1142), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1164), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT120), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1220), .A3(KEYINPUT57), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1210), .A2(new_n1211), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1202), .A2(new_n776), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n886), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n777), .B1(new_n201), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n224), .B1(new_n256), .B2(G41), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n784), .A2(new_n252), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n334), .B1(new_n1040), .B2(new_n359), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n213), .B2(new_n800), .C1(new_n806), .C2(new_n789), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(G116), .C2(new_n865), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1068), .B1(new_n229), .B2(new_n798), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(new_n1033), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n400), .A3(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT58), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n780), .A2(new_n1031), .B1(new_n784), .B2(new_n1175), .ZN(new_n1235));
  INV_X1    g1035(.A(G125), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n797), .A2(new_n1236), .B1(new_n1035), .B2(new_n786), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n811), .A2(new_n1181), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1235), .B(new_n1237), .C1(KEYINPUT119), .C2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(KEYINPUT119), .B2(new_n1238), .C1(new_n882), .C2(new_n800), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G41), .B1(new_n1240), .B2(KEYINPUT59), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G33), .B1(new_n790), .B2(G124), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n876), .C2(new_n798), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1226), .B(new_n1234), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1225), .B1(new_n1245), .B2(new_n824), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1194), .B2(new_n827), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1223), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1222), .A2(new_n1249), .ZN(G375));
  OR3_X1    g1050(.A1(new_n1142), .A2(KEYINPUT121), .A3(new_n775), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1153), .A2(new_n826), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n886), .A2(new_n219), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n334), .B1(new_n789), .B2(new_n1175), .C1(new_n1031), .C2(new_n786), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n801), .B2(new_n1181), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1035), .B2(new_n784), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n797), .A2(new_n882), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n804), .A2(new_n876), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n780), .A2(new_n224), .B1(new_n798), .B2(new_n229), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1038), .A2(new_n339), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT122), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n865), .A2(G294), .B1(G97), .B2(new_n811), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1040), .A2(G107), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1070), .B1(G283), .B2(new_n874), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(KEYINPUT123), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(KEYINPUT123), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1262), .B(new_n1268), .C1(G116), .C2(new_n801), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n790), .A2(G303), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1260), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT124), .Z(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n824), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1252), .A2(new_n777), .A3(new_n1253), .A4(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT121), .B1(new_n1142), .B2(new_n775), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1251), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1149), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1142), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n987), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(G381));
  NOR2_X1   g1081(.A1(G387), .A2(G381), .ZN(new_n1282));
  INV_X1    g1082(.A(G390), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1285), .A2(KEYINPUT125), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1220), .B1(new_n1219), .B2(KEYINPUT57), .ZN(new_n1287));
  NOR4_X1   g1087(.A1(new_n1217), .A2(new_n1218), .A3(KEYINPUT120), .A4(new_n1209), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1248), .B1(new_n1289), .B2(new_n1211), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1187), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1286), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1285), .A2(KEYINPUT125), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(G407));
  OAI211_X1 g1094(.A(G407), .B(G213), .C1(G343), .C2(new_n1291), .ZN(G409));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1279), .B1(new_n1149), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1215), .A2(KEYINPUT60), .A3(new_n1142), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n722), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT126), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT126), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1297), .A2(new_n1301), .A3(new_n722), .A4(new_n1298), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1277), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n891), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(G384), .A3(new_n1277), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n687), .A2(G343), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(G2897), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1305), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1308), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G384), .B1(new_n1303), .B2(new_n1277), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n891), .B(new_n1276), .C1(new_n1300), .C2(new_n1302), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1310), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1187), .B1(new_n1222), .B2(new_n1249), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1219), .A2(new_n987), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1187), .A2(new_n1249), .A3(new_n1316), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1315), .A2(new_n1307), .A3(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(KEYINPUT63), .B1(new_n1314), .B2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1307), .B1(G375), .B2(G378), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1187), .A2(new_n1249), .A3(new_n1316), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1323), .A2(KEYINPUT63), .A3(new_n1320), .A4(new_n1324), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(G393), .B(G396), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1283), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(G390), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1326), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT112), .B1(new_n1030), .B2(new_n1057), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1061), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1283), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1326), .B1(new_n1334), .B2(KEYINPUT127), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G390), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT127), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1329), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1331), .B1(new_n1335), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT61), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1325), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1322), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1307), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1343), .B(new_n1324), .C1(new_n1290), .C2(new_n1187), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT62), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1344), .A2(new_n1309), .A3(new_n1313), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT62), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1323), .A2(new_n1348), .A3(new_n1320), .A4(new_n1324), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1346), .A2(new_n1347), .A3(new_n1340), .A4(new_n1349), .ZN(new_n1350));
  AOI22_X1  g1150(.A1(new_n1334), .A2(KEYINPUT127), .B1(new_n1328), .B2(G390), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1326), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1352), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1330), .B1(new_n1351), .B2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1350), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1342), .A2(new_n1355), .ZN(G405));
  NAND2_X1  g1156(.A1(G375), .A2(G378), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1291), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1354), .A2(new_n1358), .ZN(new_n1359));
  AND2_X1   g1159(.A1(new_n1291), .A2(new_n1357), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1339), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1359), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(new_n1345), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1359), .A2(new_n1361), .A3(new_n1320), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(G402));
endmodule


