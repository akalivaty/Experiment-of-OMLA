

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(n729), .A2(n728), .ZN(n731) );
  INV_X1 U552 ( .A(KEYINPUT103), .ZN(n733) );
  INV_X1 U553 ( .A(KEYINPUT102), .ZN(n730) );
  XNOR2_X1 U554 ( .A(n731), .B(n730), .ZN(n745) );
  NOR2_X2 U555 ( .A1(n811), .A2(n813), .ZN(n716) );
  INV_X1 U556 ( .A(KEYINPUT71), .ZN(n580) );
  NOR2_X1 U557 ( .A1(G651), .A2(n652), .ZN(n654) );
  AND2_X2 U558 ( .A1(G2105), .A2(G2104), .ZN(n1004) );
  NOR2_X1 U559 ( .A1(n839), .A2(n838), .ZN(n840) );
  NOR2_X1 U560 ( .A1(n524), .A2(n523), .ZN(G164) );
  NOR2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  XOR2_X1 U562 ( .A(KEYINPUT17), .B(n514), .Z(n800) );
  NAND2_X1 U563 ( .A1(G138), .A2(n800), .ZN(n517) );
  INV_X1 U564 ( .A(G2105), .ZN(n518) );
  NAND2_X1 U565 ( .A1(n518), .A2(G2104), .ZN(n515) );
  XNOR2_X1 U566 ( .A(n515), .B(KEYINPUT65), .ZN(n627) );
  NAND2_X1 U567 ( .A1(G102), .A2(n627), .ZN(n516) );
  NAND2_X1 U568 ( .A1(n517), .A2(n516), .ZN(n524) );
  INV_X1 U569 ( .A(KEYINPUT89), .ZN(n522) );
  NOR2_X1 U570 ( .A1(G2104), .A2(n518), .ZN(n528) );
  NAND2_X1 U571 ( .A1(G126), .A2(n528), .ZN(n520) );
  NAND2_X1 U572 ( .A1(G114), .A2(n1004), .ZN(n519) );
  NAND2_X1 U573 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U574 ( .A(n522), .B(n521), .ZN(n523) );
  NAND2_X1 U575 ( .A1(n627), .A2(G101), .ZN(n527) );
  XNOR2_X1 U576 ( .A(KEYINPUT23), .B(KEYINPUT67), .ZN(n525) );
  XNOR2_X1 U577 ( .A(n525), .B(KEYINPUT66), .ZN(n526) );
  XNOR2_X1 U578 ( .A(n527), .B(n526), .ZN(n534) );
  AND2_X1 U579 ( .A1(G137), .A2(n800), .ZN(n532) );
  BUF_X1 U580 ( .A(n528), .Z(n1003) );
  NAND2_X1 U581 ( .A1(G125), .A2(n1003), .ZN(n530) );
  NAND2_X1 U582 ( .A1(G113), .A2(n1004), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(G160) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U587 ( .A1(G85), .A2(n643), .ZN(n536) );
  XOR2_X1 U588 ( .A(G543), .B(KEYINPUT0), .Z(n652) );
  INV_X1 U589 ( .A(G651), .ZN(n537) );
  NOR2_X1 U590 ( .A1(n652), .A2(n537), .ZN(n646) );
  NAND2_X1 U591 ( .A1(G72), .A2(n646), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n542) );
  NAND2_X1 U593 ( .A1(G47), .A2(n654), .ZN(n540) );
  NOR2_X1 U594 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n538), .Z(n577) );
  BUF_X1 U596 ( .A(n577), .Z(n658) );
  NAND2_X1 U597 ( .A1(G60), .A2(n658), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  OR2_X1 U599 ( .A1(n542), .A2(n541), .ZN(G290) );
  XNOR2_X1 U600 ( .A(G1348), .B(G2427), .ZN(n552) );
  XOR2_X1 U601 ( .A(G2443), .B(G2430), .Z(n544) );
  XNOR2_X1 U602 ( .A(G1341), .B(KEYINPUT108), .ZN(n543) );
  XNOR2_X1 U603 ( .A(n544), .B(n543), .ZN(n548) );
  XOR2_X1 U604 ( .A(G2435), .B(G2454), .Z(n546) );
  XNOR2_X1 U605 ( .A(KEYINPUT107), .B(G2438), .ZN(n545) );
  XNOR2_X1 U606 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U607 ( .A(n548), .B(n547), .Z(n550) );
  XNOR2_X1 U608 ( .A(G2451), .B(G2446), .ZN(n549) );
  XNOR2_X1 U609 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U610 ( .A(n552), .B(n551), .ZN(n553) );
  AND2_X1 U611 ( .A1(n553), .A2(G14), .ZN(G401) );
  NAND2_X1 U612 ( .A1(G52), .A2(n654), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G64), .A2(n658), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n643), .A2(G90), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n556), .B(KEYINPUT68), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G77), .A2(n646), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U620 ( .A1(n561), .A2(n560), .ZN(G171) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  NAND2_X1 U623 ( .A1(G75), .A2(n646), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G50), .A2(n654), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G88), .A2(n643), .ZN(n564) );
  XNOR2_X1 U627 ( .A(KEYINPUT83), .B(n564), .ZN(n565) );
  NOR2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n658), .A2(G62), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(G303) );
  INV_X1 U631 ( .A(G303), .ZN(G166) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n569) );
  XOR2_X1 U633 ( .A(n569), .B(KEYINPUT10), .Z(n1031) );
  NAND2_X1 U634 ( .A1(n1031), .A2(G567), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  XOR2_X1 U636 ( .A(G860), .B(KEYINPUT74), .Z(n617) );
  NAND2_X1 U637 ( .A1(n643), .A2(G81), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G68), .A2(n646), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT13), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G43), .A2(n654), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n579) );
  NAND2_X1 U645 ( .A1(G56), .A2(n577), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n579), .B(n578), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(KEYINPUT73), .B(n584), .ZN(n964) );
  OR2_X1 U650 ( .A1(n617), .A2(n964), .ZN(G153) );
  XNOR2_X1 U651 ( .A(G171), .B(KEYINPUT75), .ZN(G301) );
  NAND2_X1 U652 ( .A1(n658), .A2(G66), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n585), .B(KEYINPUT76), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G92), .A2(n643), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT77), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G79), .A2(n646), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G54), .A2(n654), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U660 ( .A(KEYINPUT78), .B(n591), .Z(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U662 ( .A(n594), .B(KEYINPUT15), .ZN(n965) );
  BUF_X1 U663 ( .A(n965), .Z(n634) );
  NOR2_X1 U664 ( .A1(n634), .A2(G868), .ZN(n595) );
  XNOR2_X1 U665 ( .A(n595), .B(KEYINPUT79), .ZN(n597) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(G284) );
  NAND2_X1 U668 ( .A1(n643), .A2(G89), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT4), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G76), .A2(n646), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT5), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G51), .A2(n654), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G63), .A2(n658), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT6), .B(n604), .Z(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U678 ( .A(n607), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U679 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U680 ( .A1(G53), .A2(n654), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G65), .A2(n658), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U683 ( .A1(G91), .A2(n643), .ZN(n611) );
  NAND2_X1 U684 ( .A1(G78), .A2(n646), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n710) );
  INV_X1 U687 ( .A(n710), .ZN(G299) );
  INV_X1 U688 ( .A(G868), .ZN(n671) );
  NOR2_X1 U689 ( .A1(G286), .A2(n671), .ZN(n615) );
  NOR2_X1 U690 ( .A1(G868), .A2(G299), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U692 ( .A(KEYINPUT80), .B(n616), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n617), .A2(G559), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n618), .A2(n634), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n619), .B(KEYINPUT16), .ZN(G148) );
  INV_X1 U696 ( .A(G559), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n620), .A2(n634), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n621), .A2(G868), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n964), .A2(n671), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U701 ( .A1(n1003), .A2(G123), .ZN(n624) );
  XNOR2_X1 U702 ( .A(n624), .B(KEYINPUT18), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G111), .A2(n1004), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n631) );
  BUF_X1 U705 ( .A(n800), .Z(n997) );
  NAND2_X1 U706 ( .A1(G135), .A2(n997), .ZN(n629) );
  BUF_X1 U707 ( .A(n627), .Z(n998) );
  NAND2_X1 U708 ( .A1(G99), .A2(n998), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n993) );
  XOR2_X1 U711 ( .A(G2096), .B(n993), .Z(n632) );
  NOR2_X1 U712 ( .A1(G2100), .A2(n632), .ZN(n633) );
  XNOR2_X1 U713 ( .A(KEYINPUT81), .B(n633), .ZN(G156) );
  NAND2_X1 U714 ( .A1(G559), .A2(n634), .ZN(n635) );
  XNOR2_X1 U715 ( .A(n635), .B(n964), .ZN(n661) );
  NOR2_X1 U716 ( .A1(n661), .A2(G860), .ZN(n642) );
  NAND2_X1 U717 ( .A1(G55), .A2(n654), .ZN(n637) );
  NAND2_X1 U718 ( .A1(G67), .A2(n658), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U720 ( .A1(G93), .A2(n643), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G80), .A2(n646), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n670) );
  XNOR2_X1 U724 ( .A(n642), .B(n670), .ZN(G145) );
  NAND2_X1 U725 ( .A1(G86), .A2(n643), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G48), .A2(n654), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n646), .A2(G73), .ZN(n647) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n647), .Z(n648) );
  NOR2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n658), .A2(G61), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n651), .A2(n650), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G87), .A2(n652), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n653), .B(KEYINPUT82), .ZN(n660) );
  NAND2_X1 U735 ( .A1(G49), .A2(n654), .ZN(n656) );
  NAND2_X1 U736 ( .A1(G74), .A2(G651), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U738 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(G288) );
  XNOR2_X1 U740 ( .A(KEYINPUT85), .B(n661), .ZN(n668) );
  XOR2_X1 U741 ( .A(G303), .B(G290), .Z(n662) );
  XNOR2_X1 U742 ( .A(n662), .B(G305), .ZN(n665) );
  XOR2_X1 U743 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n663) );
  XNOR2_X1 U744 ( .A(G288), .B(n663), .ZN(n664) );
  XOR2_X1 U745 ( .A(n665), .B(n664), .Z(n667) );
  XOR2_X1 U746 ( .A(G299), .B(n670), .Z(n666) );
  XNOR2_X1 U747 ( .A(n667), .B(n666), .ZN(n963) );
  XNOR2_X1 U748 ( .A(n668), .B(n963), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n669), .A2(G868), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U752 ( .A(KEYINPUT86), .B(n674), .Z(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U757 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XOR2_X1 U758 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  XNOR2_X1 U759 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n680) );
  XNOR2_X1 U762 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n679) );
  XNOR2_X1 U763 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U764 ( .A1(n681), .A2(G218), .ZN(n682) );
  NAND2_X1 U765 ( .A1(G96), .A2(n682), .ZN(n961) );
  NAND2_X1 U766 ( .A1(n961), .A2(G2106), .ZN(n686) );
  NAND2_X1 U767 ( .A1(G69), .A2(G120), .ZN(n683) );
  NOR2_X1 U768 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U769 ( .A1(G108), .A2(n684), .ZN(n962) );
  NAND2_X1 U770 ( .A1(n962), .A2(G567), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n686), .A2(n685), .ZN(n1030) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n687) );
  NOR2_X1 U773 ( .A1(n1030), .A2(n687), .ZN(n844) );
  NAND2_X1 U774 ( .A1(G36), .A2(n844), .ZN(n688) );
  XNOR2_X1 U775 ( .A(n688), .B(KEYINPUT88), .ZN(G176) );
  NOR2_X1 U776 ( .A1(G1384), .A2(G164), .ZN(n690) );
  INV_X1 U777 ( .A(KEYINPUT64), .ZN(n689) );
  XNOR2_X1 U778 ( .A(n690), .B(n689), .ZN(n811) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n813) );
  AND2_X1 U780 ( .A1(n716), .A2(G1996), .ZN(n691) );
  XOR2_X1 U781 ( .A(KEYINPUT26), .B(n691), .Z(n693) );
  INV_X1 U782 ( .A(n716), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n735), .A2(G1341), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U785 ( .A1(n964), .A2(n694), .ZN(n696) );
  NOR2_X1 U786 ( .A1(n696), .A2(n965), .ZN(n695) );
  XNOR2_X1 U787 ( .A(n695), .B(KEYINPUT100), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n696), .A2(n965), .ZN(n700) );
  NOR2_X1 U789 ( .A1(n716), .A2(G1348), .ZN(n698) );
  NOR2_X1 U790 ( .A1(G2067), .A2(n735), .ZN(n697) );
  NOR2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  AND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n701) );
  OR2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n707) );
  NAND2_X1 U794 ( .A1(n716), .A2(G2072), .ZN(n703) );
  XNOR2_X1 U795 ( .A(n703), .B(KEYINPUT27), .ZN(n705) );
  AND2_X1 U796 ( .A1(G1956), .A2(n735), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U798 ( .A1(n710), .A2(n709), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U800 ( .A(n708), .B(KEYINPUT101), .ZN(n713) );
  OR2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U802 ( .A(KEYINPUT28), .B(n711), .Z(n712) );
  NOR2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U804 ( .A(n714), .B(KEYINPUT29), .ZN(n720) );
  INV_X1 U805 ( .A(G1961), .ZN(n974) );
  NAND2_X1 U806 ( .A1(n735), .A2(n974), .ZN(n718) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .Z(n715) );
  XNOR2_X1 U808 ( .A(KEYINPUT99), .B(n715), .ZN(n884) );
  NAND2_X1 U809 ( .A1(n716), .A2(n884), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n724) );
  NAND2_X1 U811 ( .A1(G171), .A2(n724), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n729) );
  NAND2_X1 U813 ( .A1(G8), .A2(n735), .ZN(n779) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n779), .ZN(n746) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n735), .ZN(n744) );
  NOR2_X1 U816 ( .A1(n746), .A2(n744), .ZN(n721) );
  NAND2_X1 U817 ( .A1(G8), .A2(n721), .ZN(n722) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n722), .ZN(n723) );
  NOR2_X1 U819 ( .A1(G168), .A2(n723), .ZN(n726) );
  NOR2_X1 U820 ( .A1(G171), .A2(n724), .ZN(n725) );
  NOR2_X1 U821 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U822 ( .A(KEYINPUT31), .B(n727), .Z(n728) );
  INV_X1 U823 ( .A(n745), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n732), .A2(G286), .ZN(n734) );
  XNOR2_X1 U825 ( .A(n734), .B(n733), .ZN(n741) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n779), .ZN(n737) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U828 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U829 ( .A(KEYINPUT104), .B(n738), .ZN(n739) );
  NAND2_X1 U830 ( .A1(G303), .A2(n739), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U833 ( .A(n743), .B(KEYINPUT32), .ZN(n750) );
  NAND2_X1 U834 ( .A1(G8), .A2(n744), .ZN(n748) );
  NOR2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n769) );
  NOR2_X1 U838 ( .A1(G2090), .A2(G303), .ZN(n751) );
  NAND2_X1 U839 ( .A1(G8), .A2(n751), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n769), .A2(n752), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n753), .A2(n779), .ZN(n776) );
  INV_X1 U842 ( .A(G1971), .ZN(n972) );
  AND2_X1 U843 ( .A1(G166), .A2(n972), .ZN(n754) );
  NOR2_X1 U844 ( .A1(n754), .A2(KEYINPUT33), .ZN(n767) );
  OR2_X1 U845 ( .A1(G1981), .A2(G305), .ZN(n777) );
  NAND2_X1 U846 ( .A1(G1981), .A2(G305), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n777), .A2(n755), .ZN(n923) );
  AND2_X1 U848 ( .A1(n779), .A2(KEYINPUT105), .ZN(n756) );
  OR2_X1 U849 ( .A1(n923), .A2(n756), .ZN(n764) );
  NAND2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n911) );
  NOR2_X1 U851 ( .A1(KEYINPUT105), .A2(n779), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n911), .A2(n759), .ZN(n758) );
  INV_X1 U853 ( .A(KEYINPUT33), .ZN(n757) );
  NAND2_X1 U854 ( .A1(n758), .A2(n757), .ZN(n762) );
  NOR2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n914) );
  AND2_X1 U856 ( .A1(n914), .A2(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U857 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U858 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n770) );
  INV_X1 U860 ( .A(n770), .ZN(n765) );
  AND2_X1 U861 ( .A1(n765), .A2(n914), .ZN(n772) );
  INV_X1 U862 ( .A(n772), .ZN(n766) );
  AND2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U864 ( .A1(n769), .A2(n768), .ZN(n774) );
  NOR2_X1 U865 ( .A1(KEYINPUT105), .A2(n770), .ZN(n771) );
  OR2_X1 U866 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U868 ( .A1(n776), .A2(n775), .ZN(n828) );
  XNOR2_X1 U869 ( .A(n777), .B(KEYINPUT24), .ZN(n778) );
  NOR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n826) );
  NAND2_X1 U871 ( .A1(G140), .A2(n997), .ZN(n781) );
  NAND2_X1 U872 ( .A1(G104), .A2(n998), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U874 ( .A(KEYINPUT34), .B(n782), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G128), .A2(n1003), .ZN(n784) );
  NAND2_X1 U876 ( .A1(G116), .A2(n1004), .ZN(n783) );
  NAND2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U878 ( .A(KEYINPUT91), .B(n785), .ZN(n786) );
  XNOR2_X1 U879 ( .A(KEYINPUT35), .B(n786), .ZN(n787) );
  NOR2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U881 ( .A(n789), .B(KEYINPUT36), .ZN(n790) );
  XNOR2_X1 U882 ( .A(n790), .B(KEYINPUT92), .ZN(n1019) );
  XNOR2_X1 U883 ( .A(G2067), .B(KEYINPUT37), .ZN(n821) );
  NAND2_X1 U884 ( .A1(n1019), .A2(n821), .ZN(n856) );
  NAND2_X1 U885 ( .A1(G129), .A2(n1003), .ZN(n792) );
  NAND2_X1 U886 ( .A1(G117), .A2(n1004), .ZN(n791) );
  NAND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G105), .A2(n998), .ZN(n793) );
  XNOR2_X1 U889 ( .A(n793), .B(KEYINPUT38), .ZN(n794) );
  XNOR2_X1 U890 ( .A(n794), .B(KEYINPUT95), .ZN(n795) );
  NOR2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n997), .A2(G141), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n996) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n996), .ZN(n874) );
  NAND2_X1 U895 ( .A1(G1996), .A2(n996), .ZN(n799) );
  XOR2_X1 U896 ( .A(KEYINPUT96), .B(n799), .Z(n810) );
  NAND2_X1 U897 ( .A1(G131), .A2(n800), .ZN(n801) );
  XNOR2_X1 U898 ( .A(n801), .B(KEYINPUT94), .ZN(n804) );
  NAND2_X1 U899 ( .A1(G107), .A2(n1004), .ZN(n802) );
  XOR2_X1 U900 ( .A(KEYINPUT93), .B(n802), .Z(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U902 ( .A1(G119), .A2(n1003), .ZN(n806) );
  NAND2_X1 U903 ( .A1(G95), .A2(n998), .ZN(n805) );
  NAND2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n1017) );
  AND2_X1 U906 ( .A1(n1017), .A2(G1991), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n852) );
  INV_X1 U908 ( .A(n811), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U910 ( .A(KEYINPUT90), .B(n814), .ZN(n829) );
  XNOR2_X1 U911 ( .A(KEYINPUT97), .B(n829), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n852), .A2(n815), .ZN(n830) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n1017), .ZN(n859) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n859), .A2(n816), .ZN(n817) );
  NOR2_X1 U916 ( .A1(n830), .A2(n817), .ZN(n818) );
  NOR2_X1 U917 ( .A1(n874), .A2(n818), .ZN(n819) );
  XNOR2_X1 U918 ( .A(KEYINPUT39), .B(n819), .ZN(n820) );
  XNOR2_X1 U919 ( .A(n820), .B(KEYINPUT106), .ZN(n822) );
  NOR2_X1 U920 ( .A1(n1019), .A2(n821), .ZN(n854) );
  NAND2_X1 U921 ( .A1(n854), .A2(n829), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n822), .A2(n832), .ZN(n823) );
  NAND2_X1 U923 ( .A1(n856), .A2(n823), .ZN(n824) );
  NAND2_X1 U924 ( .A1(n824), .A2(n829), .ZN(n837) );
  INV_X1 U925 ( .A(n837), .ZN(n825) );
  OR2_X1 U926 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U927 ( .A1(n828), .A2(n827), .ZN(n839) );
  XNOR2_X1 U928 ( .A(G1986), .B(G290), .ZN(n909) );
  AND2_X1 U929 ( .A1(n909), .A2(n829), .ZN(n835) );
  INV_X1 U930 ( .A(n830), .ZN(n831) );
  NAND2_X1 U931 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n833), .B(KEYINPUT98), .ZN(n834) );
  OR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(n836) );
  AND2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n840), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U936 ( .A1(n1031), .A2(G2106), .ZN(n841) );
  XOR2_X1 U937 ( .A(KEYINPUT109), .B(n841), .Z(G217) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n842) );
  NAND2_X1 U939 ( .A1(G661), .A2(n842), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(G188) );
  NAND2_X1 U943 ( .A1(n1003), .A2(G124), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n845), .B(KEYINPUT44), .ZN(n847) );
  NAND2_X1 U945 ( .A1(G112), .A2(n1004), .ZN(n846) );
  NAND2_X1 U946 ( .A1(n847), .A2(n846), .ZN(n851) );
  NAND2_X1 U947 ( .A1(G136), .A2(n997), .ZN(n849) );
  NAND2_X1 U948 ( .A1(G100), .A2(n998), .ZN(n848) );
  NAND2_X1 U949 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U950 ( .A1(n851), .A2(n850), .ZN(G162) );
  INV_X1 U951 ( .A(n852), .ZN(n853) );
  NOR2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n861) );
  XOR2_X1 U953 ( .A(G2084), .B(G160), .Z(n855) );
  NOR2_X1 U954 ( .A1(n993), .A2(n855), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n860) );
  NAND2_X1 U957 ( .A1(n861), .A2(n860), .ZN(n879) );
  NAND2_X1 U958 ( .A1(G139), .A2(n997), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G103), .A2(n998), .ZN(n862) );
  NAND2_X1 U960 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U961 ( .A1(G127), .A2(n1003), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G115), .A2(n1004), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U964 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n994) );
  XOR2_X1 U966 ( .A(G2072), .B(n994), .Z(n870) );
  XOR2_X1 U967 ( .A(G164), .B(G2078), .Z(n869) );
  NOR2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U969 ( .A(KEYINPUT50), .B(n871), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n872), .B(KEYINPUT118), .ZN(n877) );
  XOR2_X1 U971 ( .A(G2090), .B(G162), .Z(n873) );
  NOR2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U973 ( .A(KEYINPUT51), .B(n875), .Z(n876) );
  NAND2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U975 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U976 ( .A(KEYINPUT52), .B(n880), .ZN(n881) );
  XNOR2_X1 U977 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n901) );
  NAND2_X1 U978 ( .A1(n881), .A2(n901), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n882), .A2(G29), .ZN(n959) );
  XNOR2_X1 U980 ( .A(G2090), .B(G35), .ZN(n896) );
  XOR2_X1 U981 ( .A(G25), .B(G1991), .Z(n883) );
  NAND2_X1 U982 ( .A1(n883), .A2(G28), .ZN(n893) );
  XOR2_X1 U983 ( .A(n884), .B(G27), .Z(n886) );
  XNOR2_X1 U984 ( .A(G1996), .B(G32), .ZN(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(KEYINPUT120), .B(n887), .ZN(n891) );
  XNOR2_X1 U987 ( .A(G2067), .B(G26), .ZN(n889) );
  XNOR2_X1 U988 ( .A(G33), .B(G2072), .ZN(n888) );
  NOR2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  NOR2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT53), .B(n894), .ZN(n895) );
  NOR2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n899) );
  XOR2_X1 U994 ( .A(G2084), .B(G34), .Z(n897) );
  XNOR2_X1 U995 ( .A(KEYINPUT54), .B(n897), .ZN(n898) );
  NAND2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n903) );
  INV_X1 U998 ( .A(G29), .ZN(n902) );
  NAND2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G11), .A2(n904), .ZN(n957) );
  INV_X1 U1001 ( .A(G16), .ZN(n953) );
  XOR2_X1 U1002 ( .A(n953), .B(KEYINPUT56), .Z(n928) );
  XOR2_X1 U1003 ( .A(G303), .B(KEYINPUT122), .Z(n905) );
  XOR2_X1 U1004 ( .A(n905), .B(G1971), .Z(n907) );
  XOR2_X1 U1005 ( .A(G171), .B(G1961), .Z(n906) );
  NOR2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n920) );
  XNOR2_X1 U1007 ( .A(G1348), .B(n965), .ZN(n916) );
  XOR2_X1 U1008 ( .A(G299), .B(G1956), .Z(n908) );
  XNOR2_X1 U1009 ( .A(n908), .B(KEYINPUT121), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(G1341), .B(n964), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(KEYINPUT123), .B(n921), .ZN(n926) );
  XOR2_X1 U1018 ( .A(G1966), .B(G168), .Z(n922) );
  NOR2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1020 ( .A(KEYINPUT57), .B(n924), .Z(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n955) );
  XOR2_X1 U1023 ( .A(G1986), .B(G24), .Z(n930) );
  XOR2_X1 U1024 ( .A(G1971), .B(G22), .Z(n929) );
  NAND2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(G23), .B(G1976), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(KEYINPUT58), .B(n933), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(n934), .B(KEYINPUT126), .ZN(n948) );
  XNOR2_X1 U1030 ( .A(G1966), .B(G21), .ZN(n946) );
  XNOR2_X1 U1031 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT60), .ZN(n944) );
  XOR2_X1 U1033 ( .A(G20), .B(G1956), .Z(n939) );
  XNOR2_X1 U1034 ( .A(G1341), .B(G19), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(G1981), .B(G6), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n942) );
  XOR2_X1 U1038 ( .A(KEYINPUT59), .B(G1348), .Z(n940) );
  XNOR2_X1 U1039 ( .A(G4), .B(n940), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(n944), .B(n943), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n950) );
  XOR2_X1 U1044 ( .A(G5), .B(n974), .Z(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT61), .B(n951), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1051 ( .A(KEYINPUT62), .B(n960), .Z(G311) );
  XNOR2_X1 U1052 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1053 ( .A(G120), .ZN(G236) );
  INV_X1 U1054 ( .A(G96), .ZN(G221) );
  INV_X1 U1055 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(G325) );
  INV_X1 U1057 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1058 ( .A(n964), .B(n963), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(G171), .B(n965), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n967), .B(n966), .ZN(n968) );
  XOR2_X1 U1061 ( .A(G286), .B(n968), .Z(n969) );
  NOR2_X1 U1062 ( .A1(G37), .A2(n969), .ZN(G397) );
  XOR2_X1 U1063 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n971) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G1976), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n971), .B(n970), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n973), .B(n972), .ZN(n976) );
  XOR2_X1 U1067 ( .A(n974), .B(G1956), .Z(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n980) );
  XOR2_X1 U1069 ( .A(KEYINPUT41), .B(G2474), .Z(n978) );
  XNOR2_X1 U1070 ( .A(G1991), .B(G1986), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(n978), .B(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(n980), .B(n979), .Z(n983) );
  INV_X1 U1073 ( .A(G1996), .ZN(n981) );
  XOR2_X1 U1074 ( .A(n981), .B(G1981), .Z(n982) );
  XNOR2_X1 U1075 ( .A(n983), .B(n982), .ZN(G229) );
  XOR2_X1 U1076 ( .A(G2100), .B(G2096), .Z(n985) );
  XNOR2_X1 U1077 ( .A(G2090), .B(KEYINPUT110), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n985), .B(n984), .ZN(n986) );
  XOR2_X1 U1079 ( .A(n986), .B(KEYINPUT42), .Z(n988) );
  XNOR2_X1 U1080 ( .A(G2072), .B(KEYINPUT43), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(n988), .B(n987), .ZN(n992) );
  XOR2_X1 U1082 ( .A(G2678), .B(G2084), .Z(n990) );
  XNOR2_X1 U1083 ( .A(G2067), .B(G2078), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(n992), .B(n991), .ZN(G227) );
  XOR2_X1 U1086 ( .A(n994), .B(n993), .Z(n995) );
  XNOR2_X1 U1087 ( .A(n996), .B(n995), .ZN(n1014) );
  XOR2_X1 U1088 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n1012) );
  NAND2_X1 U1089 ( .A1(G142), .A2(n997), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(G106), .A2(n998), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(KEYINPUT114), .B(KEYINPUT45), .Z(n1001) );
  XNOR2_X1 U1093 ( .A(n1002), .B(n1001), .ZN(n1009) );
  NAND2_X1 U1094 ( .A1(G130), .A2(n1003), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(G118), .A2(n1004), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1097 ( .A(KEYINPUT113), .B(n1007), .Z(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(n1010), .B(KEYINPUT115), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1012), .B(n1011), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(n1014), .B(n1013), .Z(n1016) );
  XNOR2_X1 U1102 ( .A(G164), .B(G162), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1016), .B(n1015), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(n1018), .B(n1017), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(G160), .B(n1019), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(G37), .A2(n1022), .ZN(G395) );
  NOR2_X1 U1108 ( .A1(G401), .A2(n1030), .ZN(n1027) );
  NOR2_X1 U1109 ( .A1(G229), .A2(G227), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(n1024), .B(n1023), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(G397), .A2(n1025), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(G395), .ZN(n1029) );
  XOR2_X1 U1115 ( .A(n1029), .B(KEYINPUT117), .Z(G308) );
  INV_X1 U1116 ( .A(G308), .ZN(G225) );
  INV_X1 U1117 ( .A(n1030), .ZN(G319) );
  INV_X1 U1118 ( .A(G108), .ZN(G238) );
  INV_X1 U1119 ( .A(n1031), .ZN(G223) );
endmodule

