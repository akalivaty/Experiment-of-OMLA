//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1339,
    new_n1340, new_n1341, new_n1342, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(new_n202), .A2(G50), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT64), .B(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G77), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n210), .B(new_n214), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n239), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G169), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G232), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  AOI21_X1  g0057(.A(G1), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND4_X1   g0058(.A1(new_n255), .A2(new_n258), .A3(new_n250), .A4(G274), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  AND2_X1   g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(new_n249), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n255), .B1(new_n262), .B2(new_n258), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n254), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n250), .A2(KEYINPUT69), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n261), .A2(new_n266), .A3(new_n249), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G223), .A2(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT73), .B1(new_n272), .B2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT73), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(G33), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n271), .A2(new_n273), .A3(new_n274), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G87), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n268), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n248), .B1(new_n264), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT76), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n258), .A2(new_n250), .A3(G274), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT67), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n262), .A2(new_n255), .A3(new_n258), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n284), .A2(new_n285), .B1(G232), .B2(new_n253), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n274), .A2(new_n277), .A3(new_n273), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n270), .A2(G1698), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(G223), .B2(G1698), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n279), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AND4_X1   g0091(.A1(new_n266), .A2(new_n249), .A3(G1), .A4(G13), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n266), .B1(new_n261), .B2(new_n249), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n286), .A2(new_n287), .A3(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n281), .A2(new_n282), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n282), .B1(new_n281), .B2(new_n296), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT16), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT64), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G68), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n201), .B1(new_n304), .B2(G58), .ZN(new_n305));
  INV_X1    g0105(.A(G159), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G20), .A2(G33), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n305), .A2(new_n208), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT7), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT3), .B(G33), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(G20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n276), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n273), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n216), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n300), .B1(new_n309), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n320), .A2(new_n207), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n288), .A2(new_n208), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT7), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n288), .A2(new_n310), .A3(new_n208), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(G68), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n308), .A2(new_n306), .ZN(new_n326));
  INV_X1    g0126(.A(G58), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n202), .B1(new_n216), .B2(new_n327), .ZN(new_n328));
  AOI211_X1 g0128(.A(new_n300), .B(new_n326), .C1(new_n328), .C2(G20), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n321), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  OAI211_X1 g0130(.A(KEYINPUT74), .B(new_n300), .C1(new_n309), .C2(new_n316), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n319), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(KEYINPUT8), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT8), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G58), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT70), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT70), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n321), .B1(G1), .B2(new_n208), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n339), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n344), .B1(new_n339), .B2(new_n343), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n332), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n299), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT18), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n299), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G200), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n264), .B2(new_n280), .ZN(new_n354));
  INV_X1    g0154(.A(G190), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n286), .A2(new_n355), .A3(new_n295), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n332), .A2(new_n347), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT17), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n332), .A2(new_n347), .A3(KEYINPUT17), .A4(new_n357), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n350), .A2(new_n352), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G223), .A2(G1698), .ZN(new_n364));
  INV_X1    g0164(.A(G222), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(G1698), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n311), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n219), .B2(new_n311), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n268), .B1(new_n368), .B2(KEYINPUT68), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(KEYINPUT68), .B2(new_n368), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n259), .A2(new_n263), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(G226), .B2(new_n253), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n374));
  INV_X1    g0174(.A(G150), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n308), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n272), .A2(G20), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(new_n341), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n321), .ZN(new_n379));
  INV_X1    g0179(.A(new_n338), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n240), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n342), .B2(new_n240), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n373), .A2(new_n353), .B1(new_n383), .B2(KEYINPUT9), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n381), .B1(new_n240), .B2(new_n342), .C1(new_n378), .C2(new_n321), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT9), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n370), .A2(new_n372), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n385), .A2(new_n386), .B1(new_n387), .B2(new_n355), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT10), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n389), .B(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n383), .B1(new_n248), .B2(new_n387), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(G179), .B2(new_n387), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n253), .A2(G238), .ZN(new_n396));
  NOR2_X1   g0196(.A1(G226), .A2(G1698), .ZN(new_n397));
  INV_X1    g0197(.A(G232), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(G1698), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n311), .B1(G33), .B2(G97), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n396), .B1(new_n400), .B2(new_n268), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT13), .B1(new_n401), .B2(new_n371), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G97), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n398), .A2(G1698), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G226), .B2(G1698), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n405), .B2(new_n314), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n294), .B1(G238), .B2(new_n253), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT13), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n284), .A2(new_n285), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G200), .ZN(new_n412));
  INV_X1    g0212(.A(new_n342), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT12), .ZN(new_n414));
  OAI21_X1  g0214(.A(G68), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n216), .A2(G20), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n377), .A2(G77), .B1(new_n307), .B2(G50), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n321), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT11), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n338), .A2(new_n414), .ZN(new_n421));
  INV_X1    g0221(.A(G13), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(G1), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT12), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n421), .B1(new_n416), .B2(new_n424), .C1(new_n418), .C2(KEYINPUT11), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n402), .A2(new_n410), .A3(G190), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n412), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n401), .A2(new_n371), .A3(KEYINPUT13), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n408), .B1(new_n407), .B2(new_n409), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n429), .B(G169), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT72), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(G169), .B1(new_n430), .B2(new_n431), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n411), .A2(KEYINPUT72), .A3(new_n429), .A4(G169), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n402), .A2(new_n410), .A3(G179), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n434), .A2(new_n436), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n426), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n428), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n219), .A2(new_n380), .ZN(new_n442));
  INV_X1    g0242(.A(G77), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n342), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n336), .A2(new_n307), .ZN(new_n445));
  INV_X1    g0245(.A(new_n377), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT15), .B(G87), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n445), .B1(new_n208), .B2(new_n219), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n321), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n217), .A2(G1698), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G232), .B2(G1698), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n311), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n294), .B(new_n453), .C1(G107), .C2(new_n311), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n253), .A2(G244), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n409), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT71), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT71), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n454), .A2(new_n458), .A3(new_n409), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n450), .B1(new_n460), .B2(new_n287), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n248), .A3(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n450), .B1(new_n460), .B2(new_n353), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n355), .B1(new_n457), .B2(new_n459), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AND4_X1   g0268(.A1(new_n363), .A2(new_n395), .A3(new_n441), .A4(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G238), .A2(G1698), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n218), .B2(G1698), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n471), .A2(new_n273), .A3(new_n274), .A4(new_n277), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G116), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n268), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n257), .A2(G1), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n260), .ZN(new_n476));
  INV_X1    g0276(.A(G250), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n257), .B2(G1), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n476), .A2(new_n250), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(G200), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n218), .A2(G1698), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G238), .B2(G1698), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n473), .B1(new_n288), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n294), .ZN(new_n484));
  INV_X1    g0284(.A(new_n479), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(G190), .A3(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n274), .A2(new_n277), .A3(new_n208), .A4(new_n273), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT19), .ZN(new_n488));
  INV_X1    g0288(.A(G87), .ZN(new_n489));
  INV_X1    g0289(.A(G97), .ZN(new_n490));
  INV_X1    g0290(.A(G107), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n403), .A2(new_n208), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND4_X1   g0294(.A1(new_n488), .A2(new_n208), .A3(G33), .A4(G97), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n242), .A2(new_n487), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n496), .A2(new_n449), .B1(new_n380), .B2(new_n447), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n251), .A2(G33), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n321), .A2(new_n338), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G87), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n480), .A2(new_n486), .A3(new_n497), .A4(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n487), .A2(new_n242), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n492), .A2(new_n493), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n495), .B1(new_n503), .B2(KEYINPUT19), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n449), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n447), .B(KEYINPUT79), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n499), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n447), .A2(new_n380), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n248), .B1(new_n474), .B2(new_n479), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n479), .B1(new_n483), .B2(new_n294), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n287), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n501), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n499), .A2(G97), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n380), .A2(new_n490), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(G97), .B(G107), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n519), .A2(new_n490), .A3(G107), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(G20), .B1(G77), .B2(new_n307), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n312), .A2(new_n315), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G107), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n517), .B1(new_n527), .B2(new_n449), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n251), .B(G45), .C1(new_n256), .C2(KEYINPUT5), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT77), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT5), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G41), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n475), .A2(KEYINPUT77), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n531), .A2(new_n534), .A3(new_n535), .A4(new_n262), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT78), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n250), .A2(G274), .A3(new_n535), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT78), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(new_n531), .A4(new_n534), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n218), .A2(G1698), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n274), .A2(new_n277), .A3(new_n273), .A4(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT4), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G283), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G250), .A2(G1698), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT4), .A2(G244), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(G1698), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n551), .B2(new_n314), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n294), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(G257), .A3(new_n250), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n542), .A2(new_n553), .A3(G190), .A4(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n542), .A2(new_n553), .A3(new_n555), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n528), .B(new_n556), .C1(new_n557), .C2(new_n353), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n542), .A2(new_n553), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n248), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n542), .A2(new_n553), .A3(new_n287), .A4(new_n555), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n521), .B1(new_n519), .B2(new_n518), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n562), .A2(new_n208), .B1(new_n443), .B2(new_n308), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n491), .B1(new_n312), .B2(new_n315), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n449), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(new_n516), .A3(new_n515), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n560), .A2(new_n561), .A3(new_n566), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n514), .A2(new_n558), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n554), .A2(G264), .A3(new_n250), .ZN(new_n569));
  INV_X1    g0369(.A(G257), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G1698), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G250), .B2(G1698), .ZN(new_n572));
  INV_X1    g0372(.A(G294), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n288), .A2(new_n572), .B1(new_n272), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n294), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n529), .A2(new_n530), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT77), .B1(new_n475), .B2(new_n533), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n540), .B1(new_n578), .B2(new_n539), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n536), .A2(KEYINPUT78), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n569), .B(new_n575), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(G179), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n248), .B2(new_n581), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT84), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT25), .ZN(new_n585));
  AOI211_X1 g0385(.A(G107), .B(new_n338), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n588), .A2(new_n589), .B1(G107), .B2(new_n499), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n208), .A2(G87), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT22), .B1(new_n311), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT23), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n208), .B2(G107), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n491), .A2(KEYINPUT23), .A3(G20), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT22), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n489), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n487), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g0404(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n600), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n601), .B1(new_n314), .B2(new_n591), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n473), .A2(G20), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n595), .B2(new_n596), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n487), .A2(new_n603), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n605), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT83), .B1(new_n614), .B2(new_n449), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n616), .B(new_n321), .C1(new_n607), .C2(new_n613), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n590), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n583), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n590), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n606), .B1(new_n600), .B2(new_n604), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n611), .A2(new_n612), .A3(new_n605), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n449), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n616), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n614), .A2(KEYINPUT83), .A3(new_n449), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n620), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n575), .A2(new_n569), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n627), .A2(KEYINPUT85), .A3(new_n355), .A4(new_n542), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT85), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n581), .B2(new_n353), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n581), .A2(G190), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n568), .A2(new_n619), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT81), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT80), .ZN(new_n636));
  INV_X1    g0436(.A(G116), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n320), .A2(new_n207), .B1(G20), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n547), .B(new_n208), .C1(G33), .C2(new_n490), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n638), .A2(KEYINPUT20), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT20), .B1(new_n638), .B2(new_n639), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n338), .A2(G116), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n321), .A2(new_n338), .A3(new_n498), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n637), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n636), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n643), .B1(new_n499), .B2(G116), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n638), .A2(new_n639), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT20), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n638), .A2(KEYINPUT20), .A3(new_n639), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n648), .A2(new_n653), .A3(KEYINPUT80), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n554), .A2(G270), .A3(new_n250), .ZN(new_n655));
  INV_X1    g0455(.A(G264), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G1698), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(G257), .B2(G1698), .ZN(new_n658));
  INV_X1    g0458(.A(G303), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n288), .A2(new_n658), .B1(new_n659), .B2(new_n311), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n294), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n542), .A2(new_n655), .A3(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n647), .B(new_n654), .C1(new_n662), .C2(new_n355), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n537), .A2(new_n541), .B1(new_n294), .B2(new_n660), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n353), .B1(new_n664), .B2(new_n655), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n635), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n665), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n647), .A2(new_n654), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n664), .A2(G190), .A3(new_n655), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT81), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n647), .A2(new_n654), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(KEYINPUT21), .A3(G169), .A4(new_n662), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n542), .A2(new_n655), .A3(new_n661), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n672), .A3(G179), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n248), .B1(new_n664), .B2(new_n655), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT21), .B1(new_n677), .B2(new_n672), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n671), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n634), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n469), .A2(new_n681), .ZN(G372));
  NAND2_X1  g0482(.A1(new_n360), .A2(new_n361), .ZN(new_n683));
  INV_X1    g0483(.A(new_n428), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n464), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n439), .A2(new_n440), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT87), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n350), .A2(new_n352), .ZN(new_n689));
  OR3_X1    g0489(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n687), .B2(new_n689), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n391), .A3(new_n691), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n692), .A2(KEYINPUT88), .A3(new_n393), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT88), .B1(new_n692), .B2(new_n393), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n469), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n501), .A2(new_n513), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n567), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n567), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n497), .A2(new_n500), .ZN(new_n700));
  OR3_X1    g0500(.A1(new_n511), .A2(KEYINPUT86), .A3(new_n353), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n480), .A2(KEYINPUT86), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n486), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n699), .A2(new_n513), .A3(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n513), .B(new_n698), .C1(new_n704), .C2(KEYINPUT26), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n513), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n558), .A2(new_n567), .ZN(new_n707));
  AOI211_X1 g0507(.A(new_n706), .B(new_n707), .C1(new_n626), .C2(new_n632), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n679), .A2(new_n619), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n695), .B1(new_n696), .B2(new_n710), .ZN(G369));
  AND2_X1   g0511(.A1(new_n633), .A2(new_n619), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n423), .A2(new_n208), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT27), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n423), .A2(new_n715), .A3(new_n208), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n714), .A2(G213), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT89), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(G343), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(G343), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n712), .B1(new_n626), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n619), .ZN(new_n725));
  INV_X1    g0525(.A(new_n723), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n671), .B(new_n679), .C1(new_n668), .C2(new_n723), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n677), .A2(new_n672), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT21), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n675), .A3(new_n673), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n672), .A3(new_n726), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT90), .B1(new_n735), .B2(G330), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT90), .ZN(new_n737));
  INV_X1    g0537(.A(G330), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n737), .B(new_n738), .C1(new_n729), .C2(new_n734), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n728), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n633), .A2(new_n733), .A3(new_n619), .A4(new_n723), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n725), .A2(new_n723), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n740), .A2(new_n744), .ZN(G399));
  INV_X1    g0545(.A(new_n212), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G41), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n492), .A2(G116), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(G1), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n205), .B2(new_n748), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT28), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n671), .A2(new_n679), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(new_n712), .A3(new_n568), .A4(new_n723), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT91), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n511), .A2(G179), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n662), .A2(new_n559), .A3(new_n581), .A4(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n511), .A2(new_n569), .A3(new_n575), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n674), .A2(G179), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n557), .A2(KEYINPUT30), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n662), .A2(new_n758), .A3(new_n287), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT30), .B1(new_n763), .B2(new_n557), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n755), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT30), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n760), .B2(new_n559), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n763), .A2(KEYINPUT30), .A3(new_n557), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n767), .A2(KEYINPUT91), .A3(new_n768), .A4(new_n757), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n765), .A2(new_n769), .A3(new_n726), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT31), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(KEYINPUT31), .B(new_n726), .C1(new_n762), .C2(new_n764), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n754), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G330), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT92), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT92), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n774), .A2(new_n777), .A3(G330), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT29), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n706), .B1(new_n626), .B2(new_n632), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n558), .A2(new_n567), .A3(KEYINPUT93), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT93), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n707), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n709), .A2(new_n781), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(KEYINPUT26), .B1(new_n706), .B2(new_n567), .ZN(new_n786));
  OR3_X1    g0586(.A1(new_n567), .A2(new_n697), .A3(KEYINPUT26), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n786), .A2(new_n787), .A3(new_n513), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n780), .B(new_n726), .C1(new_n785), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n708), .A2(new_n709), .ZN(new_n790));
  INV_X1    g0590(.A(new_n705), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n723), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n789), .B1(new_n780), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n779), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n752), .B1(new_n795), .B2(G1), .ZN(G364));
  NAND2_X1  g0596(.A1(new_n735), .A2(G330), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n737), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n735), .A2(KEYINPUT90), .A3(G330), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n422), .A2(G20), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n251), .B1(new_n802), .B2(G45), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n747), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n801), .B(new_n806), .C1(G330), .C2(new_n735), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n207), .B1(G20), .B2(new_n248), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n355), .A2(new_n353), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n810), .A2(G20), .A3(new_n287), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT97), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT97), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G87), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n208), .A2(new_n287), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT96), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT96), .B1(new_n208), .B2(new_n287), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n355), .A2(G200), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n816), .B1(new_n327), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n219), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G190), .A2(G200), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n819), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n823), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n208), .A2(G190), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n829), .A2(new_n287), .A3(new_n353), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n306), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT32), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n821), .A2(new_n287), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G20), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n490), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n208), .A2(new_n287), .A3(new_n353), .A4(G190), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n817), .A2(new_n810), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n311), .B1(new_n838), .B2(new_n242), .C1(new_n240), .C2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n829), .A2(new_n287), .A3(G200), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n836), .B(new_n841), .C1(G107), .C2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n828), .A2(new_n832), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n815), .A2(G303), .B1(G311), .B2(new_n827), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n835), .A2(new_n573), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n830), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(G329), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G317), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT33), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(KEYINPUT33), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n837), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n839), .A2(G326), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n855), .A3(new_n314), .ZN(new_n856));
  INV_X1    g0656(.A(new_n822), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(G322), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n846), .A2(new_n850), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n809), .B1(new_n845), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n311), .A2(G355), .A3(new_n212), .ZN(new_n861));
  INV_X1    g0661(.A(new_n288), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n746), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(G45), .B2(new_n205), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n246), .A2(new_n257), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n861), .B1(G116), .B2(new_n212), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(G13), .A2(G33), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(G20), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n808), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT94), .Z(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n806), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n873), .A2(KEYINPUT95), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n860), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n869), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n875), .B1(KEYINPUT95), .B2(new_n873), .C1(new_n735), .C2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n807), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(G396));
  INV_X1    g0679(.A(new_n779), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n461), .A2(new_n462), .A3(new_n723), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT98), .ZN(new_n883));
  INV_X1    g0683(.A(new_n450), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n726), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n450), .A2(KEYINPUT98), .A3(new_n723), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n465), .B2(new_n466), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n882), .B1(new_n463), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n723), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n792), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n793), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(new_n889), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n805), .B1(new_n880), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n880), .B2(new_n894), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n808), .A2(new_n867), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n806), .B1(new_n443), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n842), .A2(new_n489), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n899), .B(new_n836), .C1(G311), .C2(new_n849), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n314), .B1(new_n838), .B2(new_n847), .C1(new_n659), .C2(new_n840), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n814), .A2(new_n491), .B1(new_n637), .B2(new_n826), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n901), .B(new_n902), .C1(G294), .C2(new_n857), .ZN(new_n903));
  AOI22_X1  g0703(.A1(G137), .A2(new_n839), .B1(new_n837), .B2(G150), .ZN(new_n904));
  INV_X1    g0704(.A(G143), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n904), .B1(new_n905), .B2(new_n822), .C1(new_n306), .C2(new_n826), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT34), .ZN(new_n907));
  AOI22_X1  g0707(.A1(G132), .A2(new_n849), .B1(new_n834), .B2(G58), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n843), .A2(G68), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n862), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(G50), .B2(new_n815), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n900), .A2(new_n903), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n898), .B1(new_n809), .B2(new_n912), .C1(new_n889), .C2(new_n868), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n896), .A2(new_n913), .ZN(G384));
  NAND2_X1  g0714(.A1(new_n794), .A2(new_n469), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n695), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT101), .Z(new_n917));
  OAI211_X1 g0717(.A(new_n440), .B(new_n726), .C1(new_n439), .C2(new_n428), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n426), .A2(new_n723), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n428), .B(new_n920), .C1(new_n439), .C2(new_n440), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n892), .B2(new_n881), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n339), .A2(new_n343), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n324), .A2(G68), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n310), .B1(new_n288), .B2(new_n208), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n326), .B1(new_n328), .B2(G20), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT16), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n449), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT16), .B1(new_n325), .B2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n281), .A2(new_n296), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT76), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n281), .A2(new_n282), .A3(new_n296), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n718), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n358), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT37), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n348), .A2(new_n718), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT37), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n349), .A2(new_n940), .A3(new_n941), .A4(new_n358), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT99), .ZN(new_n944));
  INV_X1    g0744(.A(new_n937), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n362), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT99), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n939), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT38), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n944), .A2(new_n946), .A3(KEYINPUT38), .A4(new_n948), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n923), .A2(new_n953), .B1(new_n689), .B2(new_n717), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT39), .ZN(new_n955));
  AND4_X1   g0755(.A1(KEYINPUT38), .A2(new_n944), .A3(new_n948), .A4(new_n946), .ZN(new_n956));
  INV_X1    g0756(.A(new_n940), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT100), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n360), .A2(new_n958), .A3(new_n361), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(new_n350), .A3(new_n352), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n958), .B1(new_n360), .B2(new_n361), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n349), .A2(new_n940), .A3(new_n358), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT37), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n942), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT38), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n955), .B1(new_n956), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n951), .A2(KEYINPUT39), .A3(new_n952), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n686), .A2(new_n726), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n954), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n917), .B(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n889), .B1(new_n919), .B2(new_n921), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n681), .A2(new_n723), .B1(new_n771), .B2(new_n770), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n765), .A2(new_n769), .A3(KEYINPUT31), .A4(new_n726), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(KEYINPUT99), .A2(new_n943), .B1(new_n362), .B2(new_n945), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT38), .B1(new_n977), .B2(new_n948), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n976), .B1(new_n978), .B2(new_n956), .ZN(new_n979));
  XOR2_X1   g0779(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n956), .A2(new_n966), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n754), .A2(new_n772), .A3(new_n975), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n888), .A2(new_n463), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n881), .ZN(new_n986));
  INV_X1    g0786(.A(new_n920), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n441), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n986), .B1(new_n988), .B2(new_n918), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n984), .A2(KEYINPUT40), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n982), .B1(new_n983), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n469), .A2(new_n984), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n993), .A2(new_n994), .A3(new_n738), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n972), .A2(new_n995), .B1(new_n251), .B2(new_n802), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n972), .B2(new_n995), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n998), .A2(G116), .A3(new_n209), .A4(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT36), .Z(new_n1001));
  OAI211_X1 g0801(.A(new_n206), .B(new_n824), .C1(new_n327), .C2(new_n216), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n251), .B(G13), .C1(new_n1002), .C2(new_n241), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n997), .A2(new_n1001), .A3(new_n1003), .ZN(G367));
  NOR2_X1   g0804(.A1(new_n447), .A2(new_n212), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n871), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n235), .A2(new_n863), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n806), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n700), .A2(new_n723), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n513), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n706), .B2(new_n1009), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n311), .B1(new_n838), .B2(new_n306), .C1(new_n905), .C2(new_n840), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n814), .A2(new_n327), .B1(new_n375), .B2(new_n822), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G50), .C2(new_n827), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n835), .A2(new_n242), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n824), .B2(new_n843), .ZN(new_n1017));
  INV_X1    g0817(.A(G137), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1015), .B(new_n1017), .C1(new_n1018), .C2(new_n830), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT46), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n814), .A2(new_n1020), .A3(new_n637), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT109), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n835), .A2(new_n491), .B1(new_n842), .B2(new_n490), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n288), .B1(new_n826), .B2(new_n847), .C1(new_n573), .C2(new_n838), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(G317), .C2(new_n849), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1020), .B1(new_n814), .B2(new_n637), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1022), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n857), .A2(G303), .B1(G311), .B2(new_n839), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT108), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n1019), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT110), .Z(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT47), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1008), .B1(new_n876), .B2(new_n1012), .C1(new_n1032), .C2(new_n809), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n724), .A2(new_n727), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n798), .B2(new_n799), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT105), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n566), .A2(new_n726), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n784), .A2(new_n782), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n567), .A2(new_n723), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT103), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1038), .A2(KEYINPUT103), .A3(new_n1040), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1035), .A2(new_n1036), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(KEYINPUT105), .B1(new_n740), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n741), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1041), .A2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT42), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n699), .B1(new_n1045), .B2(new_n725), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n726), .B1(new_n1053), .B2(KEYINPUT104), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT104), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n619), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1056), .B2(new_n699), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1052), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1044), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT103), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n725), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1064), .A2(KEYINPUT104), .A3(new_n567), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1057), .A2(new_n1065), .A3(new_n723), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1052), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1068), .A2(new_n1046), .A3(new_n1048), .A4(new_n1059), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1071), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1061), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT45), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1041), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(new_n743), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n744), .A2(new_n1041), .A3(KEYINPUT45), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n744), .B2(new_n1041), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1077), .A2(new_n743), .A3(new_n1081), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1035), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1087), .A2(new_n740), .A3(new_n1084), .A4(new_n1083), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n733), .A2(new_n723), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1050), .B1(new_n1034), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(new_n800), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n795), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n747), .B(KEYINPUT41), .Z(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n803), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT107), .B1(new_n1075), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT107), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n804), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1033), .B1(new_n1098), .B2(new_n1101), .ZN(G387));
  INV_X1    g0902(.A(new_n795), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1103), .A2(new_n1092), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(new_n748), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1092), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1105), .B1(new_n795), .B2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n749), .A2(new_n746), .A3(new_n314), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n491), .B2(new_n746), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT111), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n232), .A2(new_n257), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n336), .A2(new_n240), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT50), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n749), .B(new_n257), .C1(new_n242), .C2(new_n443), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n863), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1110), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n806), .B1(new_n1116), .B2(new_n872), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n728), .B2(new_n876), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n814), .A2(new_n219), .B1(new_n337), .B2(new_n838), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G50), .B2(new_n857), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n490), .A2(new_n842), .B1(new_n830), .B2(new_n375), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n288), .B(new_n1121), .C1(G159), .C2(new_n839), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n506), .A2(new_n834), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n827), .A2(G68), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n815), .A2(G294), .B1(G283), .B2(new_n834), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G322), .A2(new_n839), .B1(new_n837), .B2(G311), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n659), .B2(new_n826), .C1(new_n851), .C2(new_n822), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT112), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1126), .B1(new_n1129), .B2(KEYINPUT48), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(KEYINPUT48), .B2(new_n1129), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT49), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT113), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n288), .B1(new_n842), .B2(new_n637), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G326), .B2(new_n849), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1125), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1118), .B1(new_n1138), .B2(new_n808), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1106), .B2(new_n804), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1107), .A2(new_n1140), .ZN(G393));
  INV_X1    g0941(.A(new_n1089), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n748), .B1(new_n1104), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1104), .B2(new_n1142), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1047), .A2(new_n869), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n872), .B1(new_n490), .B2(new_n212), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n239), .A2(new_n746), .A3(new_n862), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n805), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n862), .B1(new_n240), .B2(new_n838), .C1(new_n814), .C2(new_n216), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n336), .B2(new_n827), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n840), .A2(new_n375), .B1(new_n822), .B2(new_n306), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT51), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n830), .A2(new_n905), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n899), .B(new_n1153), .C1(G77), .C2(new_n834), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n857), .A2(G311), .B1(G317), .B2(new_n839), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT52), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n849), .A2(G322), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n814), .B2(new_n847), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT114), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n827), .A2(G294), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n314), .B1(new_n491), .B2(new_n842), .C1(new_n838), .C2(new_n659), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G116), .B2(new_n834), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1155), .B1(new_n1157), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1148), .B1(new_n1167), .B2(new_n808), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1142), .A2(new_n804), .B1(new_n1145), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1144), .A2(new_n1169), .ZN(G390));
  NAND3_X1  g0970(.A1(new_n984), .A2(G330), .A3(new_n989), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT115), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n986), .B1(new_n776), .B2(new_n778), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n922), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n881), .B1(new_n710), .B2(new_n890), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n779), .A2(new_n889), .A3(new_n1175), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n984), .A2(G330), .A3(new_n889), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n922), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n726), .B(new_n986), .C1(new_n785), .C2(new_n788), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n882), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1178), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n469), .A2(G330), .A3(new_n984), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n915), .B(new_n1187), .C1(new_n693), .C2(new_n694), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n967), .A2(new_n968), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1177), .A2(new_n1175), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n969), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1175), .B1(new_n1182), .B2(new_n882), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1196), .A2(new_n350), .A3(new_n352), .A4(new_n959), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1197), .A2(new_n957), .B1(new_n942), .B2(new_n964), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n952), .B1(new_n1198), .B2(KEYINPUT38), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1195), .A2(new_n1192), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1194), .A2(new_n1179), .A3(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1171), .B(KEYINPUT115), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n967), .A2(new_n968), .B1(new_n1192), .B2(new_n1191), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1195), .A2(new_n1192), .A3(new_n1199), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1186), .A2(new_n1189), .A3(new_n1201), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1176), .A2(new_n1177), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1207), .B1(new_n1208), .B2(new_n1188), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n747), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT120), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1201), .A2(new_n1205), .A3(new_n804), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT116), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1201), .A2(new_n1205), .A3(KEYINPUT116), .A4(new_n804), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n868), .B1(new_n967), .B2(new_n968), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n897), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G283), .A2(new_n839), .B1(new_n837), .B2(G107), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n909), .C1(new_n573), .C2(new_n830), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n857), .A2(G116), .B1(G77), .B2(new_n834), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT119), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(G97), .C2(new_n827), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n816), .A2(new_n314), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT118), .Z(new_n1225));
  NOR2_X1   g1025(.A1(new_n814), .A2(new_n375), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT53), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n843), .A2(G50), .B1(new_n849), .B2(G125), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n306), .B2(new_n835), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n314), .B1(new_n837), .B2(G137), .ZN(new_n1230));
  INV_X1    g1030(.A(G132), .ZN(new_n1231));
  INV_X1    g1031(.A(G128), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1230), .B1(new_n822), .B2(new_n1231), .C1(new_n1232), .C2(new_n840), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(KEYINPUT54), .B(G143), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT117), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1229), .B(new_n1233), .C1(new_n827), .C2(new_n1235), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1223), .A2(new_n1225), .B1(new_n1227), .B2(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n805), .B1(new_n341), .B2(new_n1218), .C1(new_n1237), .C2(new_n809), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1217), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1211), .B1(new_n1216), .B2(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(KEYINPUT120), .B(new_n1239), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1210), .B1(new_n1241), .B2(new_n1242), .ZN(G378));
  AND2_X1   g1043(.A1(new_n954), .A2(new_n970), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n990), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n738), .B1(new_n1245), .B2(new_n1199), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n383), .A2(new_n717), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n391), .A2(new_n393), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1250), .B1(new_n391), .B2(new_n393), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1248), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1253), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1251), .A3(new_n1247), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n982), .A2(new_n1246), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n982), .B2(new_n1246), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1244), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT121), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1257), .ZN(new_n1262));
  OAI21_X1  g1062(.A(G330), .B1(new_n983), .B2(new_n990), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n980), .B1(new_n953), .B2(new_n976), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n982), .A2(new_n1246), .A3(new_n1257), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n971), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1260), .A2(new_n1261), .A3(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n971), .A4(KEYINPUT121), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n804), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n806), .B1(new_n240), .B2(new_n897), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n815), .A2(new_n1235), .B1(G137), .B2(new_n827), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n839), .A2(G125), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n838), .B2(new_n1231), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G150), .B2(new_n834), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1272), .B(new_n1275), .C1(new_n1232), .C2(new_n822), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(KEYINPUT59), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(KEYINPUT59), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n272), .B(new_n256), .C1(new_n842), .C2(new_n306), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(G124), .B2(new_n849), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n256), .B1(new_n838), .B2(new_n490), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(G116), .B2(new_n839), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n506), .A2(new_n827), .B1(new_n857), .B2(G107), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(new_n219), .C2(new_n814), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n843), .A2(G58), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n847), .B2(new_n830), .ZN(new_n1287));
  NOR4_X1   g1087(.A1(new_n1285), .A2(new_n862), .A3(new_n1016), .A4(new_n1287), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1288), .A2(KEYINPUT58), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(KEYINPUT58), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n256), .B1(new_n288), .B2(new_n272), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n240), .ZN(new_n1292));
  AND4_X1   g1092(.A1(new_n1281), .A2(new_n1289), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n1271), .B1(new_n809), .B2(new_n1293), .C1(new_n1262), .C2(new_n868), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1270), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1189), .B1(new_n1208), .B2(new_n1207), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT57), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1260), .B2(new_n1267), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n748), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1295), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(G375));
  NAND2_X1  g1103(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1208), .A2(new_n1188), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1095), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n922), .A2(new_n867), .ZN(new_n1307));
  OAI22_X1  g1107(.A1(new_n814), .A2(new_n306), .B1(new_n1232), .B2(new_n830), .ZN(new_n1308));
  XOR2_X1   g1108(.A(new_n1308), .B(KEYINPUT122), .Z(new_n1309));
  OAI22_X1  g1109(.A1(new_n1018), .A2(new_n822), .B1(new_n826), .B2(new_n375), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n288), .B1(new_n839), .B2(G132), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1311), .B(new_n1286), .C1(new_n240), .C2(new_n835), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n1310), .B(new_n1312), .C1(new_n837), .C2(new_n1235), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n815), .A2(G97), .B1(G283), .B2(new_n857), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n827), .A2(G107), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1314), .A2(new_n1123), .A3(new_n1315), .ZN(new_n1316));
  OAI22_X1  g1116(.A1(new_n443), .A2(new_n842), .B1(new_n830), .B2(new_n659), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n314), .B1(new_n840), .B2(new_n573), .ZN(new_n1318));
  AOI211_X1 g1118(.A(new_n1317), .B(new_n1318), .C1(G116), .C2(new_n837), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n1309), .A2(new_n1313), .B1(new_n1316), .B2(new_n1319), .ZN(new_n1320));
  OAI221_X1 g1120(.A(new_n805), .B1(G68), .B2(new_n1218), .C1(new_n1320), .C2(new_n809), .ZN(new_n1321));
  XOR2_X1   g1121(.A(new_n1321), .B(KEYINPUT123), .Z(new_n1322));
  AOI22_X1  g1122(.A1(new_n1186), .A2(new_n804), .B1(new_n1307), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1306), .A2(new_n1323), .ZN(G381));
  INV_X1    g1124(.A(G390), .ZN(new_n1325));
  INV_X1    g1125(.A(G384), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NOR4_X1   g1127(.A1(new_n1327), .A2(G396), .A3(G381), .A4(G393), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1033), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1061), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1073), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1097), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1099), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1075), .A2(KEYINPUT107), .A3(new_n1097), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1329), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1239), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1210), .A2(new_n1336), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1328), .A2(new_n1335), .A3(new_n1302), .A4(new_n1337), .ZN(G407));
  NAND3_X1  g1138(.A1(new_n720), .A2(new_n721), .A3(G213), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1302), .A2(new_n1337), .A3(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(G407), .A2(G213), .A3(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(KEYINPUT124), .ZN(G409));
  NAND2_X1  g1143(.A1(new_n1302), .A2(G378), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1260), .A2(new_n1267), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n804), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1294), .B(new_n1346), .C1(new_n1297), .C2(new_n1094), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1337), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1344), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1339), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1340), .A2(G2897), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1351), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1178), .A2(new_n1188), .A3(KEYINPUT60), .A4(new_n1185), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n747), .ZN(new_n1354));
  OAI21_X1  g1154(.A(KEYINPUT60), .B1(new_n1208), .B2(new_n1188), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1354), .B1(new_n1305), .B2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1323), .ZN(new_n1357));
  NOR3_X1   g1157(.A1(new_n1356), .A2(new_n1326), .A3(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1305), .ZN(new_n1359));
  AND2_X1   g1159(.A1(new_n1353), .A2(new_n747), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(G384), .B1(new_n1361), .B2(new_n1323), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1352), .B1(new_n1358), .B2(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1326), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1361), .A2(G384), .A3(new_n1323), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1364), .A2(new_n1365), .A3(new_n1351), .ZN(new_n1366));
  AND2_X1   g1166(.A1(new_n1363), .A2(new_n1366), .ZN(new_n1367));
  AOI21_X1  g1167(.A(KEYINPUT61), .B1(new_n1350), .B2(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1340), .B1(new_n1344), .B2(new_n1348), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1364), .A2(new_n1365), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1369), .A2(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT63), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT125), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(G387), .A2(new_n1325), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1335), .A2(G390), .ZN(new_n1377));
  XNOR2_X1  g1177(.A(G393), .B(new_n878), .ZN(new_n1378));
  AND4_X1   g1178(.A1(new_n1375), .A2(new_n1376), .A3(new_n1377), .A4(new_n1378), .ZN(new_n1379));
  OAI21_X1  g1179(.A(KEYINPUT125), .B1(new_n1335), .B2(G390), .ZN(new_n1380));
  AOI22_X1  g1180(.A1(new_n1380), .A2(new_n1378), .B1(new_n1376), .B2(new_n1377), .ZN(new_n1381));
  NOR2_X1   g1181(.A1(new_n1379), .A2(new_n1381), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1369), .A2(KEYINPUT63), .A3(new_n1371), .ZN(new_n1383));
  NAND4_X1  g1183(.A1(new_n1368), .A2(new_n1374), .A3(new_n1382), .A4(new_n1383), .ZN(new_n1384));
  INV_X1    g1184(.A(KEYINPUT61), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1363), .A2(new_n1366), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1385), .B1(new_n1369), .B2(new_n1386), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1388), .B1(new_n1369), .B2(new_n1371), .ZN(new_n1389));
  AOI22_X1  g1189(.A1(new_n1302), .A2(G378), .B1(new_n1347), .B2(new_n1337), .ZN(new_n1390));
  XNOR2_X1  g1190(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1391));
  NOR4_X1   g1191(.A1(new_n1390), .A2(new_n1340), .A3(new_n1370), .A4(new_n1391), .ZN(new_n1392));
  NOR3_X1   g1192(.A1(new_n1387), .A2(new_n1389), .A3(new_n1392), .ZN(new_n1393));
  OAI21_X1  g1193(.A(new_n1384), .B1(new_n1393), .B2(new_n1382), .ZN(G405));
  NAND2_X1  g1194(.A1(G375), .A2(new_n1337), .ZN(new_n1395));
  AND2_X1   g1195(.A1(new_n1395), .A2(new_n1344), .ZN(new_n1396));
  OR2_X1    g1196(.A1(new_n1370), .A2(KEYINPUT127), .ZN(new_n1397));
  AND2_X1   g1197(.A1(new_n1396), .A2(new_n1397), .ZN(new_n1398));
  NOR2_X1   g1198(.A1(new_n1396), .A2(new_n1397), .ZN(new_n1399));
  OAI22_X1  g1199(.A1(new_n1398), .A2(new_n1399), .B1(new_n1379), .B2(new_n1381), .ZN(new_n1400));
  OR2_X1    g1200(.A1(new_n1396), .A2(new_n1397), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1396), .A2(new_n1397), .ZN(new_n1402));
  NAND3_X1  g1202(.A1(new_n1401), .A2(new_n1382), .A3(new_n1402), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(new_n1400), .A2(new_n1403), .ZN(G402));
endmodule


