//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g0008(.A(G250), .B1(G257), .B2(G264), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n210), .A2(KEYINPUT0), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT64), .Z(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n216), .B(new_n224), .C1(KEYINPUT0), .C2(new_n210), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT65), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G68), .B(G77), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(G50), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G97), .B(G107), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  XOR2_X1   g0042(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G68), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT7), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  AND2_X1   g0047(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n248));
  NOR2_X1   g0048(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n248), .A2(new_n249), .A3(G33), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n247), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n246), .B1(new_n255), .B2(G20), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n245), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G58), .A2(G68), .ZN(new_n258));
  OAI21_X1  g0058(.A(G20), .B1(new_n258), .B2(new_n201), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT77), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(KEYINPUT77), .B(G20), .C1(new_n258), .C2(new_n201), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G159), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n244), .B1(new_n257), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT76), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n251), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n246), .B(new_n212), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G68), .ZN(new_n276));
  OAI21_X1  g0076(.A(G33), .B1(new_n248), .B2(new_n249), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n273), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n246), .B1(new_n278), .B2(new_n212), .ZN(new_n279));
  OAI211_X1 g0079(.A(KEYINPUT16), .B(new_n267), .C1(new_n276), .C2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT69), .B1(new_n206), .B2(new_n268), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT69), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n282), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(new_n211), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n266), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n284), .B1(new_n288), .B2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n291), .B1(new_n293), .B2(new_n287), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n285), .A2(KEYINPUT79), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(KEYINPUT79), .B1(new_n285), .B2(new_n295), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  NAND3_X1  g0098(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT68), .B1(G33), .B2(G41), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n300), .A2(new_n301), .A3(new_n211), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  AOI21_X1  g0105(.A(G1), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT67), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n288), .B1(G41), .B2(G45), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n308), .A2(G274), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n302), .A2(new_n306), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n303), .A2(new_n311), .B1(new_n312), .B2(G232), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(G226), .A2(G1698), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n277), .A2(new_n273), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT80), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G87), .ZN(new_n320));
  INV_X1    g0120(.A(G1698), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n277), .A2(G223), .A3(new_n321), .A4(new_n273), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT80), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n277), .A2(new_n323), .A3(new_n273), .A4(new_n317), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n319), .A2(new_n320), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n316), .B1(new_n325), .B2(KEYINPUT81), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n322), .A2(new_n320), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT81), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n319), .A4(new_n324), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n298), .B(new_n314), .C1(new_n326), .C2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n325), .A2(KEYINPUT81), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n329), .A3(new_n315), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(new_n313), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n296), .A2(new_n297), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT18), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n285), .A2(new_n295), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT79), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n285), .A2(KEYINPUT79), .A3(new_n295), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n333), .A2(new_n313), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G169), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n314), .B1(new_n326), .B2(new_n329), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n341), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n336), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n342), .A2(G200), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n333), .A2(G190), .A3(new_n313), .ZN(new_n351));
  INV_X1    g0151(.A(new_n284), .ZN(new_n352));
  AOI21_X1  g0152(.A(G20), .B1(new_n277), .B2(new_n273), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n245), .B1(new_n353), .B2(new_n246), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n270), .A2(new_n271), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n274), .B1(new_n355), .B2(G33), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT7), .B1(new_n356), .B2(G20), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n265), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n352), .B1(new_n358), .B2(KEYINPUT16), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n294), .B1(new_n359), .B2(new_n266), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n350), .A2(KEYINPUT83), .A3(new_n351), .A4(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT82), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT17), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n360), .B(new_n351), .C1(new_n364), .C2(new_n344), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n362), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT17), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n349), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n352), .B(KEYINPUT71), .C1(G1), .C2(new_n212), .ZN(new_n370));
  INV_X1    g0170(.A(G77), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT72), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT72), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n292), .A2(KEYINPUT71), .A3(new_n373), .A4(G77), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n287), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT70), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n378), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n268), .A2(G20), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n376), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n289), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n288), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n384), .A2(new_n284), .B1(new_n371), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n375), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n255), .A2(G1698), .ZN(new_n391));
  INV_X1    g0191(.A(G238), .ZN(new_n392));
  INV_X1    g0192(.A(G107), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n391), .A2(new_n392), .B1(new_n393), .B2(new_n255), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n255), .A2(G232), .A3(new_n321), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n315), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n311), .A2(new_n303), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n312), .A2(G244), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n331), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n390), .B(new_n400), .C1(G179), .C2(new_n399), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(G200), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n396), .A2(G190), .A3(new_n397), .A4(new_n398), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n402), .A2(new_n375), .A3(new_n389), .A4(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n312), .A2(G226), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n397), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n255), .A2(G222), .A3(new_n321), .ZN(new_n408));
  INV_X1    g0208(.A(G223), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n408), .B1(new_n371), .B2(new_n255), .C1(new_n391), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n315), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n331), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n203), .A2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(G150), .ZN(new_n415));
  INV_X1    g0215(.A(new_n263), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n414), .B1(new_n415), .B2(new_n416), .C1(new_n286), .C2(new_n383), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n284), .B1(new_n202), .B2(new_n290), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n292), .A2(G50), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n413), .B(new_n420), .C1(G179), .C2(new_n412), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n364), .B1(new_n407), .B2(new_n411), .ZN(new_n422));
  INV_X1    g0222(.A(new_n412), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n422), .B1(G190), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT10), .ZN(new_n425));
  NAND2_X1  g0225(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT73), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT9), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n420), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n418), .A2(new_n427), .A3(new_n428), .A4(new_n419), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n424), .A2(new_n425), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n425), .B1(new_n424), .B2(new_n432), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n405), .B(new_n421), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT74), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n416), .B2(new_n202), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n382), .A2(G77), .B1(G20), .B2(new_n245), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n263), .A2(KEYINPUT74), .A3(G50), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n284), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT11), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n370), .A2(KEYINPUT12), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G68), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT12), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G68), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n388), .A2(new_n446), .B1(new_n445), .B2(new_n289), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n442), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n312), .A2(G238), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n397), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n255), .A2(G232), .A3(G1698), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n255), .A2(G226), .A3(new_n321), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G97), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n315), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT13), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n303), .A2(new_n311), .B1(new_n312), .B2(G238), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT13), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n456), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(G179), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT75), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT14), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n458), .A2(new_n461), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(G169), .ZN(new_n467));
  AOI211_X1 g0267(.A(KEYINPUT14), .B(new_n331), .C1(new_n458), .C2(new_n461), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n449), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G190), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n449), .B1(new_n471), .B2(new_n466), .ZN(new_n472));
  INV_X1    g0272(.A(new_n461), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n460), .B1(new_n459), .B2(new_n456), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n364), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n435), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n369), .A2(KEYINPUT84), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT84), .B1(new_n369), .B2(new_n478), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n277), .A2(G238), .A3(new_n321), .A4(new_n273), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n277), .A2(G244), .A3(G1698), .A4(new_n273), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G116), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n315), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n288), .A2(G45), .A3(G274), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(G250), .B1(new_n305), .B2(G1), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n302), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT87), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT87), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n494), .B(new_n491), .C1(new_n486), .C2(new_n315), .ZN(new_n495));
  OAI21_X1  g0295(.A(G190), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT88), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n493), .A2(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G200), .ZN(new_n500));
  OAI211_X1 g0300(.A(KEYINPUT88), .B(G190), .C1(new_n493), .C2(new_n495), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT19), .B1(new_n382), .B2(G97), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT19), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n212), .B1(new_n454), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G87), .ZN(new_n505));
  INV_X1    g0305(.A(G97), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(new_n393), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n502), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n212), .A2(G68), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n278), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n284), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n381), .A2(new_n388), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n288), .A2(G33), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n352), .A2(new_n289), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(G87), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n498), .A2(new_n500), .A3(new_n501), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n499), .A2(new_n331), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n511), .B(new_n512), .C1(new_n381), .C2(new_n515), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n520), .C1(G179), .C2(new_n499), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n515), .A2(new_n393), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n290), .A2(new_n393), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT25), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT24), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(new_n505), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n277), .A2(new_n273), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n485), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n212), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n273), .A2(new_n252), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n212), .A2(G87), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n528), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n393), .A3(G20), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT89), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n536), .A2(new_n393), .A3(KEYINPUT89), .A4(G20), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT23), .B1(new_n212), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n535), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n527), .B1(new_n532), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(G20), .B1(new_n530), .B2(new_n485), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n546), .A2(new_n543), .A3(KEYINPUT24), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n284), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(KEYINPUT90), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT90), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n532), .A2(new_n544), .A3(new_n527), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT24), .B1(new_n546), .B2(new_n543), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n553), .B2(new_n284), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n526), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(G250), .A2(G1698), .ZN(new_n556));
  INV_X1    g0356(.A(G257), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(G1698), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(new_n277), .A3(new_n273), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G294), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n301), .A2(new_n211), .ZN(new_n562));
  XNOR2_X1  g0362(.A(KEYINPUT5), .B(G41), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n305), .A2(G1), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n299), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n561), .A2(new_n315), .B1(G264), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n488), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT86), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT86), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n563), .A2(new_n488), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT91), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(G179), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n566), .A2(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G169), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT91), .B1(new_n575), .B2(new_n298), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n555), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  INV_X1    g0380(.A(G116), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n388), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n352), .A2(new_n514), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n386), .A2(G116), .A3(new_n387), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT85), .ZN(new_n586));
  INV_X1    g0386(.A(G283), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n268), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(KEYINPUT85), .A2(G33), .A3(G283), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(G20), .B1(new_n268), .B2(G97), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(G20), .B2(new_n581), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT20), .B1(new_n592), .B2(new_n284), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n284), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n585), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n565), .A2(G270), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n571), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n557), .A2(new_n321), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n321), .A2(G264), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n277), .A2(new_n273), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n533), .A2(G303), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n316), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(G169), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n580), .B1(new_n596), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n284), .B1(new_n288), .B2(G33), .ZN(new_n606));
  INV_X1    g0406(.A(new_n584), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n595), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n582), .B(new_n608), .C1(new_n609), .C2(new_n593), .ZN(new_n610));
  INV_X1    g0410(.A(new_n603), .ZN(new_n611));
  AOI22_X1  g0411(.A1(G270), .A2(new_n565), .B1(new_n568), .B2(new_n570), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n610), .A2(new_n613), .A3(KEYINPUT21), .A4(G169), .ZN(new_n614));
  OAI21_X1  g0414(.A(G200), .B1(new_n598), .B2(new_n603), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n611), .A2(new_n612), .A3(G190), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n596), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n613), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n610), .A2(new_n618), .A3(G179), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n605), .A2(new_n614), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT6), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n240), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n393), .A2(KEYINPUT6), .A3(G97), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n625));
  INV_X1    g0425(.A(new_n247), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n270), .A2(new_n268), .A3(new_n271), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n252), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT7), .B1(new_n533), .B2(new_n212), .ZN(new_n629));
  OAI21_X1  g0429(.A(G107), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n352), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n290), .A2(new_n506), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n515), .B2(new_n506), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n277), .A2(G244), .A3(new_n321), .A4(new_n273), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT4), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(KEYINPUT4), .A2(G244), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n273), .A2(new_n252), .A3(new_n638), .A4(new_n321), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n273), .A2(new_n252), .A3(G250), .A4(G1698), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n590), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n316), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n565), .A2(G257), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n571), .ZN(new_n644));
  OAI21_X1  g0444(.A(G169), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AOI22_X1  g0445(.A1(G257), .A2(new_n565), .B1(new_n568), .B2(new_n570), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n639), .A2(new_n590), .A3(new_n640), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n636), .B2(new_n635), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n646), .B(G179), .C1(new_n648), .C2(new_n316), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n634), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n646), .B1(new_n648), .B2(new_n316), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G200), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n631), .A2(new_n633), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n646), .B(G190), .C1(new_n648), .C2(new_n316), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n620), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n364), .B1(new_n566), .B2(new_n571), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(G190), .B2(new_n572), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n526), .B(new_n660), .C1(new_n549), .C2(new_n554), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n579), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n482), .A2(new_n522), .A3(new_n662), .ZN(G372));
  AND3_X1   g0463(.A1(new_n605), .A2(new_n614), .A3(new_n619), .ZN(new_n664));
  INV_X1    g0464(.A(new_n526), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n548), .A2(KEYINPUT90), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n553), .A2(new_n550), .A3(new_n284), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n657), .B1(new_n668), .B2(new_n660), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n487), .A2(new_n492), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n331), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n520), .B(new_n673), .C1(new_n499), .C2(G179), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(G200), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n498), .A2(new_n501), .A3(new_n517), .A4(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n670), .A2(new_n671), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n651), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n518), .A2(new_n521), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n650), .A2(KEYINPUT92), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT92), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n645), .B2(new_n649), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n681), .A2(new_n654), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n676), .A2(new_n684), .A3(new_n685), .A4(new_n674), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n677), .A2(new_n680), .A3(new_n674), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n481), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n433), .A2(new_n434), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n361), .A2(new_n362), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT17), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n366), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n368), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n462), .B(KEYINPUT75), .ZN(new_n695));
  OAI21_X1  g0495(.A(G169), .B1(new_n473), .B2(new_n474), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT14), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n466), .A2(new_n465), .A3(G169), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n448), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n477), .B2(new_n401), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n337), .B1(new_n330), .B2(new_n334), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT18), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n689), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n705), .A2(new_n421), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n688), .A2(new_n706), .ZN(G369));
  OAI21_X1  g0507(.A(new_n661), .B1(new_n668), .B2(new_n669), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n212), .A2(G13), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n288), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G343), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n668), .A2(new_n716), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n708), .A2(new_n717), .B1(new_n579), .B2(new_n716), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n664), .A2(new_n715), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n664), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n596), .A2(new_n716), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n620), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n708), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n719), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n555), .A2(new_n578), .A3(new_n716), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n727), .A2(new_n732), .ZN(G399));
  NOR2_X1   g0533(.A1(new_n208), .A2(G41), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n507), .A2(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G1), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n215), .B2(new_n735), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n687), .A2(new_n716), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n676), .A2(new_n684), .A3(new_n674), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(KEYINPUT26), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n518), .A2(new_n521), .A3(new_n685), .A4(new_n678), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n674), .B(KEYINPUT95), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n677), .A2(new_n743), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n716), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT29), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n561), .A2(new_n315), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n565), .A2(G264), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT93), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n613), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n649), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n756), .A2(new_n499), .B1(KEYINPUT93), .B2(new_n751), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n493), .A2(new_n495), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n751), .A2(KEYINPUT93), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n758), .A2(new_n755), .A3(new_n759), .A4(new_n754), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n618), .A2(G179), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n761), .A2(new_n575), .A3(new_n652), .A4(new_n672), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n757), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n715), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT94), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n715), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT31), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n766), .A2(KEYINPUT94), .A3(new_n767), .ZN(new_n770));
  INV_X1    g0570(.A(new_n522), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n728), .A2(new_n771), .A3(new_n658), .A4(new_n716), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G330), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n741), .A2(new_n748), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n739), .B1(new_n776), .B2(G1), .ZN(G364));
  AOI21_X1  g0577(.A(new_n288), .B1(new_n709), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n734), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n726), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G330), .B2(new_n724), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n211), .B1(G20), .B2(new_n331), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n298), .A2(new_n364), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n212), .A2(G190), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G317), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT33), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(KEYINPUT33), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n212), .A2(new_n471), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n298), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT97), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n795), .A2(new_n796), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n792), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT100), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n793), .A2(new_n785), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n794), .A2(new_n786), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n806), .A2(G326), .B1(new_n808), .B2(G311), .ZN(new_n809));
  INV_X1    g0609(.A(G303), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n793), .A2(new_n298), .A3(G200), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n809), .B(new_n533), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n298), .A2(new_n364), .A3(G190), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(G294), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n786), .B(KEYINPUT99), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n816), .A2(G179), .A3(new_n364), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n816), .A2(G179), .A3(G200), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G283), .A2(new_n817), .B1(new_n818), .B2(G329), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n804), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(G159), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT32), .Z(new_n822));
  INV_X1    g0622(.A(new_n814), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n255), .B1(new_n807), .B2(new_n371), .C1(new_n823), .C2(new_n506), .ZN(new_n824));
  INV_X1    g0624(.A(new_n811), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n825), .A2(G87), .B1(new_n788), .B2(G68), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n202), .B2(new_n805), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n824), .B(new_n827), .C1(G107), .C2(new_n817), .ZN(new_n828));
  INV_X1    g0628(.A(G58), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n800), .B(KEYINPUT98), .Z(new_n830));
  OAI211_X1 g0630(.A(new_n822), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n784), .B1(new_n820), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(G13), .A2(G33), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(G20), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n783), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n238), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n356), .A2(new_n208), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(G45), .B2(new_n215), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n838), .A2(G45), .B1(KEYINPUT96), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(KEYINPUT96), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n208), .A2(new_n533), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n843), .A2(G355), .B1(new_n581), .B2(new_n208), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n837), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n780), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n832), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n835), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n724), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n782), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  NAND2_X1  g0651(.A1(new_n390), .A2(new_n715), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n404), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n401), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n401), .A2(new_n715), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n740), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n687), .A2(new_n716), .A3(new_n857), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n780), .B1(new_n861), .B2(new_n774), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n774), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n857), .A2(new_n834), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n783), .A2(new_n833), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n817), .A2(G87), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n805), .A2(new_n810), .B1(new_n807), .B2(new_n581), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(G283), .B2(new_n788), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT101), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n533), .B1(new_n811), .B2(new_n393), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G97), .B2(new_n814), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n800), .A2(G294), .B1(new_n818), .B2(G311), .ZN(new_n873));
  AND4_X1   g0673(.A1(new_n867), .A2(new_n870), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n806), .A2(G137), .B1(new_n808), .B2(G159), .ZN(new_n875));
  INV_X1    g0675(.A(G143), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n875), .B1(new_n415), .B2(new_n787), .C1(new_n830), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT34), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n356), .B1(new_n811), .B2(new_n202), .C1(new_n823), .C2(new_n829), .ZN(new_n879));
  INV_X1    g0679(.A(new_n817), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n245), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n879), .B(new_n881), .C1(G132), .C2(new_n818), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n874), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n780), .B1(G77), .B2(new_n866), .C1(new_n883), .C2(new_n784), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT102), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n863), .B1(new_n864), .B2(new_n885), .ZN(G384));
  OAI211_X1 g0686(.A(G116), .B(new_n213), .C1(new_n624), .C2(KEYINPUT35), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(KEYINPUT35), .B2(new_n624), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT36), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n215), .A2(new_n258), .A3(new_n371), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n202), .B2(G68), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n288), .B(G13), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(G330), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n772), .A2(new_n768), .A3(new_n764), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  INV_X1    g0698(.A(new_n477), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n448), .A2(new_n715), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n700), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n470), .A2(new_n715), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n897), .A2(new_n898), .A3(new_n857), .A4(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n358), .A2(new_n243), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n280), .A2(new_n284), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n295), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n713), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n360), .A2(new_n351), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n344), .A2(new_n364), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n906), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n294), .B1(new_n914), .B2(new_n359), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n343), .B2(new_n345), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT105), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n337), .B1(G190), .B2(new_n344), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n341), .A2(new_n909), .B1(new_n920), .B2(new_n350), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n335), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT37), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n341), .A2(new_n346), .A3(KEYINPUT106), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n921), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT105), .B(KEYINPUT37), .C1(new_n913), .C2(new_n916), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n919), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n349), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n910), .B1(new_n694), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n905), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n919), .A2(new_n926), .A3(new_n927), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(KEYINPUT38), .C1(new_n369), .C2(new_n910), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n904), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n662), .A2(new_n522), .A3(new_n715), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n768), .A2(new_n764), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n903), .B(new_n857), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n933), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n909), .B1(new_n296), .B2(new_n297), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT17), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n942), .A2(new_n363), .A3(new_n366), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n941), .B1(new_n943), .B2(new_n704), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n703), .A3(new_n365), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT37), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT107), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n948), .A3(KEYINPUT37), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n926), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT38), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n938), .B1(new_n939), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n934), .B1(new_n952), .B2(KEYINPUT40), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n481), .A2(new_n897), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n896), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(new_n910), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n943), .B2(new_n349), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT38), .B1(new_n958), .B2(new_n932), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT39), .B1(new_n939), .B2(new_n959), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n947), .A2(new_n926), .A3(new_n949), .ZN(new_n961));
  INV_X1    g0761(.A(new_n704), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n940), .B1(new_n694), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n905), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT39), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(new_n965), .A3(new_n933), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n700), .A2(new_n715), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n856), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n860), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n903), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT104), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n972), .A2(new_n973), .B1(new_n933), .B2(new_n931), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(KEYINPUT104), .A3(new_n903), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n704), .A2(new_n713), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n969), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n956), .B(new_n978), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n705), .A2(new_n421), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n741), .A2(new_n748), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(new_n481), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n288), .B2(new_n709), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n979), .A2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n895), .B1(new_n984), .B2(new_n985), .ZN(G367));
  INV_X1    g0786(.A(new_n657), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n728), .A2(new_n987), .A3(new_n719), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT42), .Z(new_n989));
  OAI21_X1  g0789(.A(new_n987), .B1(new_n654), .B2(new_n716), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n684), .A2(new_n715), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n651), .B1(new_n993), .B2(new_n579), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n716), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n676), .B(new_n674), .C1(new_n517), .C2(new_n716), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n674), .A2(new_n517), .A3(new_n716), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n989), .A2(new_n995), .B1(KEYINPUT43), .B2(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n727), .A2(new_n993), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n734), .B(KEYINPUT41), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n720), .A2(new_n726), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n727), .A3(new_n729), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n731), .A2(new_n993), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT44), .Z(new_n1012));
  OR3_X1    g0812(.A1(new_n731), .A2(KEYINPUT108), .A3(new_n993), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT108), .B1(new_n731), .B2(new_n993), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT45), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1017));
  OAI211_X1 g0817(.A(KEYINPUT109), .B(new_n1010), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1007), .B1(new_n1018), .B2(new_n776), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1005), .B1(new_n1019), .B2(new_n779), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n839), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n836), .B1(new_n207), .B2(new_n381), .C1(new_n1021), .C2(new_n233), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n846), .B1(new_n1022), .B2(KEYINPUT110), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(KEYINPUT110), .B2(new_n1022), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n805), .A2(new_n876), .B1(new_n807), .B2(new_n202), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n814), .A2(G68), .ZN(new_n1026));
  INV_X1    g0826(.A(G159), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n255), .C1(new_n1027), .C2(new_n787), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1025), .B(new_n1028), .C1(G58), .C2(new_n825), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n800), .A2(G150), .B1(new_n817), .B2(G77), .ZN(new_n1030));
  INV_X1    g0830(.A(G137), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n818), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1029), .B(new_n1030), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(G311), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n830), .A2(new_n810), .B1(new_n1034), .B2(new_n805), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT111), .Z(new_n1036));
  NAND2_X1  g0836(.A1(new_n817), .A2(G97), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n818), .A2(G317), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G294), .A2(new_n788), .B1(new_n808), .B2(G283), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n278), .A4(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n825), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT46), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n811), .B2(new_n581), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(new_n393), .C2(new_n823), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1033), .B1(new_n1036), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT47), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n784), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1024), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n998), .B2(new_n848), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1020), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1052), .A2(KEYINPUT112), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT112), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1020), .B2(new_n1051), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(G387));
  NAND2_X1  g0857(.A1(new_n776), .A2(new_n1010), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n734), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1059), .A2(KEYINPUT113), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(KEYINPUT113), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n775), .A2(new_n1009), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT114), .Z(new_n1063));
  NAND3_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n839), .B1(new_n230), .B2(new_n305), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n843), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n736), .B2(new_n1066), .ZN(new_n1067));
  OR3_X1    g0867(.A1(new_n286), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1068));
  OAI21_X1  g0868(.A(KEYINPUT50), .B1(new_n286), .B2(G50), .ZN(new_n1069));
  AOI21_X1  g0869(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1068), .A2(new_n736), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1067), .A2(new_n1071), .B1(new_n393), .B2(new_n208), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n780), .B1(new_n1072), .B2(new_n837), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n800), .A2(G50), .B1(new_n818), .B2(G150), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n811), .A2(new_n371), .B1(new_n787), .B2(new_n286), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n805), .A2(new_n1027), .B1(new_n807), .B2(new_n245), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1075), .A2(new_n1076), .A3(new_n278), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n379), .A2(new_n380), .A3(new_n814), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1074), .A2(new_n1037), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n356), .B1(new_n818), .B2(G326), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n806), .A2(G322), .B1(new_n808), .B2(G303), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n1034), .B2(new_n787), .C1(new_n830), .C2(new_n789), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT48), .Z(new_n1083));
  INV_X1    g0883(.A(G294), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n823), .A2(new_n587), .B1(new_n811), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1080), .B1(new_n581), .B2(new_n880), .C1(new_n1086), .C2(KEYINPUT49), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1086), .A2(KEYINPUT49), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1079), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1073), .B1(new_n1089), .B2(new_n783), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n718), .A2(new_n848), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1090), .A2(new_n1091), .B1(new_n779), .B2(new_n1010), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1064), .A2(new_n1092), .ZN(G393));
  NAND2_X1  g0893(.A1(new_n839), .A2(new_n241), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1094), .B(new_n836), .C1(new_n506), .C2(new_n207), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT115), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n846), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n801), .A2(new_n1034), .B1(new_n789), .B2(new_n805), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT52), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n533), .B1(new_n787), .B2(new_n810), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n811), .A2(new_n587), .B1(new_n807), .B2(new_n1084), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(G116), .C2(new_n814), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G107), .A2(new_n817), .B1(new_n818), .B2(G322), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n800), .A2(G159), .B1(G150), .B2(new_n806), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT51), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n818), .A2(G143), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n811), .A2(new_n245), .B1(new_n787), .B2(new_n202), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n287), .B2(new_n808), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n278), .B1(G77), .B2(new_n814), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n867), .A2(new_n1110), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1106), .A2(new_n1107), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1098), .B1(new_n1115), .B2(new_n783), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n992), .B2(new_n848), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT109), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n726), .B(new_n720), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(KEYINPUT109), .B(new_n727), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n734), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1117), .B1(new_n1122), .B2(new_n1058), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1118), .B(new_n727), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n778), .B2(new_n1059), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(G390));
  NAND2_X1  g0927(.A1(new_n938), .A2(G330), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n964), .A2(new_n965), .A3(new_n933), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n965), .B1(new_n931), .B2(new_n933), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n968), .B1(new_n971), .B2(new_n903), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n964), .A2(new_n933), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n968), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n746), .A2(new_n716), .A3(new_n854), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n970), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n903), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1129), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n773), .A2(G330), .A3(new_n857), .A4(new_n903), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1142), .B(new_n1139), .C1(new_n967), .C2(new_n1132), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n779), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n881), .B1(G116), .B2(new_n800), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n1084), .B2(new_n1032), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n806), .A2(G283), .B1(new_n808), .B2(G97), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n393), .B2(new_n787), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n533), .B1(new_n811), .B2(new_n505), .C1(new_n823), .C2(new_n371), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(G132), .ZN(new_n1151));
  INV_X1    g0951(.A(G125), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n801), .A2(new_n1151), .B1(new_n1032), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n533), .B1(new_n806), .B2(G128), .ZN(new_n1154));
  XOR2_X1   g0954(.A(KEYINPUT54), .B(G143), .Z(new_n1155));
  AOI22_X1  g0955(.A1(new_n788), .A2(G137), .B1(new_n808), .B2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(new_n880), .C2(new_n202), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n825), .B2(G150), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n825), .A2(new_n1158), .A3(G150), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1027), .B2(new_n823), .ZN(new_n1161));
  NOR4_X1   g0961(.A1(new_n1153), .A2(new_n1157), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n783), .B1(new_n1150), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n846), .B1(new_n286), .B2(new_n865), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n967), .C2(new_n834), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1144), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n747), .A2(KEYINPUT29), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1168), .A2(new_n1169), .B1(new_n479), .B2(new_n480), .ZN(new_n1170));
  OAI211_X1 g0970(.A(G330), .B(new_n897), .C1(new_n479), .C2(new_n480), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n706), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n903), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n774), .B2(new_n858), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1128), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n971), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n897), .A2(G330), .A3(new_n857), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1173), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1178), .A2(new_n970), .A3(new_n1142), .A4(new_n1136), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1172), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n735), .B1(new_n1167), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1141), .A2(new_n1143), .A3(new_n1180), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1166), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(G378));
  NAND2_X1  g0985(.A1(new_n689), .A2(new_n421), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n420), .A2(new_n909), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1188), .B(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n953), .A2(new_n896), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n904), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n939), .B2(new_n959), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n937), .B1(new_n964), .B2(new_n933), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n898), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1190), .B1(new_n1196), .B2(G330), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n978), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1191), .B1(new_n953), .B2(new_n896), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(G330), .A3(new_n1190), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n967), .A2(new_n968), .B1(new_n704), .B2(new_n713), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1199), .A2(new_n976), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1191), .A2(new_n833), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n780), .B1(new_n866), .B2(G50), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1026), .B1(new_n506), .B2(new_n787), .C1(new_n581), .C2(new_n805), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1032), .A2(new_n587), .B1(new_n381), .B2(new_n807), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G58), .C2(new_n817), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n278), .B(new_n304), .C1(new_n371), .C2(new_n811), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT118), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n800), .A2(G107), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT119), .Z(new_n1212));
  NAND3_X1  g1012(.A1(new_n1208), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT58), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n268), .A2(new_n304), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT117), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1216), .B(new_n202), .C1(new_n356), .C2(G41), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n807), .A2(new_n1031), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n825), .B2(new_n1155), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G125), .A2(new_n806), .B1(new_n788), .B2(G132), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n415), .C2(new_n823), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G128), .B2(new_n800), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT59), .Z(new_n1223));
  AOI21_X1  g1023(.A(new_n1216), .B1(new_n817), .B2(G159), .ZN(new_n1224));
  INV_X1    g1024(.A(G124), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n1032), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT120), .Z(new_n1227));
  OAI211_X1 g1027(.A(new_n1214), .B(new_n1217), .C1(new_n1223), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1205), .B1(new_n1228), .B2(new_n783), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1203), .A2(new_n779), .B1(new_n1204), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT121), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1172), .B(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1183), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1203), .A2(new_n1233), .A3(KEYINPUT57), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n734), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1233), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1230), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT122), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT122), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1239), .B(new_n1230), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(G375));
  NAND2_X1  g1041(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1172), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(new_n1006), .A3(new_n1181), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n779), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n846), .B1(new_n245), .B2(new_n865), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n788), .A2(new_n1155), .B1(new_n808), .B2(G150), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1248), .B1(new_n1151), .B2(new_n805), .C1(new_n1027), .C2(new_n811), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n278), .B(new_n1249), .C1(G50), .C2(new_n814), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G58), .A2(new_n817), .B1(new_n818), .B2(G128), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(new_n1031), .C2(new_n830), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n800), .A2(G283), .B1(new_n818), .B2(G303), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n533), .B1(new_n807), .B2(new_n393), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n811), .A2(new_n506), .B1(new_n805), .B2(new_n1084), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(G116), .C2(new_n788), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n817), .A2(G77), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1253), .A2(new_n1256), .A3(new_n1257), .A4(new_n1078), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1252), .A2(new_n1258), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1247), .B1(new_n784), .B2(new_n1259), .C1(new_n903), .C2(new_n834), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1245), .A2(new_n1246), .A3(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT123), .ZN(G381));
  OR2_X1    g1062(.A1(G390), .A2(G384), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1064), .A2(new_n850), .A3(new_n1092), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(G387), .A2(new_n1263), .A3(G381), .A4(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1238), .A2(new_n1184), .A3(new_n1240), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(G407));
  NAND2_X1  g1068(.A1(new_n714), .A2(G213), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT124), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G407), .B(G213), .C1(new_n1266), .C2(new_n1271), .ZN(G409));
  NAND3_X1  g1072(.A1(new_n1203), .A2(new_n1233), .A3(new_n1006), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1230), .A2(new_n1184), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1203), .A2(new_n779), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1204), .A2(new_n1229), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1202), .A2(new_n1198), .B1(new_n1183), .B2(new_n1232), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n735), .B1(new_n1278), .B2(KEYINPUT57), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1236), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1277), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1271), .B(new_n1274), .C1(new_n1281), .C2(new_n1184), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1243), .A2(KEYINPUT60), .A3(new_n1172), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT60), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1172), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1285), .B1(new_n1242), .B2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1284), .A2(new_n1287), .A3(new_n734), .A4(new_n1181), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1246), .A2(new_n1260), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1283), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1288), .A2(new_n1283), .A3(new_n1291), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(G2897), .A3(new_n1270), .A4(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1270), .A2(G2897), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1294), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1292), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1237), .A2(G378), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1274), .A2(new_n1271), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT62), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT62), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .A4(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1300), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1020), .B(new_n1051), .C1(new_n1123), .C2(new_n1125), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1264), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n850), .B1(new_n1064), .B2(new_n1092), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1310), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1312), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(KEYINPUT126), .A3(new_n1264), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1309), .B1(new_n1316), .B2(KEYINPUT127), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1126), .A2(new_n1052), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1309), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT127), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1319), .A2(new_n1320), .A3(new_n1313), .A4(new_n1315), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1317), .A2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1056), .A2(G390), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1316), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1308), .A2(new_n1325), .ZN(new_n1326));
  AOI22_X1  g1126(.A1(new_n1317), .A2(new_n1321), .B1(new_n1323), .B2(new_n1316), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1304), .A2(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .A4(KEYINPUT63), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1327), .A2(new_n1300), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(G405));
  AND3_X1   g1132(.A1(new_n1266), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1303), .B1(new_n1266), .B2(new_n1301), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1325), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1266), .A2(new_n1301), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1303), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1266), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1338), .A2(new_n1327), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1335), .A2(new_n1340), .ZN(G402));
endmodule


