

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776;

  AND2_X1 U364 ( .A1(n389), .A2(n387), .ZN(n379) );
  INV_X1 U365 ( .A(n584), .ZN(n577) );
  XNOR2_X1 U366 ( .A(n762), .B(G146), .ZN(n495) );
  INV_X1 U367 ( .A(G128), .ZN(n375) );
  INV_X1 U368 ( .A(G953), .ZN(n767) );
  XNOR2_X1 U369 ( .A(n485), .B(n495), .ZN(n664) );
  AND2_X2 U370 ( .A1(n525), .A2(n577), .ZN(n566) );
  XNOR2_X2 U371 ( .A(n489), .B(n425), .ZN(n755) );
  XNOR2_X2 U372 ( .A(n423), .B(n422), .ZN(n489) );
  AND2_X2 U373 ( .A1(n403), .A2(n398), .ZN(n397) );
  XOR2_X2 U374 ( .A(KEYINPUT78), .B(n607), .Z(n688) );
  NAND2_X2 U375 ( .A1(n635), .A2(n626), .ZN(n766) );
  XNOR2_X2 U376 ( .A(KEYINPUT72), .B(G110), .ZN(n420) );
  INV_X1 U377 ( .A(G210), .ZN(n373) );
  XNOR2_X1 U378 ( .A(n394), .B(G119), .ZN(n423) );
  XNOR2_X1 U379 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n616) );
  NOR2_X1 U380 ( .A1(n615), .A2(n690), .ZN(n368) );
  NAND2_X1 U381 ( .A1(n753), .A2(n488), .ZN(n345) );
  NAND2_X1 U382 ( .A1(n343), .A2(n344), .ZN(n346) );
  NAND2_X1 U383 ( .A1(n345), .A2(n346), .ZN(n480) );
  INV_X1 U384 ( .A(n753), .ZN(n343) );
  INV_X1 U385 ( .A(n488), .ZN(n344) );
  XNOR2_X1 U386 ( .A(n418), .B(n433), .ZN(n753) );
  BUF_X1 U387 ( .A(n664), .Z(n347) );
  XNOR2_X1 U388 ( .A(n348), .B(n349), .ZN(n567) );
  NOR2_X1 U389 ( .A1(n668), .A2(n630), .ZN(n348) );
  NAND2_X1 U390 ( .A1(n437), .A2(G210), .ZN(n349) );
  XNOR2_X1 U391 ( .A(n592), .B(KEYINPUT19), .ZN(n604) );
  INV_X1 U392 ( .A(G237), .ZN(n436) );
  INV_X1 U393 ( .A(n705), .ZN(n414) );
  INV_X1 U394 ( .A(n717), .ZN(n382) );
  XNOR2_X1 U395 ( .A(n417), .B(KEYINPUT64), .ZN(n763) );
  INV_X1 U396 ( .A(KEYINPUT4), .ZN(n417) );
  XNOR2_X1 U397 ( .A(n479), .B(G137), .ZN(n762) );
  INV_X1 U398 ( .A(KEYINPUT65), .ZN(n402) );
  NAND2_X1 U399 ( .A1(n401), .A2(n399), .ZN(n398) );
  NAND2_X1 U400 ( .A1(n473), .A2(n402), .ZN(n401) );
  NAND2_X1 U401 ( .A1(n630), .A2(n400), .ZN(n399) );
  NAND2_X1 U402 ( .A1(KEYINPUT2), .A2(n402), .ZN(n400) );
  INV_X1 U403 ( .A(KEYINPUT111), .ZN(n565) );
  XNOR2_X1 U404 ( .A(n564), .B(KEYINPUT30), .ZN(n370) );
  XNOR2_X1 U405 ( .A(G113), .B(KEYINPUT69), .ZN(n422) );
  XOR2_X1 U406 ( .A(G140), .B(G110), .Z(n506) );
  XNOR2_X1 U407 ( .A(G137), .B(G128), .ZN(n505) );
  XNOR2_X1 U408 ( .A(n504), .B(n350), .ZN(n508) );
  XNOR2_X1 U409 ( .A(n582), .B(n364), .ZN(n728) );
  INV_X1 U410 ( .A(KEYINPUT41), .ZN(n364) );
  AND2_X1 U411 ( .A1(n406), .A2(n414), .ZN(n405) );
  NOR2_X1 U412 ( .A1(n392), .A2(n391), .ZN(n390) );
  INV_X1 U413 ( .A(KEYINPUT22), .ZN(n385) );
  INV_X1 U414 ( .A(G146), .ZN(n426) );
  INV_X1 U415 ( .A(KEYINPUT106), .ZN(n381) );
  NAND2_X1 U416 ( .A1(G234), .A2(G237), .ZN(n439) );
  XNOR2_X1 U417 ( .A(G113), .B(G122), .ZN(n448) );
  XNOR2_X1 U418 ( .A(G143), .B(G104), .ZN(n451) );
  NOR2_X1 U419 ( .A1(G953), .A2(G237), .ZN(n447) );
  XOR2_X1 U420 ( .A(G131), .B(G140), .Z(n481) );
  XNOR2_X1 U421 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n428) );
  XOR2_X1 U422 ( .A(KEYINPUT96), .B(n519), .Z(n707) );
  XNOR2_X1 U423 ( .A(n763), .B(n416), .ZN(n488) );
  XNOR2_X1 U424 ( .A(n432), .B(KEYINPUT66), .ZN(n416) );
  XNOR2_X1 U425 ( .A(KEYINPUT5), .B(G131), .ZN(n491) );
  XNOR2_X1 U426 ( .A(n420), .B(n419), .ZN(n418) );
  INV_X1 U427 ( .A(KEYINPUT89), .ZN(n419) );
  XNOR2_X1 U428 ( .A(KEYINPUT16), .B(G122), .ZN(n424) );
  INV_X1 U429 ( .A(G134), .ZN(n458) );
  XNOR2_X1 U430 ( .A(G116), .B(G107), .ZN(n460) );
  XOR2_X1 U431 ( .A(KEYINPUT102), .B(G122), .Z(n461) );
  XOR2_X1 U432 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n463) );
  NAND2_X1 U433 ( .A1(n396), .A2(n354), .ZN(n395) );
  XNOR2_X1 U434 ( .A(n393), .B(n438), .ZN(n592) );
  NOR2_X1 U435 ( .A1(n370), .A2(n586), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n566), .B(n565), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n508), .B(n507), .ZN(n513) );
  XNOR2_X1 U438 ( .A(KEYINPUT42), .B(n356), .ZN(n775) );
  XOR2_X1 U439 ( .A(KEYINPUT32), .B(n352), .Z(n650) );
  NOR2_X1 U440 ( .A1(n542), .A2(n587), .ZN(n365) );
  INV_X1 U441 ( .A(n358), .ZN(n646) );
  NAND2_X1 U442 ( .A1(n408), .A2(n409), .ZN(n678) );
  AND2_X1 U443 ( .A1(n411), .A2(n414), .ZN(n410) );
  NOR2_X1 U444 ( .A1(n388), .A2(n695), .ZN(n387) );
  NOR2_X1 U445 ( .A1(n501), .A2(KEYINPUT83), .ZN(n388) );
  XOR2_X1 U446 ( .A(n421), .B(n503), .Z(n350) );
  OR2_X1 U447 ( .A1(n743), .A2(G902), .ZN(n351) );
  AND2_X1 U448 ( .A1(n386), .A2(n365), .ZN(n352) );
  XNOR2_X1 U449 ( .A(n513), .B(n512), .ZN(n743) );
  XOR2_X1 U450 ( .A(n638), .B(n637), .Z(n353) );
  AND2_X1 U451 ( .A1(n630), .A2(n402), .ZN(n354) );
  AND2_X1 U452 ( .A1(n628), .A2(KEYINPUT65), .ZN(n355) );
  INV_X1 U453 ( .A(KEYINPUT83), .ZN(n391) );
  AND2_X1 U454 ( .A1(n728), .A2(n606), .ZN(n356) );
  XNOR2_X1 U455 ( .A(n522), .B(n359), .ZN(n358) );
  AND2_X1 U456 ( .A1(n379), .A2(n380), .ZN(n357) );
  NAND2_X1 U457 ( .A1(n379), .A2(n380), .ZN(n384) );
  XNOR2_X1 U458 ( .A(n570), .B(n569), .ZN(n617) );
  NAND2_X1 U459 ( .A1(n617), .A2(n687), .ZN(n572) );
  XOR2_X1 U460 ( .A(n521), .B(KEYINPUT97), .Z(n359) );
  NAND2_X1 U461 ( .A1(n412), .A2(n410), .ZN(n409) );
  NAND2_X1 U462 ( .A1(n407), .A2(n405), .ZN(n408) );
  XNOR2_X2 U463 ( .A(n360), .B(n361), .ZN(n653) );
  NAND2_X1 U464 ( .A1(n537), .A2(n597), .ZN(n360) );
  XOR2_X1 U465 ( .A(KEYINPUT77), .B(KEYINPUT35), .Z(n361) );
  NOR2_X2 U466 ( .A1(n600), .A2(n581), .ZN(n570) );
  NAND2_X1 U467 ( .A1(n545), .A2(n391), .ZN(n380) );
  NAND2_X1 U468 ( .A1(n378), .A2(n382), .ZN(n377) );
  NAND2_X1 U469 ( .A1(n377), .A2(n384), .ZN(n376) );
  XNOR2_X2 U470 ( .A(n362), .B(KEYINPUT74), .ZN(n600) );
  NAND2_X1 U471 ( .A1(n369), .A2(n371), .ZN(n362) );
  INV_X1 U472 ( .A(n386), .ZN(n545) );
  XNOR2_X2 U473 ( .A(n478), .B(n385), .ZN(n386) );
  XNOR2_X1 U474 ( .A(n496), .B(n495), .ZN(n638) );
  XNOR2_X2 U475 ( .A(n498), .B(G472), .ZN(n574) );
  NOR2_X2 U476 ( .A1(n776), .A2(n775), .ZN(n363) );
  XNOR2_X2 U477 ( .A(n572), .B(n571), .ZN(n776) );
  XNOR2_X2 U478 ( .A(n559), .B(KEYINPUT45), .ZN(n631) );
  NAND2_X2 U479 ( .A1(n631), .A2(n627), .ZN(n629) );
  NAND2_X1 U480 ( .A1(n358), .A2(n383), .ZN(n378) );
  XNOR2_X1 U481 ( .A(n376), .B(n381), .ZN(n539) );
  XNOR2_X1 U482 ( .A(n363), .B(KEYINPUT46), .ZN(n367) );
  NOR2_X2 U483 ( .A1(n734), .A2(n733), .ZN(n735) );
  OR2_X2 U484 ( .A1(n747), .A2(n636), .ZN(n693) );
  NOR2_X2 U485 ( .A1(n675), .A2(n746), .ZN(n677) );
  XNOR2_X2 U486 ( .A(n366), .B(n616), .ZN(n635) );
  NAND2_X1 U487 ( .A1(n368), .A2(n367), .ZN(n366) );
  AND2_X2 U488 ( .A1(n404), .A2(n693), .ZN(n662) );
  AND2_X1 U489 ( .A1(n404), .A2(n372), .ZN(n674) );
  NOR2_X1 U490 ( .A1(n374), .A2(n373), .ZN(n372) );
  INV_X1 U491 ( .A(n693), .ZN(n374) );
  XNOR2_X2 U492 ( .A(n459), .B(n458), .ZN(n479) );
  XNOR2_X2 U493 ( .A(n375), .B(G143), .ZN(n459) );
  INV_X1 U494 ( .A(n678), .ZN(n383) );
  NAND2_X1 U495 ( .A1(n386), .A2(n390), .ZN(n389) );
  INV_X1 U496 ( .A(n501), .ZN(n392) );
  NAND2_X1 U497 ( .A1(n567), .A2(n712), .ZN(n393) );
  XNOR2_X2 U498 ( .A(G116), .B(KEYINPUT3), .ZN(n394) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n668) );
  NAND2_X1 U500 ( .A1(n629), .A2(n628), .ZN(n694) );
  NAND2_X1 U501 ( .A1(n397), .A2(n395), .ZN(n404) );
  INV_X1 U502 ( .A(n629), .ZN(n396) );
  NAND2_X1 U503 ( .A1(n629), .A2(n355), .ZN(n403) );
  NAND2_X1 U504 ( .A1(n413), .A2(n415), .ZN(n406) );
  NAND2_X1 U505 ( .A1(n412), .A2(n413), .ZN(n407) );
  NOR2_X1 U506 ( .A1(n526), .A2(KEYINPUT95), .ZN(n411) );
  INV_X1 U507 ( .A(n527), .ZN(n412) );
  NAND2_X1 U508 ( .A1(n526), .A2(KEYINPUT95), .ZN(n413) );
  INV_X1 U509 ( .A(KEYINPUT95), .ZN(n415) );
  AND2_X1 U510 ( .A1(n699), .A2(n500), .ZN(n501) );
  NOR2_X2 U511 ( .A1(n698), .A2(n699), .ZN(n530) );
  INV_X1 U512 ( .A(n631), .ZN(n747) );
  XNOR2_X1 U513 ( .A(n480), .B(n484), .ZN(n485) );
  XOR2_X1 U514 ( .A(KEYINPUT24), .B(KEYINPUT93), .Z(n421) );
  INV_X1 U515 ( .A(KEYINPUT71), .ZN(n613) );
  XNOR2_X1 U516 ( .A(n494), .B(n493), .ZN(n496) );
  XNOR2_X1 U517 ( .A(n515), .B(KEYINPUT25), .ZN(n516) );
  INV_X1 U518 ( .A(n746), .ZN(n641) );
  XNOR2_X1 U519 ( .A(n424), .B(KEYINPUT70), .ZN(n425) );
  XNOR2_X1 U520 ( .A(n426), .B(G125), .ZN(n446) );
  XNOR2_X1 U521 ( .A(n446), .B(n459), .ZN(n430) );
  NAND2_X1 U522 ( .A1(n767), .A2(G224), .ZN(n427) );
  XNOR2_X1 U523 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U524 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U525 ( .A(n755), .B(n431), .ZN(n435) );
  INV_X1 U526 ( .A(G101), .ZN(n432) );
  XNOR2_X1 U527 ( .A(G107), .B(G104), .ZN(n433) );
  INV_X1 U528 ( .A(n480), .ZN(n434) );
  XNOR2_X1 U529 ( .A(G902), .B(KEYINPUT15), .ZN(n473) );
  INV_X1 U530 ( .A(n473), .ZN(n630) );
  INV_X1 U531 ( .A(G902), .ZN(n497) );
  NAND2_X1 U532 ( .A1(n497), .A2(n436), .ZN(n437) );
  NAND2_X1 U533 ( .A1(n437), .A2(G214), .ZN(n712) );
  INV_X1 U534 ( .A(KEYINPUT86), .ZN(n438) );
  XNOR2_X1 U535 ( .A(n439), .B(KEYINPUT14), .ZN(n442) );
  NAND2_X1 U536 ( .A1(G902), .A2(n442), .ZN(n560) );
  XOR2_X1 U537 ( .A(G898), .B(KEYINPUT90), .Z(n750) );
  NAND2_X1 U538 ( .A1(n750), .A2(G953), .ZN(n440) );
  XOR2_X1 U539 ( .A(KEYINPUT91), .B(n440), .Z(n756) );
  NOR2_X1 U540 ( .A1(n560), .A2(n756), .ZN(n441) );
  XNOR2_X1 U541 ( .A(n441), .B(KEYINPUT92), .ZN(n443) );
  NAND2_X1 U542 ( .A1(G952), .A2(n442), .ZN(n726) );
  NOR2_X1 U543 ( .A1(n726), .A2(G953), .ZN(n563) );
  NOR2_X1 U544 ( .A1(n443), .A2(n563), .ZN(n444) );
  NOR2_X2 U545 ( .A1(n604), .A2(n444), .ZN(n445) );
  XNOR2_X2 U546 ( .A(n445), .B(KEYINPUT0), .ZN(n523) );
  XNOR2_X1 U547 ( .A(KEYINPUT13), .B(G475), .ZN(n457) );
  XNOR2_X1 U548 ( .A(n446), .B(KEYINPUT10), .ZN(n509) );
  XNOR2_X1 U549 ( .A(n481), .B(n509), .ZN(n761) );
  XOR2_X1 U550 ( .A(KEYINPUT73), .B(n447), .Z(n490) );
  NAND2_X1 U551 ( .A1(G214), .A2(n490), .ZN(n454) );
  XOR2_X1 U552 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n449) );
  XNOR2_X1 U553 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U554 ( .A(n450), .B(KEYINPUT12), .Z(n452) );
  XNOR2_X1 U555 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U556 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U557 ( .A(n761), .B(n455), .ZN(n656) );
  NOR2_X1 U558 ( .A1(G902), .A2(n656), .ZN(n456) );
  XNOR2_X1 U559 ( .A(n457), .B(n456), .ZN(n535) );
  XNOR2_X1 U560 ( .A(n461), .B(n460), .ZN(n465) );
  XNOR2_X1 U561 ( .A(KEYINPUT9), .B(KEYINPUT100), .ZN(n462) );
  XNOR2_X1 U562 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U563 ( .A(n465), .B(n464), .Z(n468) );
  NAND2_X1 U564 ( .A1(G234), .A2(n767), .ZN(n466) );
  XOR2_X1 U565 ( .A(KEYINPUT8), .B(n466), .Z(n502) );
  NAND2_X1 U566 ( .A1(G217), .A2(n502), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U568 ( .A(n479), .B(n469), .ZN(n738) );
  NOR2_X1 U569 ( .A1(n738), .A2(G902), .ZN(n471) );
  INV_X1 U570 ( .A(G478), .ZN(n470) );
  XNOR2_X1 U571 ( .A(n471), .B(n470), .ZN(n536) );
  NOR2_X1 U572 ( .A1(n535), .A2(n536), .ZN(n472) );
  XNOR2_X1 U573 ( .A(n472), .B(KEYINPUT103), .ZN(n715) );
  NAND2_X1 U574 ( .A1(G234), .A2(n473), .ZN(n474) );
  XNOR2_X1 U575 ( .A(KEYINPUT20), .B(n474), .ZN(n514) );
  NAND2_X1 U576 ( .A1(G221), .A2(n514), .ZN(n475) );
  XNOR2_X1 U577 ( .A(KEYINPUT21), .B(n475), .ZN(n696) );
  XNOR2_X1 U578 ( .A(KEYINPUT94), .B(n696), .ZN(n524) );
  NOR2_X1 U579 ( .A1(n715), .A2(n524), .ZN(n476) );
  XNOR2_X1 U580 ( .A(n476), .B(KEYINPUT104), .ZN(n477) );
  NAND2_X1 U581 ( .A1(n523), .A2(n477), .ZN(n478) );
  XOR2_X1 U582 ( .A(n481), .B(KEYINPUT76), .Z(n483) );
  NAND2_X1 U583 ( .A1(G227), .A2(n767), .ZN(n482) );
  XNOR2_X1 U584 ( .A(n483), .B(n482), .ZN(n484) );
  NAND2_X1 U585 ( .A1(n664), .A2(n497), .ZN(n487) );
  XOR2_X1 U586 ( .A(KEYINPUT68), .B(G469), .Z(n486) );
  XNOR2_X2 U587 ( .A(n487), .B(n486), .ZN(n579) );
  XNOR2_X2 U588 ( .A(n579), .B(KEYINPUT1), .ZN(n699) );
  XNOR2_X1 U589 ( .A(n489), .B(n488), .ZN(n494) );
  NAND2_X1 U590 ( .A1(n490), .A2(G210), .ZN(n492) );
  XNOR2_X1 U591 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U592 ( .A1(n638), .A2(n497), .ZN(n498) );
  INV_X1 U593 ( .A(KEYINPUT6), .ZN(n499) );
  XNOR2_X1 U594 ( .A(n574), .B(n499), .ZN(n587) );
  INV_X1 U595 ( .A(n587), .ZN(n500) );
  NAND2_X1 U596 ( .A1(G221), .A2(n502), .ZN(n504) );
  XNOR2_X1 U597 ( .A(G119), .B(KEYINPUT23), .ZN(n503) );
  XNOR2_X1 U598 ( .A(n506), .B(n505), .ZN(n507) );
  INV_X1 U599 ( .A(n509), .ZN(n510) );
  XNOR2_X1 U600 ( .A(n510), .B(KEYINPUT81), .ZN(n511) );
  XNOR2_X1 U601 ( .A(n511), .B(KEYINPUT75), .ZN(n512) );
  NAND2_X1 U602 ( .A1(G217), .A2(n514), .ZN(n515) );
  XNOR2_X2 U603 ( .A(n351), .B(n516), .ZN(n584) );
  INV_X1 U604 ( .A(KEYINPUT105), .ZN(n517) );
  XNOR2_X1 U605 ( .A(n584), .B(n517), .ZN(n695) );
  INV_X1 U606 ( .A(n524), .ZN(n518) );
  NAND2_X1 U607 ( .A1(n577), .A2(n518), .ZN(n698) );
  BUF_X1 U608 ( .A(n574), .Z(n705) );
  NAND2_X1 U609 ( .A1(n530), .A2(n705), .ZN(n519) );
  BUF_X1 U610 ( .A(n523), .Z(n520) );
  NAND2_X1 U611 ( .A1(n707), .A2(n520), .ZN(n522) );
  XOR2_X1 U612 ( .A(KEYINPUT98), .B(KEYINPUT31), .Z(n521) );
  INV_X1 U613 ( .A(n523), .ZN(n527) );
  NOR2_X1 U614 ( .A1(n524), .A2(n579), .ZN(n525) );
  INV_X1 U615 ( .A(n566), .ZN(n526) );
  INV_X1 U616 ( .A(n535), .ZN(n528) );
  AND2_X1 U617 ( .A1(n536), .A2(n528), .ZN(n684) );
  INV_X1 U618 ( .A(n684), .ZN(n529) );
  OR2_X1 U619 ( .A1(n536), .A2(n528), .ZN(n589) );
  AND2_X1 U620 ( .A1(n529), .A2(n589), .ZN(n717) );
  XNOR2_X1 U621 ( .A(n530), .B(KEYINPUT108), .ZN(n531) );
  NAND2_X1 U622 ( .A1(n531), .A2(n587), .ZN(n532) );
  XNOR2_X2 U623 ( .A(n532), .B(KEYINPUT33), .ZN(n729) );
  NAND2_X1 U624 ( .A1(n729), .A2(n520), .ZN(n534) );
  INV_X1 U625 ( .A(KEYINPUT34), .ZN(n533) );
  XNOR2_X1 U626 ( .A(n534), .B(n533), .ZN(n537) );
  AND2_X1 U627 ( .A1(n536), .A2(n535), .ZN(n597) );
  NAND2_X1 U628 ( .A1(n653), .A2(KEYINPUT44), .ZN(n538) );
  NAND2_X1 U629 ( .A1(n539), .A2(n538), .ZN(n541) );
  INV_X1 U630 ( .A(KEYINPUT84), .ZN(n540) );
  XNOR2_X1 U631 ( .A(n541), .B(n540), .ZN(n558) );
  INV_X1 U632 ( .A(n699), .ZN(n619) );
  NAND2_X1 U633 ( .A1(n619), .A2(n695), .ZN(n542) );
  NOR2_X1 U634 ( .A1(n577), .A2(n705), .ZN(n543) );
  NAND2_X1 U635 ( .A1(n699), .A2(n543), .ZN(n544) );
  NOR2_X1 U636 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U637 ( .A(n546), .B(KEYINPUT107), .ZN(n645) );
  NAND2_X1 U638 ( .A1(n650), .A2(n645), .ZN(n553) );
  INV_X1 U639 ( .A(n553), .ZN(n550) );
  INV_X1 U640 ( .A(n653), .ZN(n548) );
  NOR2_X1 U641 ( .A1(KEYINPUT85), .A2(KEYINPUT44), .ZN(n547) );
  NAND2_X1 U642 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U643 ( .A1(n550), .A2(n549), .ZN(n556) );
  INV_X1 U644 ( .A(KEYINPUT85), .ZN(n551) );
  NOR2_X1 U645 ( .A1(n653), .A2(n551), .ZN(n552) );
  NOR2_X1 U646 ( .A1(n552), .A2(KEYINPUT44), .ZN(n554) );
  NAND2_X1 U647 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U648 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U649 ( .A1(n558), .A2(n557), .ZN(n559) );
  OR2_X1 U650 ( .A1(n767), .A2(n560), .ZN(n561) );
  NOR2_X1 U651 ( .A1(G900), .A2(n561), .ZN(n562) );
  NOR2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n574), .A2(n712), .ZN(n564) );
  BUF_X1 U654 ( .A(n567), .Z(n598) );
  INV_X1 U655 ( .A(n598), .ZN(n622) );
  INV_X1 U656 ( .A(KEYINPUT38), .ZN(n568) );
  XNOR2_X1 U657 ( .A(n622), .B(n568), .ZN(n581) );
  INV_X1 U658 ( .A(KEYINPUT39), .ZN(n569) );
  INV_X1 U659 ( .A(n589), .ZN(n687) );
  INV_X1 U660 ( .A(KEYINPUT40), .ZN(n571) );
  INV_X1 U661 ( .A(n696), .ZN(n583) );
  INV_X1 U662 ( .A(n586), .ZN(n573) );
  AND2_X1 U663 ( .A1(n583), .A2(n573), .ZN(n575) );
  NAND2_X1 U664 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U665 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U666 ( .A(KEYINPUT28), .B(n578), .Z(n580) );
  NOR2_X1 U667 ( .A1(n580), .A2(n579), .ZN(n606) );
  INV_X1 U668 ( .A(n581), .ZN(n713) );
  NAND2_X1 U669 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U670 ( .A1(n716), .A2(n715), .ZN(n582) );
  NAND2_X1 U671 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U672 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U673 ( .A1(n588), .A2(n587), .ZN(n590) );
  NOR2_X1 U674 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U675 ( .A(n591), .B(KEYINPUT109), .ZN(n618) );
  INV_X1 U676 ( .A(n618), .ZN(n594) );
  BUF_X1 U677 ( .A(n592), .Z(n593) );
  NAND2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U679 ( .A(n595), .B(KEYINPUT36), .ZN(n596) );
  NOR2_X1 U680 ( .A1(n699), .A2(n596), .ZN(n690) );
  NAND2_X1 U681 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X2 U682 ( .A1(n600), .A2(n599), .ZN(n651) );
  INV_X1 U683 ( .A(n651), .ZN(n602) );
  NAND2_X1 U684 ( .A1(n717), .A2(KEYINPUT47), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U686 ( .A(KEYINPUT80), .B(n603), .Z(n612) );
  INV_X1 U687 ( .A(KEYINPUT47), .ZN(n608) );
  INV_X1 U688 ( .A(n604), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U690 ( .A(n608), .B(n688), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n608), .A2(n717), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n614), .B(n613), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n617), .A2(n684), .ZN(n692) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n620), .A2(n712), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n621), .B(KEYINPUT43), .ZN(n623) );
  AND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n625) );
  INV_X1 U700 ( .A(KEYINPUT110), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n625), .B(n624), .ZN(n774) );
  AND2_X1 U702 ( .A1(n692), .A2(n774), .ZN(n626) );
  INV_X1 U703 ( .A(n766), .ZN(n627) );
  INV_X1 U704 ( .A(KEYINPUT2), .ZN(n628) );
  NAND2_X1 U705 ( .A1(KEYINPUT2), .A2(n692), .ZN(n632) );
  XNOR2_X1 U706 ( .A(KEYINPUT79), .B(n632), .ZN(n633) );
  AND2_X1 U707 ( .A1(n633), .A2(n774), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n662), .A2(G472), .ZN(n639) );
  XOR2_X1 U710 ( .A(KEYINPUT112), .B(KEYINPUT62), .Z(n637) );
  XNOR2_X1 U711 ( .A(n639), .B(n353), .ZN(n642) );
  INV_X1 U712 ( .A(G952), .ZN(n640) );
  AND2_X1 U713 ( .A1(n640), .A2(G953), .ZN(n746) );
  NAND2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U716 ( .A(G110), .B(KEYINPUT115), .Z(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(G12) );
  NAND2_X1 U718 ( .A1(n646), .A2(n687), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(G113), .ZN(G15) );
  NAND2_X1 U720 ( .A1(n646), .A2(n684), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n648), .B(G116), .ZN(G18) );
  XNOR2_X1 U722 ( .A(G101), .B(KEYINPUT113), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n357), .B(n649), .ZN(G3) );
  XNOR2_X1 U724 ( .A(n650), .B(G119), .ZN(G21) );
  XNOR2_X1 U725 ( .A(G143), .B(KEYINPUT116), .ZN(n652) );
  XOR2_X1 U726 ( .A(n652), .B(n651), .Z(G45) );
  XOR2_X1 U727 ( .A(n653), .B(G122), .Z(G24) );
  NAND2_X1 U728 ( .A1(n662), .A2(G475), .ZN(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT88), .B(KEYINPUT123), .ZN(n654) );
  XOR2_X1 U730 ( .A(n654), .B(KEYINPUT59), .Z(n655) );
  XNOR2_X1 U731 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n659), .A2(n641), .ZN(n661) );
  INV_X1 U734 ( .A(KEYINPUT60), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n661), .B(n660), .ZN(G60) );
  BUF_X2 U736 ( .A(n662), .Z(n742) );
  NAND2_X1 U737 ( .A1(n742), .A2(G469), .ZN(n666) );
  XNOR2_X1 U738 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n347), .B(n663), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U741 ( .A1(n667), .A2(n746), .ZN(G54) );
  BUF_X1 U742 ( .A(n668), .Z(n672) );
  XOR2_X1 U743 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n670) );
  XNOR2_X1 U744 ( .A(KEYINPUT87), .B(KEYINPUT55), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U746 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U747 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U748 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n676) );
  XNOR2_X1 U749 ( .A(n677), .B(n676), .ZN(G51) );
  NAND2_X1 U750 ( .A1(n678), .A2(n687), .ZN(n679) );
  XNOR2_X1 U751 ( .A(n679), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U752 ( .A(G104), .B(n680), .ZN(G6) );
  NAND2_X1 U753 ( .A1(n678), .A2(n684), .ZN(n682) );
  XOR2_X1 U754 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n681) );
  XNOR2_X1 U755 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U756 ( .A(G107), .B(n683), .ZN(G9) );
  XOR2_X1 U757 ( .A(G128), .B(KEYINPUT29), .Z(n686) );
  NAND2_X1 U758 ( .A1(n684), .A2(n688), .ZN(n685) );
  XNOR2_X1 U759 ( .A(n686), .B(n685), .ZN(G30) );
  NAND2_X1 U760 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U761 ( .A(n689), .B(G146), .ZN(G48) );
  XNOR2_X1 U762 ( .A(G125), .B(n690), .ZN(n691) );
  XNOR2_X1 U763 ( .A(n691), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U764 ( .A(G134), .B(n692), .ZN(G36) );
  AND2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n734) );
  INV_X1 U766 ( .A(n728), .ZN(n711) );
  NAND2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U768 ( .A(KEYINPUT49), .B(n697), .Z(n703) );
  XOR2_X1 U769 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n701) );
  NAND2_X1 U770 ( .A1(n698), .A2(n699), .ZN(n700) );
  XNOR2_X1 U771 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U775 ( .A(n708), .B(KEYINPUT118), .Z(n709) );
  XNOR2_X1 U776 ( .A(KEYINPUT51), .B(n709), .ZN(n710) );
  NOR2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n723) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n721) );
  INV_X1 U782 ( .A(n729), .ZN(n720) );
  NOR2_X1 U783 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U784 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U785 ( .A(n724), .B(KEYINPUT52), .ZN(n725) );
  NOR2_X1 U786 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U787 ( .A(n727), .B(KEYINPUT119), .ZN(n731) );
  NAND2_X1 U788 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U789 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U790 ( .A(n732), .B(KEYINPUT120), .ZN(n733) );
  XNOR2_X1 U791 ( .A(n735), .B(KEYINPUT121), .ZN(n736) );
  NOR2_X1 U792 ( .A1(G953), .A2(n736), .ZN(n737) );
  XNOR2_X1 U793 ( .A(KEYINPUT53), .B(n737), .ZN(G75) );
  NAND2_X1 U794 ( .A1(n742), .A2(G478), .ZN(n740) );
  XNOR2_X1 U795 ( .A(n738), .B(KEYINPUT124), .ZN(n739) );
  XNOR2_X1 U796 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U797 ( .A1(n746), .A2(n741), .ZN(G63) );
  NAND2_X1 U798 ( .A1(n742), .A2(G217), .ZN(n744) );
  XNOR2_X1 U799 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U800 ( .A1(n746), .A2(n745), .ZN(G66) );
  NOR2_X1 U801 ( .A1(n747), .A2(G953), .ZN(n752) );
  NAND2_X1 U802 ( .A1(G953), .A2(G224), .ZN(n748) );
  XOR2_X1 U803 ( .A(KEYINPUT61), .B(n748), .Z(n749) );
  NOR2_X1 U804 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U805 ( .A1(n752), .A2(n751), .ZN(n759) );
  XNOR2_X1 U806 ( .A(n753), .B(G101), .ZN(n754) );
  XNOR2_X1 U807 ( .A(n755), .B(n754), .ZN(n757) );
  NAND2_X1 U808 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(n760) );
  XOR2_X1 U810 ( .A(KEYINPUT125), .B(n760), .Z(G69) );
  XNOR2_X1 U811 ( .A(n761), .B(KEYINPUT126), .ZN(n765) );
  XNOR2_X1 U812 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U813 ( .A(n765), .B(n764), .ZN(n769) );
  XNOR2_X1 U814 ( .A(n766), .B(n769), .ZN(n768) );
  NAND2_X1 U815 ( .A1(n768), .A2(n767), .ZN(n773) );
  XNOR2_X1 U816 ( .A(G227), .B(n769), .ZN(n770) );
  NAND2_X1 U817 ( .A1(n770), .A2(G900), .ZN(n771) );
  NAND2_X1 U818 ( .A1(n771), .A2(G953), .ZN(n772) );
  NAND2_X1 U819 ( .A1(n773), .A2(n772), .ZN(G72) );
  XNOR2_X1 U820 ( .A(G140), .B(n774), .ZN(G42) );
  XOR2_X1 U821 ( .A(G137), .B(n775), .Z(G39) );
  XOR2_X1 U822 ( .A(n776), .B(G131), .Z(G33) );
endmodule

